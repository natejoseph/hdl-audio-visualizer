��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�p,f�9��+�<~ፘ�Q�ԁ2��eQ\����gP�T��J���£?oc@����T�Nr|\R�K�E��D}�I�z��i�)�}	S����L�={��H,��?��F
�Q��ݛr�I҆4�J�:f����<BeB/&�R������m[�4^�4bw1��r�>�
�I3£P�%/Ź���M���[�h�1�
߈�|t�e)J���i��opX����7*��.�y����P!C�������&�9��I`�nt6y��ϺC ��ʗ�훕oK.,�)u(5N�LǾQ4N�R)F��tRԋ3��qiI�!�^�$�u��iS�'�MŲ�����*ocƃw�]_��)��Q�+���%E�G�H�!�B]�$�ɅR�0��p�m�4E0�h��z��$4>렰�
�ߧ�X��:�]*D����1@�H�VNa�F�j��,�f��S��е��IA����2��1�i�s!��2ȃ���i�z�9'�������A�8�w���L��19b��_���Ȟ�>�`*Ͽߎ&-���_�'��Pj5	��Cc���~}o���eqF��N˘]ޝ'��?��X&�@���2P=��r��E�hɮw�?(���*�����[���@�;�����IQ���y�[T��co�U����3ȃ�*�H�O��@�f,n�I�'�j�Š�b����,�
�d�I)���]�l<�w��� �rՋ�"��e�z�[�$+���q��U�%�?�)�IϪoa�;V���� ��=�,G^F�FX��h�_�]F�~�nܾ���H*��r���Z�Rv��Ow�L)�	�ꡊ���o�"{����Y+���i�)�5P�8���K� ���p z_��&ɨ�'�L�A�bJ�	on��"@*t*��C�C>�`A�W�#ܮ�=����U���BT{��;�t�#鯇��Y�S�n{�d�m���מo��}7m����Q-pJE�^��0(�k�Avy	l)=W���;� t��T�U&CA�XX��RLN� ��c�|lQ�.�$r��7AC�$I��ŉ�Q��6�����*���������keS����UtK��d��E?���<EɄ��6R�јf~ҙ�����ӼQ�Ou7~��}�4��Qz��)FE�5c�ߚP[Rڊ�y�z���V�Hl&��0����Rڿ�D����K�Ѕt�}�	L��D����Ψ;z��O�)H��xܷ�Z�FP8����q��^��e��-S��팶Q -K5t?p?���##˖ (�件VÔ�[��˖K��]*��*. ��
�W�-ـ�{1ja����^_���Lڙ�m��p`G�B�v�_��,M���S7Z/�mM���A��xn�alf�I��x�鎯��j�9o�nZ�s��	��e��T|+������{��oLH�=>��S���,�ex@������C���(r|��*���%�O�T���T��ȷ�@w�%do/3���<"�5�v�k��@+��z�k_�X4���<�p�q*SLB��l�3�>�?#
�cf��;�p`�[��Є������]i,�Ъu#l����ڄ^�1��M��:�IRt廬�\���s����ar6�i�T��7��e&W}��$��Y	�	���`K�`�YO�t5E�L=L�O��yIY?p7S�=+[�j�s��+6<���<ޯ��D��ʝ4�h����|�88�])?r�:����r�E=�?�V��mꌭ��| J:#:�͛V���Ԏ �ӻ�o�~��Q�t��������P8ku�T��C�S�qP~�y{�Z(�4�I�}>�M�n�����g(u�R�CL�\pH!Y�� ��닔�І�B��^�h���&_A��S\�w���i���m���xpk�+SD�CUs��rP5�Q�f��c�> �9zE�����y֞閦�T_�]� n��ȣ�oi^�c�w*]��)���ѹ�,�U��F��(�BXk��HH��TOj�5���5��<� ����k{��a���L����g�5Ex��Q#���!�Fh�F����!拹�(�*��ľt���ȼLY�L�.�T�C��~<S��
�yO��Ԇ�J����õ�L�&Py��mS�*�p�YDh���`5�La�ϲ���EDĐ@}���v%Zd�������:��T��J�-�֜X���+���ѐ4�^t��&���T�c3u7!�}�w�$����
��;�~��>iӳ>�f;kE%��\�pH���Ș���sI�f"M��(E!���*�	�XMu��˂M��3��{ƌ�y��ƣ�
Qz����?_��0f�k]�_Y1�,�(���wy2.F�:�y<�O(��<��<�;����I6<�S�0��s�IC!�h�Í�ޚ���C>�0._�����e[l�NF�|NW�Ĺ)x�-�2U#Q!\�@5���:p�ЫA��U�c� ]�dT{��+�bVMG���7��ȢT�Z���Q���.��5H�o�-g/���h��d�w�	4&:�D�`=/�'`Q����ߠ7I���-��aDQ!t������L��av��N)��-	�!���'�:�¼V���T�b#��(r���V�wN����7e@6t���l0� C|�]ߐ�X����|�HOJ�(su$��-Ke�%B\���
�9uV��l�ŷ�	N<�{5C�A����]@��e%��{(j��VB����}���r�'luI0 'X�ڰEq��-˓\�0���bw_ m�������c%���u�uabr�����aD�DbV�}|���6�.�b��~^_7s9�ZX��͕詘���6dHG?�[6 Ua��u�:�'�?��r����֋Y`�v,�~2i���z���jktjj�<VV����f���0^;��z**��!��И���2��9.�}��6�o�R�00�&񐼶�I:=�Oj·֠���:/��E�e�Z���L%���.)@`4��/�p�y:c�bα%�8�#F2��a�f'�ю"���3��64�	�T;͖J�+P��r����Z<Rn��5ږny�e�h��l��ߞ���L���P��`�7J!���M�51�$u�'
xZ0s�B�ڎ�$<��>1|�a�k�Q��Aj2�N�R�;�hp��&��� ��/�W�T��HQ�l&y[A�<�pͧ�A	Cb)8u
���������R��0�#��ol���� P?|c2�Bw�=b�4�Ӳ��k�b/��@���HT���)mDG�T�ɓDL)P>��3,�m�G��CN�c7{3�|�c��&��^�/�����@�-�w�C@h�!]�
�Pd�r����*�Xv4n~�6L|])+�{��VK�6��͜��On������|y�'�>x2`�_����i��<�)�o�J�Y�"b�Ct��̟^��B�XP}Z~<�1 2d�nm5w�<�%�MΆB{�Z��Vy�CQ�Q.���Db?'���H=��j����%w�Vpp$T˪��Ў�ok��]!�L!�w��?`3�ƺ/P4S��� g~��g�S҈J���\�U���52W���d?ū)U��/�uCRF�>S�Tq�ר8�6�:sVaX%l�A���ܗ冪�|�KZ��e\/u!!���:��{�ڒ5γ^eZ��L��m��;	7�L "�~*+���`	���Ȭ�t�DI���˛�oKYɚM��߃<Y"	;z�%c����
���2|��£&����Oh޽�e�����I"�S�
+���0���0�(�FF�լnb#5�Vњ����j1�U*��S(���8G�jx%Ӊb��ou�h�����<0���"���<y�v��;[oSā�,n�u�I���e���Z^��rU�>N��#���zej��N�.��s�2EB�GU�x����%�B)c�@0�/{
bA"*Fݕ2?L�F�S,��3�j˼����(���[�t�oWƽ�V�u��	}e�t��(~�� ^!yj��ma줴�fR��<3���aY���2s7��D@Y��Ӈr�FV�o!����j�n#u��4�P�ē�C&$�8oÂ�K�@�j2�$�4�n����!'m�!�o*f-�S����Y��{JϒA�^G���٨�/�5�XF*{*fe�3J�z��@�������hѯ�ٲ��d�U�������<��יC���%J6Q��*�_�
�1�a�6�3N[�4����J�	q�S`�=�g�d��V��:�p}���A��cRh������Z��>���=�Ҁ)r�I�~PL˟��<������T����<-=�l߻ǒ��4��5q�꠻A��$�%�?�t������.�e�?��[��U(���χe�oX��6�����]�x��R���>���\���@Z�QLB(�*�F�b�G&/"���=:#d:����r,	!���Q:G��Z���3�����I҇�����j��D�	��i����=������>���J�o'���#�b��_
@6(H=k�7�"���?�6 ƃ�0�l*��X�����1)J�X�<G��0'V7��@�O��fp�$J�eQ����Y*�*/χ��u2'7YY�̐��F�W��8\�J��m��f`ix'�����Ս3i0�2�.�.@�r9�!7VG�~Z�Y
�dP)���q�,���B��q���Y��$��Qב�;�6��$T��?����%g��qPt� �Jż��B�2\W�P���<�^xޑ�gk�:�ޕ3�p�1�EP @��C�]������u��Ǟ��0��'�A.���
��O#)�eVLl��S�jx������[���C~_��H�����&h���{���XI`�� ^�����J�tF���6SuG6"��ۭ��H-�Z�n��0*�cZ� ��bn�5x&�m���|�]��}�ފ���=v}�~�ՓB.l�4�4�D	)���I�B�0
5�U�oD{���\����O�e�3�枷&�VIH�6�(9͵�8o�O�T�^΁~{ޱނC��:�킲tSS�9Q^B83v���ź�8f)��W�׌�R���� ��G~Q$Ar�dj��Ƹ�v) �#�n2�.B.�ˠ@�Д�n�v�N:�lD�"p��1�"g%'�.�ٖ����h��:�8Ѡ�����	�����t�봶#��[oشV�؀�ebP��d3�Ѧ���1x�K6Bq���vEy���>s�BU���J�or,A�I�յ�z�ΘV[��.�Ү�QiKp�ES/F�`)��+�T��ׯ@@,�F�S`��w�����v�!ͻ�My֌S.��$�H��`��yX�6lb���4|)%Ǖ��L�*��:̓�f��EB�T��t�|�a	�e{^|n���1����C�,dن.�v��^j��v�Lw�p�l��d/&}�������T�H�P�r�<��i&�A˹�P1n{�����6/��^�;J��Y�y��Fy�k�'��c`#�ɂh"��e:_�N.�r�V*����,��Z���U�<v�S97X�S	A��fY����(�MCx�@��d�\��[���ŧ�⃻��%�0��r--DwG�X�9|�5�h}�Iq���.�yn����,-��Y%D�u������L�b64�>�T Pڝ�&��wKa��(O)��M	q0��G<�4�lZ8�������?Z�Ϻm�l���dj�&�b5���dv��~�4�/�r�����AYZ�+jg���L�^�f�FqtDDm۾|*y�7w�����Ź�'�0��q��7��ͽ�.g��څ�q�;���U!=d!�H�hQ���hETs��A�]3����{x=0J���+�ޢ�B�3�.Q�^1D��6�.��Ea���.X�\]Ã�h>`���t?���ʵX�a1{ C�Ǒ�����@c�6e*���o�)�\�t�H.;=;�:���э��t 	�~�(�9�tR�9�rA�H:�
����s]b) .�����c��k?�gaG���ǐ᳊Aao3����y���%�� w������WI'�Cf���`1݌2q"P�$$8�d��GzK(yg�����6ޕ�}�p% ��|:'�*��*�؏�����cQʏ���5A�N1o+��B�Fh��0�����]N�=����9'� ����P�448Ĥ�JvP��O�O�8�|��U	��m��&@��3
?��P��"�.����;��&,.<��I���`��a{�9��h񘈸��Α�Ԧ�p��Y�b�������8�^`�_���*.9A�;J��Yt��9�����;�#���rۙ����5�D�Ӳ?��="sEd��]�䇱��m��l8V�k?�x�%�̴�6xR�����.%���R�o����`�Ĳ�O��肽�}+�|"��1��"K]����_�~>_��9���f,6��Jq]��5�������i��I�������m�/�h^D���o�|���N:	����`L��ڠ?Nt���	Ó\A�6;q<�\>#�/i�z�������Kb��Xl@%�=���ʭ�H�H��i,����� �
J�nG��Y�)�`�b>X��	+(|�d�S&�>�I�q�RD��"�[��8il��~RI�^��|�h.���P&�$��8�8�/�q�\�8��Zf�+]�p��UL�ymQ�*){�$�`6h0u��,?z(���,�n�Ҍ��2�6%�p&�e=�򴽠dA�hd�!����.ʁݨF�;|jRCr���gU�8�.���`ݺ8$� 8n~��^#"����h������x���*p���=R)���D�����Ur�a��,��\]آ�����
�m����T�����0�XY��a���d��ғP^@�{Q�p�$B07�]e�P=��hYx]�hA���v4�V2*�`/V��i��4���&�:)�Wk�E���3e��zٓ��U����xfNq/�$Y<��� ��:EE���P����u8i_,�������pК<J9AI$ɖ4  9���J�0�nĳA�H�d=dq�Pѥ1<��ݻoˁu���h��U�Kj�h<ނQ׹���Ou�a�>����������v��鴏��aǸ.Aǣ`��u�vŧO�rsa�b0-��$��S�&�?ȹ>�����fI&z�l������6|S���X�f�y�5�-��-����AmU�+�o����)�N����P�f����	�loZ���]�1��?%���w��_����\�/n%q�5�W����V�ۓ�o�!�H�2P̌r�%֛\��sL�W�g���Ja���$���	2��6��wB��Ro�B�n�系��ٹ�,b�3����GO`Q�"a�J�>-��$Zz�A�c��lB#ϝxI�q���Z#	xƶ#�bpA�}^|_�0%�;~�⹃)�F�Hq� ���I�$5-��}����I@Z�yy

 '2?�E�i�*��&c^�#�дX{s}`E�'��W���k��]Q�\-z+�7�̺7&t�G7�Z}�-���Lg�t;��c�vs:D_T�<##K���M�S@�yVT`4<L��s��k��tז	H�[���2�_