��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��,:��z��I�$^)BQ�}���T�xɥ�g)b]����������oCX�,n��4�cA~����qhL%H������[mPX��({'zR��e�y�c"��A{��[��(>nT��@���������Y����aCj2�W��=c�
�v�ۏ�||��y�$F�g0�{U&@���(���ҨT�tD�����"�}|�Pն���Q�?� �l������±�b�bi�Ʊ�Nxlu��#�(��]V��DR/����H�V�pU5]�2����T�!sf^���߷��1'�ڱ�Z ��z��������U�N�F�\��N�р�$���a��2��s�K\�m8�DT?.�J�Gh�#�o�/U7��W���W�TY�&4�8\P0�|gՀ'jK�����
Ӓ�߽���(o�d�Og#�џ��""�gd:wr��\ph���Si��(�#����5~%|�#xZ���N�Q��	r�g�CQq���ב��->�`�X#Kqo
��ܨ{� g�����@�`l���q�O\�C���"�+�]Зv���K���[8^����1��~1��O����Cy&�g��t�u hw��ඍy̽�d�ڈ��
[C��k����"|�>E͕Ҏq��>q?^����1��n-��A-��H�W���^r͢���5�tvG]2�r��Oy&��~҃��R>�[؜_���o�^ 	��+�Q⟵�1�`�̻1x|���>���
n+1CJ�eZ��%�l���|�Z *�`�M�D�D��4����M��%F�[��ME�:ܹ?��ӭ4ivVش�����տ?�Qb��%��*`�v��a�R�#�A�鼖�(o�C��g�t�p��>~�?y����z����J`]xB��Q�m��%��d��]�Ҫ��ۚd_�:ʛ6�&�1`����@����$��M�#� �伔����"����gpF�=S�p�-��f�Y��� �r��V�; 9�V�J ���]�~�7f��I~�������=+B��	L��� �����eϕg�Y;MΏh�#%���� ���6�]���À9�1V&dK��͵I�qx&���R�]b��B�> V��c*=�� �2(�q��o@�1�C���+�թ�9�d�x��?�S��<������GY�[�4?��+X��\ ������/A;�����au��s�G͐���s�\�T���#�aI&�'
.˸�\�c�;�H�5��>�+�υhO�����\����8ZQZJB���a6�����O��Asԏ���E��(�ֺ�"���O5�v��v�l4@�㎉��㓓OA��ʉq��%=�� ��ԭJ�M\`�1Ș2��kNJ ��_,� B(�~֏���<e�5���\HKb�����vĳ�J])��SI<7&{�˖f�斳��y����`��z⃙��ҨN��x�c�ˆ_�;9W���Lc����VR�V|zH5�`�W��!�$ι���J_;�R��,��_����5�s�]��P6_P�V�<���C��{E"��\�(�l����UI�Ŕ���uv��M�躋P�݌�?Zo��l��=v,%Ը1�wwB	���f>3�'�V��l�"V3.�#���ܗ]Q�f�}�g~�A�0��-t��x6s�`Q�Y��p�Cr$���9�-I�jB�7�9�`��Ju�
~|N����G�B"�?I\�^'�^���v,H��+�LMR�k6��f	�ٚ% ���r(��~;�/ �e�Ǫ������h����8w@��u��Io��]�|ݏxਫ਼��aPLy�&yڮ	�� �,A�ď���m���3$�V��\�����մY9ZK�$�$��$c�P��׈�׷P�������և���Ϥ�J>:qAN�Dr>�+�⍥���9�;߈B�ƫ�aB�-��}�i䁐>�0�P$/:	o�����p�[YӓO��.�Q�x?�s�"9�p�0�4Px��������G�V�	�O0�)��rU�s�e��d_Ȼ̯�`�GBM��u����[��:�E�1T�!)e�P�3�|�'A�)���u����m�Gm�@�_���/��=ͻ��dޢ^1�c�Aŧ۞N��4tM<�r��=md����.G�5
4D��HW�0%��)C~�H����fP�Q�v��e6���n�=t��i���ϙ�L�R��ׇ�:�@'P���4��u�J�b
�˰��J*���p=�ٻ������X|�I-������к*�`(�i	~Ni��A���(��^N�\n<�ڶp�1�����o�4��}�D��f�b Ü��0i�Ԝ�;���ׄ;�"��I�ϒ����9q��j	�>��c	]�	�|�K
��	,/%�Dz�T@ ��
dc�ޟ@\eր0�UnAu&g~`���O5J��v&(�Z9Ն�xU�a��N�:�͚(Z�4y,c]�+6?^�k+��B�������v��_c��m�xI��#g�s��̱_y�Q����	g�F���I��{B�����+��!���`Lޮ�TsL��r�$�!�{��-H�`l� 0��%}����X�O�i!�U��m0�f3�a�����H���C�=�v5�&�Wc����6��¶7͔&�!�N��Ġ�^���)(�;.�[�k�7w����؍�q���H��I�7'k�$��]����*AG	��9��i���MeG_�3�C�A�A?��Y�U��s5󑷵��m���6D�b�
���{Nub1mK��J���S�9�ф&���_ N��^ݹĵ�1�&F
a���ш���ߖ·�oa4�ǚ4wVa��O��<���l6��w��V\��ZhK%�Rq0��r�Y�^-�>��W�����6�!ˇ����8��r��o����U����AgPeE2����+����ɬ����+l�w���:���ɰ	#qX7Ht�ͳn���R��B&��1�s�nJ�i�xr��d$���ny�^?��U3�����X���L87�U�1E3;t��{_o�f�lk��h��ǵ.j�-y���&^IS6L�`+A�Tw��P¤�d���x�P�G�]H߳�xm���%{�|��l������]*A���[_�M(�$�?�GP��Ύm��;݌e�W�$���Y�O��jZ�]�8�.��S�;��zȈ���[�AI 9�HvnF
Ϻ�7��x�W��6�4�.'�֠ԌC�ו瘟�@J��)��?����K�E<�]���qf��ƣdT�x1�9���ԍ�B`Lz��[ǀܬ�TN��)J�P)��1�-��R����P!�r�]X��d���Bp���0�1�D��n�t5�R����>�H�g v�Ј���{�$q�\���"f�C����3���r#И�hr�f!���ۣ�W�G��^�^m棲M��\�_Ud�g��y��s*8�>ЙK$�P46��޹&p����IN�`�sD�'�4�,}��%O0m`���p����G�����`�Q�0n���lKR�g����[l�ʊ�N~�j�U���m�	���q6�yz���s�k�c嵐��c']�8=�mT�5N(�)"-V�$������nQ�PҴ�|ge��AN{���1&o�,�\�e��h"���gNԅv��.-�)��ؙVSܚ�l�R���G��򆀁�;3��Q'�^.��~�c��#�#y�1Zb�C�)���� 0f%����%S�;�=�Q%=�vI�k�<���I�T_���gT/���'7�ʰa�m��0m��e��,mН:��0JVI��˱��J�v�Q{�2���Y�3�z�|=�}3N��I@����/̤��2E��1�V�t����#'�&8���4V�\-����X��9����H�z�m�@�	��Nu��e0%�==�q���/R��k�˴,��o"�<\R&})�\��$�Y'^sM_�Z}dF �g`���X˾ΊM<��^�6�/?�慖�>g��v��]Wq5�]m3�?�KA�J��ʣ�W�)0��ۍ�^��X��K�C&Oؤ8�[,xV �ֵ��!�5wM,B�ϟ�8h���a�I��(��X2v'� ����zw�����u|�¹Q�(�Q �8G���j�u�0.�sԹR+�ΔZѭ����ZH���1Jp��W/�xFI<����Ϥd�ő�Fx�Z�0y mM�ޅ�Y�%w�X4 ˆ�}z�b9�˩F�"i�?�?:���x���T7���.:��C$|����JzR$��C�k�q(�.�]�g	�ۺ�C�HRE(�b��!���yEǰ]�gVx'F.ӱT>����ȯ�̒p�6Ͻ3E�c�>�E}�<��.l[ȵ���_IH�Y�[|C�C�?7'jwL�'U��n��ޯ���S����[���Ϩ&��oJn?�}���t�:I}�i�
=�Gc��D?��>Bq�%�=��J��,��P���^P���lG����ɯ���t5]�r�����i��bI2hg�g�TF6d��:"KP��A4c6'�{\x벀F���qPy �x�X���trȗ�OF�I��#��-�CV,t�3�I�|V5�	���#A_ *�E�Ԡ�yCV��wm�qM���(,�zK1��@�0��9�ʅ��֙--��:ŃaXW��T�v��y%����� o)fF<paL++��S��55�0>R-�l�0��G��78j0o����q[+"8��30R/$ӛ�t��Y�.��z��Y�|z�7%'h��B�Wv��=��۩奀���z.��
wU��`�ߘ���n{QmX4����1�~s�\[�c�L<C�кZK	���@tH]�@6�T�"��O�'���n�m�W����78=Ejd<t	8��3��d3Ff�l.K��mm��8�a�4 {uf{��TɒΧ�r����m�u[�˖�G��J��a��Mч�t%���I��(�Z�a3��ݖ(�_�L^�̦	d�ہ�Q�C4��ǔ�y����I0Z3߯Y�ag�W�t+�oF�Ӯ�C���k�hU��	,{0M�_��2h�F�����7`��#$�����F�	�C�²���D�u�Wۜ9��j��S���#�b�1VJ��l��9ޤ�%s�_��-d:W��#+vk�M�B��#l>������.�#��
�O�­�ƫޭ'2lc�pFy{�+������qR�M ��e�#��x� �p�5��th�f�N��z^ͬ�)�m��5�3~��1��}T�i]�۱�f�uqo��;�3ђxR8��s����e4����ƌ�]	��,�2F!� �cj������)֥��kĸv|�����)x�ܣ�d'L˚�@�����<����US�=&E=>E����ۗ�˴:ؔ8�u�6���]��_�$��-O��o�?���.�h �;��xX?���}6r�t�8J��j�@��%�fp8�ݐ���$(9�����kТ����>2D�yݴ�N؞#>�"�9�j	oX���Wf��
�Iy	cv���+��/����%��N���bop0���V��X��,1Їk�oF�uxԬ>���x:�Pf��~yH�Q_�����ED��r1�Z�P��ς۠�K��J?Ճ�k��,ܲz����^,���(�z�="q�RL�r��D�� �|��	���I�3-���8!���B$���m�;q�7������>
'���Ϭ�-N����{7kfrG޼"=)u��?�*Yi)`��Ke�U�Y�K$3��n;q��#��|��̰��m����mf��k E����R�~V;`�oE�Hsj����iE'h��ŞΓF�%`\�|��G�od�%���6C�g=�1���t�[�G�%cE�}Z��kUͅ���ġ^5�.q�u�م��xt��E̸���U�G�A	��{
=�&�������~Kw���F#�$*VF
�P�w�J(���Q]�C�!�����x'�&�Ȓy,σmI�|i'���i�}<�U`�/R.N�C5¨A��\��G��׸>N��T[{�+QO�rM�$z�ZM���9��k�zo ���Чe�5���5d�����T��]P4~��+��s��"H���"%!�z�K`�|'�_79��{����ܳ�~�s�M��eS��7�
n`��,����L���k~��bA�s�j��K�~��!�K���V�Z阰�b<��<I��C���.�Щ��k4C%�a{3�+o��e�*T=38�^������.ȫb��ř�-I���
9!d9��Iw����g�ݵԽm۳�^�֊D�DD���8�%��r=�R#�w�ry����Ɣ�a���(�_m�t�4x�f�yxI<p����?��y9�mC>F�����H��$���T���j0��zDY����pu��9���"}R�B��%,lo� �H[!����)�R+\~q'
N�|`�ͮ-u�6:J�MV��E}��9��}.t���a��6�虜vWH��K������t֕�M���;��*�S��,���^�=�sc�S|I�!T1���d�]����{�f �\OU�;ZI��h``��~n�z4:o�����YU
�>/��zHxm4ep�y1���NdO͌��"�q���˯(��SR2B|�qᤊ�OGJ�c��P_@�[b��U��Π|�;�e}�U�JU�w8�lK���$���&���y�>���e;B�vP��܊�fc�J�Y�i�˙I�y��_�x�mq��FĹ}�=&��s�񺟕�� �IIׂH��HPֽb�J�7z�6��)ܬ�͈x�O�$M��w~�!Q���0JD�����C�Ih�T���`v�f'O,u�U�0�;�6V�7R�U����+��8��v����C�ީL��5�k�ĸ*��|��;���Ǵ��pҚE�1?���֞�RhI�֠X����?_Mu�$
��&+��*MuK
�}
N�|�^��:��I�q/RMTg�0c�wvO��Q\���~~���)��SM~��)�F�b~P[�y
ETc���FRr���K�������&�b%���S�����LP�ĀVF�iM?Ęn��p�#LcGO�\��A��Β�N���OPB��0��<bk)~��
�O����H��C"/�8�
V
��.��='Ck�ϰ�q��%^^�_h�3_���#_,�����i�%��i8��2S�!�G�ĺ�����j���H�;.�Ř�{Tۜ�@�3ɇAw�W�%�ܮ�qƟ0��@�JZ8,�U e���v��2�2=Ԟ�L�~r���sWV�v*o�k��"�� *驲2o�u�u|�MO��Y��H񔜿�wF�hWL���B[�$9<UCJk�w֯�l�Aw4��sX\�z'���]Z{vٍ͖�c�����=�S0�J\�r�xŵ�Ij��!�F����,�;�l9�q"c���ׂ3���btF���q��ɭ��T�ݙN�����K����y�k�dX���k�Ab�5����'��������F�! H�x
���LEi��dE3��B�㓴7��m10��
�ճ ��C�qiB��j�2�؞�]��NP\i�W�fzK/�j�dm��W���Y.S2�
��DQ�B_]s!�N�sI���r�(�-k��K� ��.�a�v@p�O�/�=l�,� ���*���r>6V�`U�Ǖmhjxg�g���&(�'73�u���Ys�f�@)�J9�ڡ�f�{@�Cp.e$txK�c�����{�H ~�S�3U�S��"N��3ަ���g%6l�:D\��$����~_�0�A�jI\�_�w����ƅ��B��i6�0~��_���;�
�bE4{k^
4�;��D&��R2����iW��L�{�j+`f5�i�Є�b���%�Z�L��&9g�d��Ob壵/z�Nl�?��D�A��۲D@e�f{"��������j%�aU;\��)��PK�0J-I��'C�:%Ħ�������-��W#���D<�3��7����>m"��2���F=��w�~&t�]�ɹ�Y+h���b;u����r�h��BȽ��4T�
b�;h�&x�~N�Ed�f␒�^䀗����4=��3d�(_���9�{��I<`l�.󭯴Z�8`�{�t���F�Xph}g'G8�[3F��O�p(F����+�'�
&Pi9U�W�o=��J���x�D�� ���)vT ��=B� w�*�:h8�7g]u5����5�xuG�dHUX����j;|o��:�Ϭ��~�����R���$�6��.��#��0�Ȇ
5UV��Q#�����dq�AA����l��y�t�'�[uס*���,zo��xb�q��JÐ���Y�����K����"���T�NFQ�P� :��B�a�鼄��L��yŽ5u�/��ۇA��lud����u���kZ-���-'*  ��K: K���pœi��j���V�jk�'���0����=`����Op(�ME��4О�:ѾMrl��>���[~�=U����"Cl͆���u�,�n��C��B�ǵ�b<"�}zu3h�(��Μ4	➈߈x�O���̗��I���}�!���8k&�Sh������I��s�4
�1t'nM��S�X�m��-���� go	�Jޘ� �Eҗ�g��s�c�t� ����f0�O^���q�X�0�Q�{
��ʜ�D#c�]g������J�߰�i7����ݤ��a/���n�f���Iz�b�X(U��W��f�8��~@��R���#�E����H~�]����AJC׸VT_� eP/&XjB���n<��!nr�jx��J���v������ac�KD�e�-%VB��x���(}k([> H��i��	xz<�F`�^s�_d�|&q]Xl`y��$h��s�CG*Xxe���x�-���.�>���O��i�Q^@V��y�B�t�r�峩�W�L�������&�R�b[A���M��3���m��]��r<�f��=Ve�a��.5