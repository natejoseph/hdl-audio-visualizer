��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�@�{�ʩ���.�l�e�ir��Rjnג��V8���Ჯ����EQ�ى86�����8��_ғ&��.�L̇�#@27F1V������i8�,o)��ɦZ��_(".v�9(l��&fO,Z����Uof�~|�M��ߎ���i�HoCїp#�u�_bN���́K�i�Z�T���}��r/o"�Z��7��M��U��2��n[�i!N���V!�Ic���������|'A�@x��R'#������V��K}�T�P�Z�M\=^m���c�|WU��,1���j�Y��U�\���M�}�9�buC�q���Ko���Z���%������a��� 2�T@	=���=��d���K����@tsts�����}����q���QZ�j ���{�˻�[�F`��?\OF���X����S-ڟ�O�z�D�.'��gTB���̦^"���Sa-3�"9Ki�r���Yu���q\�����r}�$uM�� 󉍕��u�L1��;���m�I$Sz��>�g���i�޻�P�%��0\J�f�"<�

�As �./����*���v�-�%�%��g�98֗ͣ\*�G��Z2JlNt[P�)Q��c�DS.)I֘��u_P6��. �l�`n`c�����C�'4�2�.���_�4�y�_�A-~�ǘ�}`���BO���U�<�;��frRc�N��҄vX��4Q��r�k��v��Oo�ɟD��:H`p����A0���T�[�v��5~XOT���3� ���V��Bwͣ� ���֝�"��8����Ƭ�;u��Y_�`��S�^aHrsMZ++;�0n&�n���&��z��O��U'�T6eo���ҫ밪�<}*�)1��&Da��hw�d�K�`2�iA�8$ى�����ɴ����T�Z�0+��aDX�W����-����^1D���e�3\�;Ŗ}���QR�a5�M���ړi蛰�	0q�'����Ya�5�WPۦT�$U ��+ŝP<�H ���Q+6����a^�-�r��G�O��A��d
�h�I���7l	���݊Wz0\��Q�X׾~��ď$~�r��9�2��(2��[O%؂�f<� Eg�=6�Lt}�s���#7M?!a��[���a	i��}����H������8��łw�PK��{�C�%38�i�����<�x��5q|6o)�X�fr�{ܡ0М>g�|ţ��^��2S��-yv�qw^s.�&����V~�����L�Z�&I�zvJ�:fbb.T��(n#:�TGz�M8�N���m���d����r�t+zʞ�ȷ&����=���,(+�0w�0U|0��S�)c	 �B��������I%�� � ��^�l:تK��ğ`�L��'tK<�Q˗%Efhac/\�Zm&�,��%]�s���R������]�i�����)(Y��Y�2e3�S'r���?Q�L� 4���X���z0.�ָ��/���ș�Bܣu�����ӿ�e� �2	0|�봳�0â]a�Qb�hm�R}�~&�V�x��]�ؙ)��,s�x�)�(�n���V�~v|��v)SH�Z]2P�9}�]�ɐ����0�4���,��q����De��ԂX��(3��+��
ё��`��@G&����u�-���9W2�d��W��c�(تi΂<�a��W�(�@�J��G�L�~��ͽ[�����LZv�& �J�?ub[��i��Կ,Y�\=`�,��}�b�Y
:Tb��:�I�s�=��|AM)��֭X��ļ�X��vb{�4�7��j��Y}��za��7SWpY�.�fl�߷܊�BL�p� ������I8ߴ�)��s��ѧ��^����)��f9�O�C��(�Xq�I���Tڒr<̛��W$�>��U6�;��oO�B��ذZ�y�;���9-ʅfc
Or�a*�5�H���4�۾��Yba�2��^��޽/�E��6*�P|i�`d,�Ѻ-=VO��"йO����,;��op����)c���l� l�K���wk>�.S�2���>8~\|x�Bjb����6<�跭�s�&���eU�vC��Ƅ��1�]�8�J�K��ym�805�
�{Ds�&���5�5`�����9���D��k`;C���`�,�SH-�ޝ�)�4LI{b���#F�fKp���'3�T3Ea)b�[V�r�����b��s�e+ũQXUY5�k�]��*k��j��82�y6 �f��4�9�o+E�yEG:��H
�~ռ��Fl`!���ZD�Ҫe ���h$*���)������<���
鎯̵m��J�M�b�8�yA��{*�5�wv�c;�������ef^a(A�7�/(<����v��-��%}��ٓw��6 }�% �_�\	R�'�<C$�����:�9h�-cW;��G�J��>8:� #a��/��iά*r����`F�Y��.$P���׺"�)6�}E�=c����ˤV�R1��m�[>�� .��E7��W�,2^�vdsh��R��}��*{]���0�k��t����]^�:�k���IP�M��t`8�_"��"E�>9��vX��5�����S3�]\�-}�I�Mu9\'�#*\z:�}t2�-3D���Q9:S_ey�sax�~,�I
�M�Xx�р���Ĝ�׃mVع�����DEc%�������>>}�]���i���TW���徒LG45"�ڧf�lc�N"�ذ�r�csFm���0��0�1��V�%ʽ�R�����'����dm_چ:;�yv[V�1a4}��q�ZUoZm�m���[�f���t�y�z�Y��N�.�Ð��{>������r�(�(iG~�۶�2�����0��U@��[�s~B�G�;��'e�
�M�G;��;� s*�\���1VK}
nZ?��S�.����b;I���|��|ʃ ��z𻓷��=��*���d��y+��6j��@}CN�z?�'m��u�Yd���ɫ�1ѺD���)=��x�(��:-pAj{�xEu[��U'0��	
TZJ �]��ɦ���4�(J��pR�}����E�g
�6��IP�th��v5l�(���t}ݩ����rF{�W�\�@�[�.>�38<�d���U�� ����u�V��%Yg���m�L%B�����d[�Pc�5p���To�e�e���t�j�u#�6a�0��P�	�yW
-���ZOvo$�򄐀H��AU�]������d�	w���qZ2UB:���&�N�\R�ҽΟX�r�v�O��r�iR��<��Gu�i"R!��)Ẍ��M<o�m�����y¢�"�)�_������ᛩG�������jQ@1m��r�#�����w����w�^�k�xP�%FMz�lm�6�B�v^|�M�j2&�ejK�
^FY���ē����&\��B4/��Ԝ=K��\�~l������̈́]=�OO��S��ʌ\M	̅޹��&� ��Gd�/�X�Ý9��8M�ٌ�gTG��Oك��,�̓��8��ױ�^�l[M�cJ���t����G�_��ɔ��+������ɕ/V��l��Հ��q:���e��`�U�e�PʚcLb���f/Au5�F3!�����w"N*��)KǺ6���5h���K�3���~���\=oS��@�J���u ��۞@0�g�&B��I�_ ��������l�;�B�`N��vY,  �Iս�dV�]E�.8̺x��*KY">M�OvcL�����TaTC>�'0m��$���d�MnYt�&�0/�������h�
뵣n����~t�iR}��l,�nt�����̂��H��A:��e�A�d�|��A�S�*rm��I��1��N�Z��5@}!t���䀌��Y�d�����M(L���|,��aIA�b|9k�9~7�s`]�Ǒ>+O�?~U�{���!���{c���������f]�@yT��&�:�c?�s`^�gež�ʨܑ�������t��BQ��,F�͛^:S�81n QF`�n[�"�q�?��8�}�:�EَViQ�O���k��N{j�i��[N����HS�-�/��pu�V���<9�]>����#�䯬��ȇ�ލ�$ztw����ØUۻI\ے]�Ք�1�u�����?#S�R�~���Yȏ��TՎ��w�*H���+�|���~]��U�S����&�Ⲹ��v7-
A�+7�tTkc��H�U��V��~+��4Qw�k`x��-E?�I7�������͖�͊F.��.����7��0��o�]�>��D�X�f����Q���A,��Q��6D �4�L/��m-M?��1���p	��#�2�~�Y0�e��s��R�p��X�2��,,c����1G�b�g`�l8�����+���M��h�7ٮgI4�$!c�;-�]İ���|�?3��\3-�����mVq�Q�M�EF���#�V�>Wc��@d�,|�H����_�<Cr�г�sB�fR,#"D~A�$9�g�%v�% ���n����h�Y
(�2ł24�=���$q1C抪��vp=�z�u�?��\��Ǵ蚔�>n0���ܨ��P溲]���+;�C�iV����Z/9�@�c΂t(��<Rt\�8$G|�̴>�K��7FR����1�j�e�cU�5�Ɗ�OB�4�ܜ���SGș5���zP^���_�|Hqs�V�yQKG������d�w��.=��n��Ϩ�� ��D+j-bR��01���,���6Qz���KzfW�<]�:�#��h&x�>�/�=-<��bLM�c0y���lq�z��Q��Cb`&]�$�9*3�ɵk���M���F��y����3T0�ҡ(U����*����w��{*9_ �i쬚��#]r�&�@Ǎ�=����,7Hߴ8�R
;�����</n4ڶk�@�h)��[���x���P�d �	}�m��'B�*B���n��^�c��}?'��20����I9�J?#!"�4�-�d\1Zfx�$53	��q[﷐� "�N\��������бڼ~>��2�"��Ꮠ���Ѿd��L�&�V�[�~�0ڕ�-�oJD��'bq�S��u�y�ƹ �ܜBm���3\iYcB�B�bD�����P�н��1���,��jĮ\���������z��� �sX��I��sgR����f1�ISf���)�nF��@W=HZ���{2���L梪��+�i+eՔLy¤�~-�6��|zC��f��G���n�Q4�~^������~�Y�E����뾺���lH�j4fm�x��	˾z����`�"�X�(��Z�W�1Ѐ8y$���!I��в���ثn�������A���ϓ�����9��ޛ�+Dp}"�`'*�ä��f���є���w�
�,��,�h-0�hW[[yR��������4"�������'ڮc�}������ˇ~u��Hj.�<̃�ܙ�õ$�{��^ro,d
��B��ll�>ުl-=���хI��,:A��l��D%E�D����g�qZ�&g�؎"�7Ͷ���Q�ȯW�v�@��d$6�+�?Kn�x&m!�k�A}�ga�c�`��y�8��J� �1	�6�� �/�N���u�����+��ݴh��/z�j,�XD�2�o�cX:�+&��7$j�ԫm?q�y˄�4�Cu����}��Uվ��$��8�u���a��x!�O$��<� z�8����؅�=&-�����O�@t����KP������jٻݪJM��/J6͢Ԧ���X�D�͒�d�Uı9�o�Gg� ��F�e�"п�N��v��n\�E��)�LC��QX���3|�˫�	?�r��>Ed�s����]`�\ezH�꼏!�#��
3��_��� �r�[.�o{�y������HnG���(Fv���{T�oW��<��,s���V��vWY�
3	���k ��q��y���R�V�_�2�ǖ���no�m ��ק.�G��Sy��c:S�՘���BP���E�3�~#��gߦa��)��C)��i��T-+�i,R� �y��˺Ư�O�oH��e��5���- N�ֈT&��m�s�#}������pO�P�n������9~���D���D	%qS�/(c��z��߂�"�sp@�5����xc���[Фd<�q�8�R'������i��|���5{�����{R����]���#A��<u6n���O|����D=O$Q?��3IJ�j��f *9���� K'���l�ƭ�P;Lҳ�r��@��V�R�Gy�����D��Ț+���Q�i��΃�pb�/����/������ ޏ�=�5��M��q\�גe��S��lնW�m�;Ҡ�H�>Zr��i�3^�sw�l�p����/�󷼦o&^aw8{ !�r�t���z�hᓱ��˹zr��@ɧ�2J�ڼ�zŦ�+/x���+� e���{�r�`�������7	�sg?jF�d��>�����I�׀�xS_�ږ�jk�K��d�A+�D��lT�F�]������v��u5^?J��{9u�	D�2��:v�q�+h�[��ܶ�u����6�Fjdba�6J���m&N�21���ݰ{BL��g��Y��Y]�p�7}�]���	��n��s�.ߦ�dTl�($��@���gD��[Q�/4(���p$/tk� $�T�g9��H���H>�Z9;�FV(�[6y�����{����Σ:�W{JZ:�o柬�H`%76W�֛��) �7}���y�}\y�)-�P1�e�;�#�-�Ѩ�)����Q�N�sDة}���O�d�2o�M��뽨;�2��Gmž]7T��N=[0�0}�V���9:ۄ��>\+����&��ͱ��!�Ԣc,~Q$�CW��gZ�K��i�uC��'as���7%j� NM���
��%S�T7{�����nn�ʽ��_K���?�L�?e��#C�Y�t��L�]'�)o�w�N���	M���뙧۟��L������+�g�2+��eJ��7��~����d�e��]d%]={SO	�Q&d{�;u��(��z�����&�!��ħޫA��/���x3,��R蟛��*>�0o	XD�w�r [[�k1�ك�p�C}L5x�
��m�#�3 ���"��D�h 㽓K1��E�-�R=?�����kJ�z�5(���i�
��	��p����J�րܕ�� �H{�"�B녆��aݰ;��0���y��A>���4�Z���l[�,R(o�x�IDpER\��b���FK����ġ�L���ZF�ywV�|�͢���9� ���yUor.�!�C�CH�m����E �D@:�2_i/2���f+��}����?+n���j��n � �f^���ViV�4Q�6,���lә���"��E��I�	��?�3����f�SE��1%�z�_H�Ez��}�Aa�A��ʰ��o¡9�|{�A�du�R_U�W]۱5ߠ�욪�v��s�a�J/,�3k��R�!ت7s7���?��O��4��t٪�;wc��:H��̀`�bu~�Ő5^���6�K �s����#�+uR1A��)b����hÏ�n&!XO������n�?!:��#]�}����5����n�[.�8E�.����9U%N�X�����w-!I�mV�ԟ�Fw��.Y�4N�/��(��LVXƵYC�ubF��V~�Y���+ľ���&�@�����^��~x�ȵ��a��HM�k�~��X��'I���v	�Ҿ3��:�d�K�U����d".8c��MI�a���G��#���M��B��$���K|&�
(t㛀pSԁN�6�ם�柂���)�����@gk|�be2y��˼�\*����핤.�
 :l$J����6��!c�d��^S��P��թ76Q��xxA��m�S�K���, ,����,fu��Ӭ1��)�Z��=e���٪�" s�,�COqJ�����YL��������w>puw/ ��$��jP�ai��(ɗ��[0�Q��h%ەa)�+�頦17V6<���Fr~���=N'�!�d�Y��v�W?o.a1c>��?-r
��<
z��{��#�  Zi��e2�vU('�Fi�t\�Eu-E趤��Q�� ��f�:MY��N��N����W����?����LQ�	�}�)Ô ��[O� �X��$�?g���� �~r
U��x�WMu�%�,��2v��i�s��Y#����lˢ�E4(ڏU�����DWܑ���.���k	üPB3���9�Ѧ�+Eq�{��cv�ZQ} �v|Uߨ��������	�bl�C��\ "��3n�^uJA�����{η � *v������@���`	���K�'�7�S2닒R�.������gb �6ISʕ�&���b�#�[��<�o:*��0q��Y,X���Bv��@}��կ=O�j�ރ�z5qa��19S����>I=�S��0����ڠ*��󋷕�N��@�4ZM�K�a��2�C�L�_0�L(�<"�.`b��x.�{Z5�7x�8�UX�tX�J/�F�B�//n�%���N��� ��V������@]�u%�br�Y!Ƹ�lD��<�{������p،/����v�*�� m�W�R�
�0��E/s�ʮ Ї0z�_�Z2�p�y���2N����$*=T��{P0��z���>�5�V:��������>(���Th%��Vr� ���:��X�{�|%�У���Z	�,�9u1��m�\�0��l�%�#a ��s1�>�!����Bap����-�!�n��;]U͏C�n��F�LS!�*��U0X_tFF�N�w����&$0|0�ݗ�y�S[ƕ/�4%-w������s�U:��	��k��y O��fk$��C͓i���،�\��%�w�EW>"�&��ϡ>d������X����4�]�E�Ե�$q*9�^����4�Nk6��Y���>��m�b�'�U��8�]���ʎ���t�t%�bW#�Irj+{M׬���j`����Z
Ɖ�7Y�)�.X�h����W�o�V���Ts�x�]K+f�׵��W!SL�,֘�*������/Fr�cPA����
���	������q�E���JAa�W'�Ua�#����4{o�������rL����2��)^����a�v��}]��9j����([�ն�M�����#$�yh9�^�zC�?��)Щ�@�-�l&�P�>�)�-�.�I}�#�0a~ב��
��J��LH����[���*�����=�J���c��a��z��s~��ґ��򬖔���)�N"�=-7D�rTF��5��m��h �ӳ*ޅH!������{�
��d��t�f��t�
>}���c�MJ�CI���cV�o�d�l�����{E���M����|p��;��|Q�Iul�I����DC����{7��e�!���@`G"��V�wI��v����2��֚?�up���2~�������t�Z��0�fDC��VhT>Q�%��0I�Fx�rIܢi�'6}��E�8��^�_5�V`��\c�b��M��h��<���Mt<��T{s�L\-�� a�Ҟ�at��Zq-BW4=Ԏ�x�,"�T�.�wN��v̐j�D{6TR��r8]p.�P��JM%@�J�����\�ƲK��\��r�|c�U5�R����ϣ�v����8ym�X�p��A6��oA��Nx��BZ�F���CJ���4�&?��5EݭȈ�Z���G� �:*P��Rܽ�;Ϲ��z1'��� �!�-�=/�E��e��d��v�m#a�_��J�i#�v/�������ָ���k���/����a�ՀMB4��;\���%1;��i�G޲������ԯ.�a�g4��*S�uW�K��ە����3��2+b���^Ar_KB8"�L?/s�<j��z���&�@a���f�!��7C/���G�{�$^A�5� Ԅ�]!˛�
�gj�u�w�.V��dy��#l}	Ñ��:��tQ�I�)Yr��<R]������.�}5���G�����Na%�"ic�׵�F���i�?.|�ֻ�慷b5ݰ�P���p����F�������@E��cID>[�u�`."�GoV!֕u��=�N�Y �Q�N4N�|�@�D��o�F��p�F���/
�U0^i=o ��9h��E�������y�	U��G$U�-PHX��.�W�4�[+^-h�� )_+$�WІG�"ߋ�^�k�d�h6Suh�ά�4��Ej���T�ːl���"��,���K=/Nk&B�7��V͞iRz�L�j)�I;!)�!2)~�i�$fcR?�QZ����#A�|b�|8$�`\�������D܋e}؟�2>�i�51�1�]2K1�{Z�ܟ�wU�o���J.�%AUSL���ZU�+�T#imJ�B�|2�d����)Fd�O ��T�,_��"
ao?������b���;��NX&��g����u�<� �sQ;zU����SE��ą6=���h����ڲ�7Qy��K���Vo���o��>�`�}��9͜Ru�
V�~sY]}�au�ρ���$�l��'�˂=-L�آ=a����	�OO��;��X�f!����\��Z4�`{�\uo �w���4�3�,�3�N��G�䄙��"��$�ْ�׉�<y��R��4؟��%�����)�	��2�2�f�.W�(������_"���_�m�Yw+*�R��Z���R�~�J�q�xW��+�+}�g��E ���ǒ3�8�a�#�r2HBP�������$Βְ�<�(5�]@	��|�}bYq�͔�E�
7��/W���ꁉ�W�Ѕ1��O$`p_Mqo�b"��f Ai�|�t��[�ڶ�d�wS��8��c�~!`�B��;�x��O�ho�dせ�m�S��PhȤ�!��LgS�k��
�-q�(��wk���_�l��v��o��2D��*��H�|��<ud_׸4�W�u9��g�i�7k��r~��r��"� /䔎�	�]�o�~��s���gW�w�`A�VT���_����"�hT���|��=�毚?T�iX�U��b�C/#���I7��b7��:Yuk�q�}ǽ`�c��1����d�P�A�@�Td1!FZ&���Z)>��aI�I����R"�4�aKx�   �h���K�� �n�v#���a��4�ᙼ=&LU����`u�AM��q����(�� �D�qh6ĕ^}Q�)#�y��������;�Mm�(΍�S2�P.,�2]�8q�й�\hxp#���,�!5��a�����K�\�"`����z_I>b�Q}�g%2�Y�)�~��z4|���-�z�����N���C2p�q�/Oy9���=� K�!3S*k�Pa"�;�<�&̗����K�G٠c!<���AX�����!����
�&����N'�.gڼO�-uIKhT� �櫧��Q�j���T��0h����-2����R�(z{my@M�m{⢙8��:"��������1,��ܙ�
;��ں*�y3�"���Ŭ�ְy~g��]��[ ��y�@n}�sc��۝�DC��xSq������5������[5�Dz7�C*��př����{�3Fz��2R�ukQF �sޓ<�`(�Zt�L�,dJ.r���=�c}�W��kй��G!��]��ӽ��s�%�Aa� RX�G"����f���|�7�f� �>�;d2/	G�Y(R�凴Z  ���d��+>��2x�ٴ LYΝ�:B��˸.�A	e�����?�����D�J��������7t�n+�ðs0�]�yaE<$s��
?�
Xd�#l!���e�⨆�/�֡	?1<��c�!��jf����-��55��a�=�D�Yȫ�c=�Ԃ|�����,?�*�;"
�xόo�c>	G������w�9� �1j$�!��1+b#��}aX���������nn���L�@j���JO���g�dO��.�YrX����	�H����X4��]���']��/���F���w�{d���uZB�8����c��*@�b�W��@2W
o�ϻF��%n6�m��3K5�-O,�D��>ĺr��m��=79Oᔯ}�0�B1�����C�|�^l��t��#(㡐yok[$��@$�	+Q+���q�F�t�W�׈��V����-��ұ������5\A�j��}��h��������~�dH�f~�!d�����[*�{Qש���c�!�u��C�N�i;�	�Da��l� ����)����|B	�-�{�Mz������j�%3��g,�"�/�:��s䨠,��GDi��dkj�%Y�*�M�scic�}T�Dd2��KFs�zM��V�ʸ�";?ɇdCB�י��Sԟ(աe��l��4���b�3,��S-Vؼ� Z|LS��G�KM����"��ND,�<��ev$K�6��yi�:�� ���4���4X1tz�!�����1�b�@>t��]�Ŭs���p�m��-��x��x�"�|�0M�5�;O/�Pv�3p�����o�I�%4���1� ��~���1;R��vz��G���������7qَ���$���X��ġg�v	��JM��
^�
O+���
r��&�e����$a���~a|qi���С[�`ˣb�,N��:���C�p����VT�`D"
>XЧR�9��x��R'�]�[[�E�¸s���˩`M�5C�Is��~427�`�{�H�N�i��k�{%�6mJ�.�3���J���2c�c���O��YHe����v�;�M>t��w�lQ���v�pĈ
��Qwo
D�T+c����R�kk�0��Z�n�%>� ��D�0J�w�.˭�¯f2����e���ƣY}�(�����f�ɬ�\p�32�;	��S�F�'���Ϣ��@0��u��u�U��t�
�a��L}�D�b�^���R��v@N��tvz���iTn�Z��>��}�W��\�c<�j奷�)��%r�x^�
(^=Dz-�8�#��λ
��Q.�nm�Ro��a�?��fm,����z3���j!�|zS��(�J6����^Ej[j��j����
;��>5�A]�"�i�F�Tf�HYfE}d�8�CZ�T*�4���85B �#Ii*�D�F�){ٷ�@1IUܵ�$���W�`���C�՛!�����qn�"�h�ۈ��GF���[����ڳ/�iG/,��4�x?��z�6D�M��ɅI��Uq!�c���f�������� �NE$�zF�כ[ŀ�][��=�b��\k��ĳ�s4	�f�=±�D���)Þ�;rɵ��E�����ă��W+hO���V�$ӳ�ⶻ�r~�;��vЅ�$�0�J�ä��,�2����%R�6�%�;���ڌ�(�DQ��A~a�݂�������(�P^�2���7�F�d�P�Z�dwlįH
V�	V�˄D\V�=.��@U�씔%�m�`�d���>8�l ��>����Vοs6�V�.k�	8�Ա�
(��:CK)�̯����ᵙ:���:�1 �U�x��;p��������8#Ӛ2�~Jg0����s�}#+-:����/���M�gw9�d�Q*4]��`�j��}�;�f��7�&��q`�ꄂ���ɉ:�V\�˧{����Qg�?�9_Y�N�(���{?uƿ�s.O8�=�5�����M�EӘ�l�өS�zCƵ�`V��pi��[=OJD�h���|3�L��>b3*��D�T�;Ǽzk4���|�;�O�$5 2|��������A�.Ъ]>mQά�N�OR�� !Z��+M�@qz<1�F����5	�l��?|0c_��:�o�t��¯���X�h�i��4NW!H���a����9>C󥚳���֏������u(tҩԙt��k�?+����߰�SY!~���Ot��i������x�����p�*�ڸ�G#�x۵J���f� ��!������3��(hTw{���쫂�'�D�m@�Ɏ�n��\`P��xO�}�2�"!���U3J��ӑP��_�$��z�R�&�A!�arhqҋIุ%v���[Y�6���ݴo�3�I�Cy]�d�e��|r&	a���&���A�nub�鐶��b��W�e� k�rZS�^�rN��L��u��[�%6����m����'��̚R��$��E&*�F
�nM������^"��v�@�e �hV"x�B�+ߣ����<&fr�b���3����v&�`�n�㼨���$�@��Y��?�l�r���i!��G?�B ��+��
,\ ��PwSD�'v��+�xE�c�W�~>v�Y���+.�?6��oB6}��cy{�����R���3�+:4-��K,e���j�k�i�L2�Dȿ$^�5��5�����t9��������1�9��GVR�b�� �����m/+I�^�t��f4�7�<�Q�A��ӭ��2{m�����/�I��������x���x�u�S ��<�v�W;o`F9E)���<%�N5��F���
��v�։��˙b���)�"��:|��{����֫A�x�׌є�R�S\:ɸI32�*
T�ፃ��I,�8����#����D�����}B�,�x��B^4�V�֑�����8%L:l;h�w+A�BK��|��z8��ଗ�爈%�� 7k�7z��4Zց3qL������0q��y��B��W�]I��LG�,����x��p^����l{�P)���M� ��A7��ˮ/7�����+���;��ܒ�4�cL+t�����Z�De���8&��L���=�k�����\Q��,�[k�hsLB�:�)#V���P~Q"��Oٵ��� ����]����� L��_
1�o�]#,>���R�v�R.1s��~�����}�SF�~:���}�
5pʂ�1�:�^YIg���SR&�'��v�Ѝ���M0@KD�hZf��ehZ>o�3I��.}�o�ǓL�ka�:]]3��8^�&x,������lB�S���k�~��D�`c0B� �ueL>/� �M��Ց��)������2l��g[��D�����T�"*֌Ԅ���ļ�do7�W�pH�����°���.������=\#xs�Bz��^YWB
�i�v�}��J؀����{�S� X\,�J�,�O��J8���ß̮.�ՔE���Oҋ���B���!{v*�!ۼH�S�J���:O����-�_%Iƍû�M���*�)#Bt1����x��DU*n�y�m�
�x4a�+:`��q�<0�����%�}��%�d1yq�[�Tl�!O��O�q��ks�0��I�mA��cYt}�����,Gk'ȟ�G��S��K����2H;�������!�uJ��l�-�����V)&�R�`a�/ PI����U��r��#U�s�Y� Ƈ4��#���ì��݊�B@�+�:G�>�M|Ah\�Z�\�{��,���E{��ɀ��h쓜*�w��2�M��_k��?��x}"G=M��G?�����;4���h(E�ZդO���h�?[�����	0��G�$�v�N�ύa���5�o,�'y�6�ҥjeR����А�~w	��T���T}'k԰r��'�`�c�e�^8I@2y�%I�K�p�;�7�c�/��f&+V{yeO��ݯ7Ȋ<�X�-��Qp8�)�eD]Ö��JD�{�d�$!.�ĳWmqg1J�