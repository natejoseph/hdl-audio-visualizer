��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O����Q��VT$��~��(��p�`�i&��ҵ:F�����M��[�͔��g�׬�퐕��}:�p�C!�,�����D0d���{:EAA��z���^4��)�?k\���g���ydB��n��N�@���-��>�i�	����e�fc/9O6Y��W5������z8���9F�������)"�?ؽs��wʂ»!Χ�=vj�2��:��:u�U�Br�-��T���m%䇨LM�����9��Vn;�L�]��|����i;ж��lK�����z,�.�+�Ā�/%u[i`�o���H�D��6�`1��"�$}R�SM���/my@^�8����Wi�H���.)�m=�/D������)��e�:�����0��`~#V�R�B�~�?�>�Ir�k�Cy����"�$}�l�M���w���$����2_�xC�����׺Q��Ў,r�J�e���)��7]�f8�yɸ������_�O�c�F�b4jE�9`ք5q���8���豘�c{3X��7���w��[��V,������?�ӧ �>�j��n�����k��͐z�\��'����c�͔{u2H�ߗbJG�!tB_�e�c5�.��L^8�wEb��.�C�՛�Rc�7����23��S���,�Pg�/���:2��z�n'�j&k(ה�<ŕ+IpRgAj\��&�@Q&�n�N����4��pH��O�����FE�Y�}���O����
U"����wR}}����sA�Yn�`f��	�`��$e�0w��!�`F���	�pa������=�Ǔ���;� �G �^�X���{��۴�e8�Me��7毓m_f�;���ְ&zS�ņf��Ѷ�"���Q�	�_��8�	OO8YJ�5|��߬g)�������>�����2m���~��?��������H$�8Z]�M�=_��D�c<-i��&Eh��?�]Ѵ(�"V7ED���X��!���5��M%�_�,��>A��]~�����R��+���B�@�`�^E�Q�6������8��,54�~C��1��d�R�����7����#�H]�8�EK�R�JG�e�,���e齽����e_ɴ}�>6R4�z���͔R�<ܤ�MS� <��P���D�>�'R�rw���e�f�j�9� pV�ۖ��}��I�qЬ+�\My^m8۠(����OHs���.p,L��?a�#�v����?.��-����8��O��w9�EM�'�6v�GGX��4+-�V/$>� 8"��у`�0�#A�?%��[����S�������d例���BR#.�B6�G��"�$�Ӝ����b0����K�1�D����-[>����إ.!�HO�M]:e
��}���26t�/iIP�Z6Ѓ�� �N=�@����_��_��*fJ��O*�� .�E��LP�Xz���9 ��;-m��X��\�������}���ߤ�heh#�h��g0H�.��B[�Nᚩ@�@��p���t�_�4�U~�j�7�Av�,����}F��L��0'n%���A5X]c�P��(f^��D&d''�?5!Ab~�'	��:��Tl�'���~��,l���YM>3�8F8t�D�^i�Cv �3�Ĉ��o���_X4F%�af�x�m0�K�c����9���|ˁ�
9��ȾG*n:��R#Ì�b�+����8"�8���B�v8k��Qe�Po'䉅w�+͚��cgn,q�˯ku�t�M�˹�i�F����q�E��S㙑��v����HÓ楘��7˨
!��5w`�3�Z��lZ��~��^l��)n"���*�5���,zr�--9�[)�x=2��&ҝp߫��6����Щ`�H���8J�p'{��ћ�ÌR�Ύ�����7��5�K��S��M� �l��E���=b����s�����~������Xv�j��rI#SǢ��f7���W1��#S��N~�<�NR-~�������a�iu>�5X�U.�
���C���y}��:�kz@�:�	���vaG��؂�]��%d�¯�D��x���B7�q}��8E�Mn?n]����X*\���� �|�=�	��{�O��w�O�e�p]�����h�ϣ�?bS<�"2]������s���X�$�^7.�B�� ��j{�7���Ց둩FG������=�~�a�������uJ�c��s���Nṏ�����S�d��SX�l�F.%��Z}8� ��ҘO�<�joĪ� j�*���AB�U�-���AH��V��1��,Aq�79[�bШ�v�H0فV��,����{�!�?��^������ox6R����~|"@��<a@���E�����e�F��$�����_��>��L�mmΓ�֫u�`蟟+�&o+�/d���n�J�pViM�F����/�2�����,]�)P��*��7!!�B�n�? ��Q;5�~�7~x�˳L���N��E��z"ᣵ'd�\*���v�vm�	���)N��C:�u�#y�ǆ�a�rp[��E��u����ʩܧ�[n?ܾ4���9ӂ�^��X�2�$�8:�R��ä�.t|%0���@�w1�_��=^V|���UNoL��l���Ժ��x�_Z��G���׫ <���E�< �V�&{�p�ׯE]5y~$Z��W��2��&5���R�g�@;}�Ҍ�V�~�dY'W�a<u�|g���X��Y*���z��F�b
+̤�<��nn�SȃL+�G*���}�q@��ҡ��G�Y.���k���}�i�)�N�W���vp�We�l��Z������P#��nE$��O@��������y˥�!��B�����w������5�;�x��,��ކc�onS��"r�{��ib�`��������ӌ�fz+�$��*�~�Yc��??����
�J�=W��?��7w��w�cþX!���[�� �p�]4�	�BȤY������z�?�V=��:TR#α��!w��D��(9��񅢌�Ч'�E�+�l�u{�������S4V^���:X6F��#�Q��x�h��`�\���}7cCc��3k<,�K4��T%��n������zXc�i:�"֪P�Qߏ�2LN?E��;	��;#���n!�M(ɆX�hn�pp���@�������U�0�w�x��QP�P����4#�P����t0)	��g�N�٭�����w���_H|.�G�m�l�h�N+_lDʍ��*(���<jlWa	�h�_��%��Ce�l1eX��oC}���2��5�C/uF%i��8��~���	i*�(�Q�KY��,��}K�xw�h0VR�s?�f���`��_qrq�!>��gv��ȢU�Qh${q�%a�5�L��r��������c���,�5[���E��@FԬ;Qm��I����O��/8t�Z�:o	�N�Ad&
~[�x�`;�����H�G1V�Q+���-�mK�K
�<����Gql�)u���ą�!w֭�[5�hf4>5�����wI�sc.H��Z@��AİW&W�[���#��U,�_�#o�M(?�>�'��V�ِ짪|�8`���o�>*ƆF���}L��l��q`D���F�� ?���{�+|r�!��3��v&rп�4��\�8�$Z�Jc�2��A�QZi��7�����Tޝ�ب�&tDq���v�?x~�;�)Z%�v9^h*���o
�h���+WL+����u�D�EGC��(>N�	+ r���ϡ6���lXY�}q��<�nOU1f��I��69,�d>0��b� A^-��[r�ظÈb�)�D�������3E־�4�܀�*�O3|��Mk]+��-(�6Y�oϘ�:΂< '�:a7=A:�.�m�u.����mP�K�.d�'pIƑ��_Op�5��d��+t'�ے�7�d�A�1=D"E�O�ϱ>�?��K
(�x7��m]��pKY���F�����p�O/�T�ąQՙ��g�uw-R]���?�L:��E�c縊;�T;�
1FY�W��[ �Z����[9N5xQ�_�q8�Y*J)[�׼�᪁<�6�=Z��3� q�k��Ȝj���_�Q`G��wBv�L�r��N�����(&Vj�p�^�O-Ț\����I�Ïu��r��1������������$���(�o���^�_��e��Yg����9�����Fv\�!!�+�&g�e.s�r�5��r�ȓɅ e&��4Lm̾��7nقT��dQ�V��P�A�ʵ/�qV-&8�l@zT66E�ni�d?Ш=�����~���o4�>�o�A���dc�؝7�?�|M��V�4�u9���#.qә}�-�����[�N�����p.`������ǭ�B�K���j�1-.|'w UV�>�dNp	�W �Ŀ��4�A??�޿)4QR�&bñ�Z�&:g}P�:@�>y��w��m�/�'A6���Wv^�g��Ц����R��`��>���fC���'��uy,9�y�$���ʯL����]�~�,�d�dҖ��Y��SL@K�]��A��3|�g"%#���j=�-BW���Z�q[s��ЄeG�U�:	R��.fd���P�YK}�V��������r�@T��I�77�1��ӧ�ȧ��XU���#��ޱ�� ��d��v�C��z�0��\(��0I�;���8�(N(��0�[cq��};�^�dp1�����a/��n:�J�$��1��-����b(��7~k��mGZ"��x�[hM�9��z�QhFv
���T�����[�$�K���ql0�A4Ȇ� ����w��<jw>�Oٷ��ٶ���ص����N� ���\ݔ�^<=3aj�IUJ���L�&�dK��l�����7J�ĝ����{�%y���Eg&����,��4/�d��*k�t�ɔ�tg�ZT�}1�L4q���4��ZhC�����'�T�AoY��]a,�F4��x۳ 3��	gU� ��P��B�]4޷���؁�>A&����wsj�
c�6^T>y����=� ��T�g�3R��~�l�y��CU�5~���[�r��7����a\���"�xdEm�1Bi�)�^p��V#a�n�)�1��~�
�n�^���]�^�I���X`q���W,����ե�+?'���J14�G��y8��/�/У(�d���>+@_�.�����K�pji���4C���k��R�\�[����Es3X<�L�zL��|w-R_������������U;�7�
�=��?s��Y�C�Ip��>��+�:�D��-�6ʔdt̊it gݒ�qԈ]���Y�V�>����m��IS�Z�\�!g1��r�T�Y���6I `/�´�ڣ��n�L�3�n�o�7H�_4h�|��:���X�r�d��1��DJǃ��!���i���0\(��� �^�Ϩ?-�&IC���2nصq�:��f2�m�$ܤ�K.e��6�R��Ӆ���s����t ���+ݓ����g9�7gr�X��cFƪM)����d�u�V��Y*��HDIb���u:{r��gH?������WÌA�K��<	z���}��l\8��*�@G��0��]8��{R!��|�����?�;���@��yq��\Y�*J�B.XRU�s��7|��x�RB����P[�k�ZPL��7��bҰ� y��
��6���[��$�)�73hI�ReѨ@��-�T�:��u��c2�K�?�F��tU��?9	�=�E�,�!�ey<Yd_5=ݩn�r�%�ξҝ-��M�q�ަݏnB��+�E�
�:�����C�����~=<ſ7u��:�`���)}N��_��6��bw�+_���1�q�Qe���E͛#J���N�#z�f��CJ�3Zo�V�7���G��Ȗc|����t9y��8ŷ5��U�3�M_�ֶ�6)|ܘJ���\���HxsN'x{:�Ts�5�'#�,��jX�����?��<Z���St�v'�Ղ�R�]���2���S�G�[�� 11hu�H�B�������%a<x8\�>Q�>���㪺����zƗɑHu�\-��dM7����ce�fp�v
U��vi�8\r)����=쎑�i{������m�f��	e��W��6���*�eMm)f�� �S1�k]��Äy/S��1��N���k�<�F�Ά�`����w�ݚ��楨�SpQ�?)�S��>����	�����Z�j���N�{��S��VoR��Ź��a�g���y��p�����~,�]b�Ӏ:��F�<��9�|;�w�PJ���A=Y�C�	QCG��;Z�H�w\��f����i��,1���u�3ŀ>sAק3?[ݭ��^�b�U��10�v�ʔ����j�����ײ�����,&m�^��E�q�!fW;��O�Էv���i�5h��8�\���Q��v�ˇ�,��#��wb�v߇��x>����(ְ7yGi9��vg�U ^���z����v�@�ѡ;��T�{|fef�ֶ�2��MJ�S�PF���>$$�QL�oT=�*�sp򏘱���HaD�1nl�l("��n������F��[E�V]�E� w�/��1�cF=�h;kh�Q�ư�R�U���v�_��R����|����}��Cq��7��ݟj�w�dnK	hk9�0�0��ؐ���v�z1��\r~��*vB</�q��T��q	��>����׿��pTJ�z���ցT�i���ʆ8E�k�����c��o[0	!�O ����|ݔ���&��RѲ!7p�DF;��5��'�����EBb�2Sy@��#�P���[����Ȣ�)h�d�95nw���LQ.�����YgKH������i11_�O�`5K�P!$�Q�dN#����¾�(Q7��^z���v�5kxjf�aD���b��]�{	l�a!�|�=��K�֒Y�+�\�e>�M	���O�+�<O��$
��\�d���������%Y���n��<���[]p:w�m6{�Ku ˧�ت$��6��;7�T��T�U�^߬�]-R�4!�ڢԁW��C��T^���@/�{=���-&���'|���	k���xu1t29����PB�	X��1s��K��T��+�30x���܅�@�]]����RhW�����'��;�`��q��]	>x�Q�J���6��8�ǿCUJm� ��ѷB �����.�F�G2>*��֮��g������/��Č��kbO4�:����� ����hI{cy�Q}�vS��m���w�7{-�h�УD�w��䵄K6��ȩr���}�M<-����߄����rp�M]q�r����C`!x�)�J s��X�Fj��܉���Gr�0v�Y��u�=�{�`��Iܖ�.�ٔa �I��D��w2*�`�zS.������4Y��)QF*��a�("+�yEx�E��������'Y8ȼ;]4�Z�a���E)���~?ؠ�[���/w*�{�,��26�+x �f�}ݼ,����h��#�W��'D(���˅��R?�bk}Ќ�c:��b悃\���Z�ɘ�b�yP
Q��h���ApEb��������r=��(���	�Լm;Z��P�5 �,�������+9�ɼ/��_�&ؖ����.֨�ڙ]��tќ|���p�	^���0���?���"�[����Թ*^��f{�g׍�Y�+v�9���ߺ?����