��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�v�-Q�π���*���t\�D�8��ؽ��N�'���W�)8�k�!�g�ì
G���ޜԂ�rq���6�
+�fp=<������;�74�m_\���ka徤�p��ا��q�)��ęŚ ��3��t�v�N@���
�ҟ���j��T����s���5���H0.������.#���[`�����:|���j�
��	Z�����JŪ"J���£~8�j�.��@X"d��Q�̍�*-r�ȶ�&�����T�L��(���� �����Գ'��|��cJ�1�`
���!��I��mn��U�࿭;[ߘFz�#�0�SU��C-��(�a�t��Z���)0a�^A����̴�=1W�&�.q�.�{�n���H0�j( �U}R�U<*#�|>��Af����a��&��/eNv�k�:�d�j*ŵ��ׯ��M��
�F�JN��Ӧ������`�}��u� _?����RV ��eǍ� �%G2af?�§w��KӇ ƺ�U���2�N&HǬd�<}��
�S���>�Lp.[�h_k�4��|�~��J����B��h�_�w�bn�/+������8����ԤGX_8ΐ�������w�B��b��猶(�H�/���9}�%ҍbE���  V����
�kuo5��6~��d�Ay���?�&\�Z�!�MȀ�p�J��9���{���+e��������Tn]��� ���u�g��t���O�L�xX���=�bE�n���Bs� >Bv��ťt���gUȥ{ 0��G�y��ih&�o���H�%��9�3�to,�X���V;'�">���tAɿP�U�I�/g�t)��[�"m7�<Z8��*�j3�S!vK�
s��r�R��̑�@�$ۓ ���Q3�x yC-�e2�4	�5Jڍ8��O�w�0��B�{��� _�`�ۨvCOk��TgsK�o�xUZ	��}��܍�^�L&lT��u�i?bP��p�C扞�n��{�^M���=��,U)�����9�K]rs`�h/!���#�\Q�;���{�:��ޫ�Ɲ��B��w�Jw9��M5~1��l�]�%z(Sb�s���X�艧 :��kT�)Ec�N�+���?t�6�S����`����F��鈖vcK�$BCl�G��_�y�B�/�oDx�|��s{cS!��6����	������:qWĈ-���ts� Ռ`f�xD_�S��^7�q�FJGy�kW�-zb��i�[��
�� ���r��]�oJ��=SvW�y���/>D���k�:�UIC��MP�w`�y{m|kS�CA�@<�=�L���������"����K�v*\�����_�SE�z��`3"֖�o�R���b���C��pf��x��h��%�o�Z|��u7��~��[�oH.���y*���M�����4���$�T#��v����j/Y@�s:s�SCQ��ct���7�nH	!%���|�D��Q��\u��Ā�C���~_k���@0��/TГ�����u�֛��N.쮦 1�(����c _����S���^a�0ݻ)�� vM����<�B
Bʜ����b�f'#��l�*�p<��*i�{���|LP<��Uī�:�j��s�oi�B����"�V�A��|P�"\-Ο*��t���I��b@��}��aY�;R͒��d�(B�>���hq���`Ȟt�cbq�'����ܣ_9��~�ed�`t���8&�"w��/�x_sь%�72�E�x2���d�k���^ڛ���,��g�o���$؞ &�E���Yw.�A��\��"8�xOwH�.>�O�-�ENH`�(T$�(͑��9��G��dD!��q&�:�	V�$2YUxM5��T|}�`�-���P������]K����\4��Ru0;�;ս����(C�.'M� @]����ʱ2ؒ���w�z�Z� ��oި�-j�.�ZX��0�r�ַ�K3⚿}6J����L�������0 �	�8��{�����Y��mXvo�W[�Pd#�vw�3�6{��,��O��8�� +A�g��x4��i���Dl̽:���ɹnH�od${����2B &��9����k���u='�%B�v<��]�(_cF����)n�<���a:�m���!V&� c;:<�H,B=>8��PA�օ��i�l�G��Q4[��-q�M�H��e���ۯ�? Y8`)�Ӊqȝ��r�m��2u�|��>�������4F��k[��]�7m��5�a|��R��?����=U�� 	�Z�$��2o`"Ȇ5�T3�_
�%����x^�[����]�|8"�
��$YF��*�-���C�����G%�Ǎ�R� `R�6X��׹6��j���+۴��|I��p�ӽ��Y�gs�y�c+���jXg(�3�f6��H�̼�"���
��mi#�晫�O��$����R�Q��`r��ޟ���=y:�����AU=�X�t��҉��I��Qu��.�\�t<^�*��(��Mbm��&t����V_�a'�u��)�~�n,�phPR��>��mjM��0���0�tW�ŏ�^U������j3�ΚfU�|��xa9�TF ���`� �M�u�L��	
������Ĝ�U�f�ı�1a�JF%������#(���ۿ �08��r��#'�gz�8i�N�9�~��W �x�%�}z˄I�(�8���přL��|v�����7|��L��YvΑ��PI)FD�GV-
EC|݊D4���;��-�!?�=�YP{�ʵ����{ߩ2�/X��y�O)�z�[@�ʏBF�%3� �`�>��k:�l�x,e�oZ��;���".��c9g>�C��3�v�Aޜ�$ݶ(Ck��M15{չs��Zr�J��7;�Y��#��K����0�nS�?S�|��=��M��'�`׸��t{��Pѩ�֣�TbH���>�[����%N���S쭴J��$�W�B)C6�k��e/��:�Y*���X��P�]-�P/8�b�?�,��_�
nz�����^M|t����/P�܅��u��<��gټ�p����7�������b̃r�p(N �Ǒ��d��I��P�"�K~��hԐ�dlH�I���8\s�[�U}c_.�&
h�i{����C�@�0��HvhL!y/Ǖ'��+��-Cz3�!G���f��k8+M��җ�����uu�D����Ȳ� �y�T�\�6�)�ݙ)&�
h�0Ń�����z�A�q�k��gSp���p٬� ����'.�Z�%�v%޼I2-DgM��������
��iy#!���������)��'B��L|�\�jN�hJ�q�+����D�Xyc|,檳�T�:��T�9fT�	�^����+c��������u>����(�"�A�K��l�?�h�����p��KښEJ��ԁX�C�*n
�?�AKY{�o�sB~j�~T����皊�V�b&�1�`zrT�M��{�������� n��^�����o�B-��_�)9;�t�A��u����*�
�j�6����7��D�.�ij,�VZ��ͦ�J<VYl���n��3���*�ȳ�2TZNHY��&��'�
$��wɭR"y��m�V ��F¬��Q^s���vX��P�<y�p��i6d�S^�Am����R�Đ��P��^��y~����l�_��a�Γ����8�g��kL40q!���iJF�!�9��1z������:@t^�G����D>#R�
&(ď�Q �9.�!�9��r�d�L]q��p�5Q�84�L�Rk�)�s��j(�/��>�G���#(��&�'��z��{�	.Yr�EMY(4��[`_�<^M�:��<��n@-�6������F�)6��&���8f)y������V�殘y�w�M��k<�P��#wB��yFPؠu[Zy��;Sȟw}G��Փ�J�]�	Z�J)���_����^5�3p~�}A��8�C.u���dh!�&U��e��D��'jj�om��o�q�ԺıOM�5��"�q_me/z������Z<��2Ͻ���5DG-*�*$BIs{�����P�O�P���6�;R���\W쌌��i~`Q�VτA��7%�?h+8���0~�Q>a�"�V�R�d�J��Z� n��}6��XUL�7�L`x%����Ɉ:��q��������~��7Fl�����r|�6���iH�	I������M����1{�q�"��((+�=�G����G8�_�#�K�m�j4�	V�kvI���k42�Z#�8�SUZ	�ߖu'-b�����l)G<3(��X7��yL�/��g+<'�\�s��qz�t��<P�M1�ۿ�=_���Q�7﫣��ۻ�=�Re.*��/�D�)s�O3�J�7mQ)c�11�.�~nK#oڝ`��,�y��K�L5T��U1��;U�����|����36- ����7���<E4���������w��-cȧ��z��0��!�1]R�8F"C�}�y��K{s���Զ�;2�܊�U�|����J�5Рi���z��">J���s����j����p��Z��=w�Q�6����}8�ڳP��Y�jN��U)�axUL�ňS�ض�.2%��[%�'jV�~p��Q����)�,%
�E�s��eE�ܭ��C8m9�]|E�Q/���P }����X��K�ܽ�k>eV��!�Z��e\v~]t��o勶bӟ���S�FQG��� u7�/��je�E�s���%I������<�6�A}-�l�=�yC�;��1e�/�c��{��㯌Oѽ�U��v�M��%MqOэw�GU��-�1W�f����cY�P�:�j�3ֶ�9��a�,�.'`Rk�CE�i��m���2�:�
<l����n���U�V{�2#Y���c�a�A��HDE�*ƚ�)Jm
//ڤjvպ��Q�O���,cQ��&��O���p��y�∽��k�`�h��	Wɴ�o�c�gd-�,̰pb^,����4�$�MX��}��B�x m��M�b��q������(�G�9��b��ò�����A�@.H��(˗�B��n�.(����^�r2E�K�M�jX�/:��lhε�d�$�/u(m�1����C�>���Y��.M��-fnEW�NM��]�v��W�j�x�6!=��~�,RZ�u�`*T�Tehk�2)���F�b0�G���2������(g���^+Y�X�!��/��.6=EUk�Z�L���D3���LD��(�<��>����ȉ�3��AL�YD2��y�]�b	~X�܆!B�s�qB��p�O%ƽ`�Q>������h`Ƶ����l��`�1�u�9�K�P:#�Uݻ%ϱ4hn�3�	�K�xt"�����0���M�D]��ҚlM��@&݅��Rз���^I�CG<���ժ�<򵭉dݔ\9/-! ��� �SY�W���ZT��?:8���b���
Nt7���M7"G`z�}g�
��,�/�M2��p�M'_>�{��q�p8�e ��/0Lb&|�\��{0T�w�x6w4��bx���z�� �i�W�G �2�D���Aj|[d�}���	�����U��Biu���NΝ u蛅)���{�C&ԓ���C�����|������,a�-���Q���sV�n`��o�k&������(F�F9	S��BH�2�J��`��a�D���3l��ԩ�W���DG�=�-R�L�A��A�Ǐ,@v�����3{������9��Z�0�t<a�I��酳,!c$�3�EM'j�u�O�UU��6�x��0[�;�~����]h����s��H�2ء�7L��=v��E�_I!j���{ٶ�� ��\�>4p������Qާ��S�Yͼr�܅��<�l��U�k	�ui}Hk�bKRnlkΙ���ݗ�1tm��0"|Pd�$ʧ��Y!u��s��ͺ�*�YZ7%��C��iY{�w���X���}�[s��9өi��0���a����	".����@�0n�����+X��N�u &V ���K�,Ǖ��l4��?aMaU�0ۃ�=n�t*oP��|q6Y�z�汫��B�o�_�Kb(��>E�ݻ7\�d��Q:�Wv���w���
8.E�d�w}�Rp�\�G=W���r ���,A�������DH�R�J�u!�����x����|8b����8�Gc�?�9��)lV}旓�n��G`�"�"a�k�tJތI��:y��=HH�y3@��6����U���9Ki���ѡ�����w��%�&��u!e�'��|XN4��N*���g#`�_�Siȣ�r�W��m{B�n?Bn���'r�0�_	9�xI����%d���Dt�Gn5)p"'t���׭�x�C�������ow�n����R]���0�Q��脡�D���'�pw���ŹvI/,N)��|�Ƥ��JM�N6��p�qT��r�/��O*��ya�E kc*��&mo�E�����(7?3a��ix���3����������n�80r[(���br"f�XQ�'ϟ���K&\��)���ZW��X��$?��&�͉��-cq�#�,�0��e�Ck��q���#�m
0GWY��9`!H��_c�)8��X����ЍqFRZX���X�>����dy�e`D�)tRONR��a7#��ӫ�{%���D��&?�p*���w�F��V��S�x֤m�ra8Ǧ�[�r˦jrޤ���rJ�BX�����4	�-��W�m��o����c���`�h]�9A�kS<�~2�nʺ?�~�h ������QS	K&~m#m|9��z�&?5�=�ڨ��_,4{�5^jI�ɥհ!�ذ�C��ٳ�g1��Z]v�
���/�&jލ�*e19zY�	��-c����yQG��/�2]���C
?�L���� �|�A��<��̋]���C���kSHD�bp�k%?��gO���>�Wcy�1M���:-�m��rJ��d|Z��� �����b�y�*�ݞ^��#�F�d�����������!+c"�(��τm���P�Ί<o?�������J�Q6���#6h3�ϛ�%�o��?����;�e��2�֠�O��
�|LHV�ڠ��z�C��@B�H41���_��U;��9�^�^d�Ã�\di�#�/w��Bz�����&h�t�-��1��ǹ�_)��	f������m������������R�O}v��)��O�� M�*��`9=s�yq1���h%s��yc�[J"�S�QӢ�_�:����sn����RXj֡��'� ����$m�i�B �x.�M([�1�ˊN�F]����·JSۓ?�rI��#��u֐��[T�2��R�����K;��8ލ��~A�K�tq��x����%���1h�:G`�\����Ƭ�Mѫ9�3e��s�R�V��r���ԅ>��s� ��k�N�\r�)�k<?e�o"�m��!�ǿK�Q��`Dp�i��VN!�W&�/��3����]��W�������ثH������~3`���>��־΁O�U��HC�r�W8�$ɠ�6��j���*�-�ܰa)����X��blO��u�R�>��@�_/�Lq��K[�$/�tUf����`�ie��`h�3b��f��UWԐ��,퓞v's����W{������I���ci�9���H:74cEh���a��n��g��_�1�wL��
F�.�=Q��oD�)���XϢM�|�@ǳ\��do0_xs��(���M��*�1�h�f������$K�����F ��0M&�+��M|xO^QjY`�=�"���߃󲉪|��gmd���_��J�!UI�Hg��
ə�#~������� ���'�e�օVt̂c���ǐ�:ީ2��Ш3��^�E]+���'����:k`�ߠ��kh�6��g������7���סa]�[�޿ ��
�_2ݪ�t'wZ�/�~Y�9-��1)��)�!�����A-�V�AP9Ҝ���	J>P�=jE9���T�:�*��yO4�^TF���dbb"> &	�-�w8�`w�=��g�>o%=���낱.�$b@���E��E9��|��.*��i��'�D�ù5��y������W��߸�9��'�\)${�0�s#J�C։c�J���2Ai��l��/�4T(��S-����L���k3J
��J�F��O�4�|=�'��s�BƯ$��<C�NŹх�5_m���G�Lc��L��֊h� ��;ekn��X�C���KBq8V�鍝�rW�V wO�n<�������P�=2.�ޞ^��Ycb��N�5�8�l�	��E�C�y�:��]�"63w�%�i7ȓ`. �����`�s(���66^��풸1�R�����1%z��#�kI�_4���R���mM��}n�!�h��M$D��b^'�2������L,�5<v��������t5Չ�ɺ/�����M�!t�dѯ5:��:6�N%�p��"}zv�-��[m��*i
��?Gx��kΏ�X��&�(N�fl��(���$MO����,����[27�����s�Њ"}#ǳ`73��ʕ�D1pH�ke��c�,N��ne�
�+�Z��t�Apd;CQ�T#�n�)K�Wc�u���<& ,Z/���3�����P��-�\:m�F��w��<�A0��<�=#����iN�xjWW��7�M����i�� �t^�zr����h���7��˝