��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K�&	UT.y�J6��}԰�c�"�� �.ŞtG%��\�&l�@%[(q��
�-Ћ3�E���_'�0���RqVw�{�v{D�|��*��C�HP����h�����+�>����6S�>'��]��U�7!���Q+~p�xʒ��2H-}�z�(��h\7����@|/D�͡n��!�h��e!;�<��8� ~YL�@�S�u	@�ܚ�Wmer�P���J٣)V�)���ه�����:�6ZtY���'��@�p���׺V9�9��/e=�>��`0�H�[�
���xi�ZcZ��ka�A�ϛ���.r��ş|��0U�L���܄@�`��o�J|>�~�����-E�ύ����S�֚��Sy�S�+�y]�P+_�I�&��;>�qW_�G#��-�,��}3�R��j4^T��h\X=!B ��K[��Ⱥ����
V��9?�����J+W{2��RR1�Rm��;���h�\��9s+}s�Ojq:9���{��{�\�F�V)�Yb����J������A)��	ה�d��� 
�jp�B�S@�F��>|�U��ہ�2�K�|
D*�4���ΡH����%�6g��݇Y��_x���P���r17���%K�9�x}�7��y��*�N�u���@'DZq�� �{����(N�+�}K��h�������ُ�磿��:u_�+8���gC���?0�̶���5:�M){�0ѳ��f0�z�^ǔ�D#ue���u׀��U��>��,��Q�m���Eg�����ԑ�I��PV�4[�af|��|���6��M��Y��p&������#e�䵅�G�������ƞ ������\n��n�`Vn�Ƭ�?���ђqYy��x��Ϫ�r ���n��2\=�����Y�w����xs E����	�6+��jL�@��|�\-ڹy�q��a��W�=Sp�P����"XvJ;�����c~�q0tB�P
��ڬ�CΞ�5}�����ѿ�`�kJ4Sȿ
HkE_?�)ݤ$�bgT�M��F����.j�3���USU:�)W-�0�^�Y3$�Cԓ��-ѓ7�����>i�6�ҶH�Y�6P�D�0^4Z�r����EO��5d�$�+��d MP�sA>M���#�f���8U�H�<��qu�y�3�'�M�:F��Tk�=�/�a=�+���C�y�[��!x�������+J�ڬaNu��W�`��O����^�)j��E+�r�����j��xb��*͢2�xeR��U��_�e@]9J:c�>y+�n�	-��~M_����L2���%���e���D��q�	]a�����PE�u/ȰN�:��0A#U�Vt��W��_q��*�u&lq�F�ƭ�m������5|���k�4{���e�;�n(� ����b~Z-;O�S�`ĸ;gX�*JќdA �^����pN�������7�`!��Њ�v�g|E*Y�*͠-/W�흍���V�R���5�~e@���$(��e8	��jĺ2u>�m%R����@X��|�S1�ؠ?��mG�#���_�(��
F�_��ok1okɌ��$i�iz�M�4� �{����N�*��I�~��>��Ϡ\zP���O5-A�f�8����%Y;Qk�u�&�˨x��QF �g���{%~=I���<C��#^� �I)l���|�Sv9!�C���(j�k�R	U�B�X��IS��&��Z�=�0�B]�)gt�y�@�l"�c��O�����x�7�}����ּS��3P3H�//�<�>\���cA_x�Noż
�4#5�kQ�fNz����}��ѫ58cJ�.e1�A��6k�ey9ƫ!(��Y˭V��v;�so�~Ɯk>�������)�?��7f��nk�

���O����i��F�K"�T�MK����si�)��@�����g�|&N�oó��⤈?����ʣ���B�}�	���/�?��b�6����BA75}%�3,�q�������ʼ0�I�C��(���V��Z�9¦tmt2�k� �Lx�9���)4���n���m��x����@uHp\xe:I�a"�f���o��;�6
,=&+�� �@�-!6MI"��e�i��^�/��������2���"�;*�X�:�e}@{*n�X0Hҿ���2�fʱ�>��}w,;���	����	��38�[X-\����� ����w�^�U`s˽/�m��}r\��ǯ� OX��ASr� ��T&��'`���*�Er� �#����)m��Q;!N�@:�>�g��\�߻���% \���/�97���K���s��k:�DK6j򙴰I�Hs�4?W�]���'��vxں��?MF�?=��׍�ru��轹�J=��p�z5�Zn��F��2�u�1Is�->u?A�[��MI�� 4#ʘ�S�!	��f쎈��(ck�f�Dw[O�$�.��Jk������8��L��q���$��)�5�а�ޭ�7��huJ	�Ln�C3Z�:2T�/`���oa6��־��O�8�s�0�����K����G�G�Ɔ��J.�YN���	\���Tbg������(�<��n�<������ Gl��^�O�aI늛I���Y�тč�)�Ej���mY��c���42+�t�W2�v>�!�X2$������ܔCj���Y8���]m�Z������(-L�J�����sA�O��Ym;�elF{	� Z!5R��P�[���Ak�#��_4S��܁~�EǕo| EWM����h�9`��޲N��ЇpDL0{�����k�9e.�_;���_�h~y]kvh"�.�������Uj�$�Ȗ�[����K&��b�X��J�Y�=�C#���a�2��j�@UZ�nǉ�1*D'W�ow!�[#0d&�w@�6��v��1GK��ל��Z�`1�\�R5�d3-(��K��86|�N�"m�q@���,'p�m9�ޢKV�f�19{!�q%ߒ[�TcDy��݆옱4:4��m��Vg��_��@/��N��.5�m#������/zۊ��P��e$w��!���#����&�b���\	 �>V�w���LA�s$i�f���z���~ܿ��6ΞXN����pSkc��l��,�6�ci�$�G�7�4Q_�D��M���� �By���zm��h�
Mh�	2P
0�`���Y�q��V��w/��!�j,�B�[P��} ���=�R[��6�Ά\Ͳ|ы�>]m�B9�}��x�o��rW_��EU�h>M�i��P��I7�6��!�\��=� �n��� CX-ڟ�r��ww*�u���%�(:��g#��Q�]�q��v�l��p��ѪM!2�>�xk�-��H)��Q�N��]'���@A��=����c�'{��"c�����5l+��^�gWVo��`C��C��^�w��C�Z\I���h��=���8o�{R���p�oz�[B�Qm���봏���	�Y�4��a<���Ϗ]5�� �@#?�7����K��St�vpH��ƞ�̦ f&��mM՝ꑎ�wr���F[����\����w=�'Ä*���?�S	��b8Rѯ��O�n�-}Ñ�o5S�����9������P��]�2��1�0��X���<zlۏ�
����޽ߖF�<QY��]pA����t�=�ǈ��p���}���=jED��٫v�Jyt��ACo���ۏt��R.F��s���6I�����M o��w���K�n������
�ؕJU`�9.���N��XB0�;��>�����F���q�nv��k��d!��2q�e��*j����7�!�²�
���sֵ�(����@@>�vS6�Ye�D��c��2
��'�?gSSx�`��VC�ȃK�uW���L���A�P�GC�׆�]��E���ȧ�����ȏOp�"Nbh��I�i��0M���&P�����x�p����.��G�qa����HYԥLګxA�s�@_��4?�K�� ���>㟶?S��S`����B��s0y�j�
D+J��W!�|��K�R��*p����w�������J�Y��B~B�ө@T�����R4MD?�dS���XܥAF�:���憔�:���#�'�.�˥�Ꝺ���;-1���/�=��n%$�+�xn�AI�@�K0iQ:�(mx=�*(��v#�y�~Z'?��;D�������HsA���f�	��ْY��H<�˸��"��ۖ>~�s�gg*�D9�p�x������H�80�"Y{��G��K��O�V_޺$4 ~���(+��"k�QI%���|$,VNI��d��X ��rL4��!f0�=�m��s����[�+�
��Dg�?O"��>L�N�_����T�7�����iG~�>|�U�9�z��|#��nIt�TK�k��=գ��Wu<Bo�c��_�6�<�d>F ���}�fvbYG�vj�����c�+ϛ�I��Lb=.I����Cލ��bM	�)�9D yB�v'�6���\i4��PX/��v?V���Z�0����Nƀ����]/뙌�JȹJ�T������.�'&9ho���-�����Y�Q� 5B��lt�&?=RG��I@�z�`u)48��M8�bX�гf�u�?�Iϵx����T�[�1W*v%���v6-y��=����wX9-��9��Ls��n�o�ܱ���t�|m�|B����{�aCh1�i{��`����H�|J���b��V��q8H;G[Ѭ���(�o��!�T�y���h)g����XD��k�
S�lS�	�_�yE�qqum.`����(�k/��Z�6�	�������?9
y-�d�X��o�:�����dV\�qç����K�5*��S���H�3���wz��q�Jj&_��w�3V&;�@nJ�%��Q��U¾��a�z2^�i�r�Z���`�����,5���A@�o+2��J[ԕ�!p%wӫ��Qױ�b��b� ��0紞
H=<��� �gΚ4�j�l*�=�\=�[>y�Ɔ�e��Ș�g��I�����I��3Xb�R-��״��Wv�z������Wc��<���0g* 7h4��f��D�ύ7�s��ķ��Z7�x�g��
���/���yF(��_�s׮n��K��-�D�`��R�4Y�i_�e/�����˩{�-J'������Jp:�jnQ�x�)S[�4�Ĝ:3,��5|;�Î��X����}ϭ�B��`�K�C���i��[4�ܘ�)�o���)��U�2y+���hzVN|�խ����a%�-�tu7w�R̫N�l~�n���VI�\�_��ye|��6�D����j���
?��LX_�������l�?v�6Pn�>������_�0��R��(��)`9�Efu
?wH�|Wu�(�Õ���]k �?V���w
e*��S���k�"^�X�R�
*���`G|�oI���؛pr��+��W4+�l���|>�AM�X�l���鶶�p{�Ŭ�T�{f�Es\a��c=5���˭�Q���z.^����B��~����^ik׹;�Y�H�iq6˗w�U˲�4~jT�̓�/~�f��rzħ��Ӻ���<K���1���}�`��6$���|2��  �C��}�/��Q��,��X�8���c<۲�fTBpߵ�E�׸���'����PLo��([��7���q����}SPf�6���C�����~f��W�ZG�Eڼ�Pd�4Z2_��±m�=`�5������ˬ��z�5,����-l�k�,��>|5*���ך�s�����B������(ݞm2'&P+�P�(ڲJ�=�D
���R6�\+��ǚM|�K�|Gusc��L-���QmG8��Y����zW���}S촾�����,���^8h��=4^�itN�/k����GL���=]!YT�n��n�6�%� 	����ќ����0my�/=7<Ob:�\D�����u����!��H�W ���Ɉ_f�Q��\�|T�dP��+Y�R�>}�2���d�u	�>��a�����XdfуoB�خT=b����et�_�T0�E���%�S&>���]B�@���'�Bs�`_�Q�.֝��n��E|BC��O�ɒ/J�~CZ����J1��<�`�/��ݨ�>LX�jj����~�LmN�!�
�8I�O��
����3�>>�C�O��ǁ᠂/���r>���0(����s�h�
f�6�$�����ݙ�-aI�I��6�'��k
�nv3^R��n� �ٙ�F�P�I�T�K_W����d�x��� �k��w���FF� ]Z�I 2��|{=��]�^����F�`.�O��Ϧ�Mf�����/U�|�"��xڀ�!��$O�lx��0ʹX���SO~퐺b�!p$�«Y�p��c�\��
�SqU?��>@N:��������K3H�j!�I��V8�l�Q��h��r$����%Bn˗��eH����Y��qT��8�&5���~�_C��-����B�L_�W��������%f�Ҽ�T�;�DS�B��B�	D��o������$� ����/,	�d_��}������Ȫ����������H@q�IY����LÝ�z��C(j*�$?XX�d}��5&�m��*v�qu��v�u8Ϊ��"M¶�e��J�
iҺ��NqZ�C�������J�\]��]�<D���ɢ��N�U)۽�j��~�[��P����]�eXq�#���귚
ٷAA��wY�����4%N��d�a\�Mg�f��L�fç�Ŭ^�#�W7?N�x�p}�y������;����[�ku�J��4��:-�4'aLΖ��$̂c̣z�Ǹ��X��<���p%�:x�}����V(ssK���*6D�20P�sO*��D��^43�9[��(o��n�)���J��L2��E!�PT����}��#�&�����M��c��䕵xPv74D��h���V�j$���teE��o�ru���鶨
|T{��i[SSL�u�³��9�$C�~o�J��۹��s�M�h���&?n�$� KLp�r�&+\������@��u�S�V�,��H��ļ��پ^��� d�{Z|���b�AS��,n	���WU��[2N���������ӌ�/c"���S�M���:�Ruc���Ji�)���T��kY�?3hY��8��,/�1���� ;��奭�����7�yf���F<Z�w0Y�s�A.�Ȯ�`����6>Y�x�я}�r3��ӱO��n?e�{�!9���4�� 6�wBԻ���n?%*��v���˼�������A�	|��n�eV��<����0P�����	������)F�1[P|���VV+���:�7�^����hT�k`�	4�=(�O֒�VI��`\�A��x���w�۴��.x�d�Gva t�8�c���mߺ:��� �~+ծg�HsH �t�����ZK���U63� țN�Ct(�+z��8j�'m����|(赾��n_�Δ,J�g�TܙG�	Ȑ�^eٯ�O;}�x���;1�zC����{�f`������P�]%S�z�%��H�GC��[?�,�
���+���c��Uc�hJ�O>��mJ��sKE���r��&=�ߐ�+�-�K���rR�|3�\5Wv_�d�Cф!�PQ�m!qPe��Ԕ)���x5���P%;wb�k�aq>������za�2z0v;�q!E���5����x��Q#S���C\��Yw���63�y��Y�C�����;��ȁ��`�zcwo�����C��0d���	%Q�[J�y:�[��H^5��e��,�5F|�%�A�V[K���h��a��I�'R곩e�r�W|3��,�%�g��gv� ܙ��wuAՄ#���+���D�GD.��:�3���g�������K#����M�!=kb~����;5�(|w9¶��-̘�bT��8ñ���;��^���ڐ���
���Ԅ��*v��Im���v���fp�����M��a�sM�L���������{
+�p����h�v9a���z┱Mg"��iF��2��
���Vr}_@lUoQĄ�XD5M��b� �%�Ӆ��$@� z�.	"0,K���}�����������i�ɓ���P���xO)�^4�I���	�ƛaA�>�hȂ����#w?pęsT������c�1�� ���� *u~��v5�<�O"��nu�K�W���`�3�T��S7�2@LuR���8d�y�l�q��^4ĈV�ie�#��,�i��e�U��>�e3Wrþ;<���6�U+	�N��G���5����r��D>�T۽r�cA��	�L�R�q?��4�ue@�%�9����e�S>�y)!�Q�G���8Z��g�X�b�z�QNL�L㡏���2�>H��\��lh��kn�
��(N�/�H`�����z%k��L���y ��qT݈�ʚ�������mj�8���kʚ�������N������G��$FlT��穵�.�w��6�p $C�"iMOQ7�J-{މ&_ƙ�[�9aS#�<o UM��сh�A_�	�|G��(�gE�1���\њ9�"�>����e��	�1��I���¬��;젽S���#����0��\��:�{ń�+B>��Icke��O^l|���������㋗���j�1d�nD�Ȑ@3��Oc��di�Z���Ã8�OAk0�"��ք�Et�C%�YaCyi���SLd�%K^�����3+��BMv�D�1X�9vɰ�|��O��k�G��rz�9yh
ևJ������cjN��+z�)�y#�	1���?asC�YƁ_���%��;�!��բ\�����a�sX/��g���2�_"3PKeҳP��z�z����nv"��&5�b����P�kܿ0-&t����*l�E�$��%�C����w^i��kR����ҕ�D��ŤJ3@/Ku�D�]����гf(5?ULt%58�R�d�P������eP��s�q<1�z-��)fE���&_[���  ���>*�X�P&�be|�`������5"�+Q��½9l:�)�!ę]�I�23uZX���H�6��.?��_��X�A�tb�+i�'M�ֵ�r�����Bˏ3��t����'e��H6�q��빪�Ya=���,�q97SX��o��{хb	!�S,�ݬ������0߱��9m� ��+�k3�LPڔ�Y�����a��:��îg�5�"��#n�Q��ÉƊ�E�3:���Y@�'�`�k[�E�O��8���L!��'�F(�1w�7�\1L��ns�X@���0 �Z�@��47�G��1���mH�΃AB�s�Ϛ�$X��F��Zp����$q�dBy�n�4
��D�t�Bpש�����,�<���66g����
U7�{KN��3�ŀ��Qggҽ���3>o4=K��Y��!. '�[��aT���e��%��"�5m��@�qU��7TT�}�á�������`�o�ZK�W X����$�� Y�g!��� ��,4,���iFarr�G��=Vu�*f���QZC����0鉍ţt.��ϕ�/=��5��2�\o�Q�F4�Je����;p��6`}7Pћ�*���B������o �VzzeU�V����I*�e.OU��"�RY68=�h��=��j[?m�ϡ��(Q�A=��^�d���)����/����4݆+9�{t]1���>����0�q��7�H���g��W�6$?�1Ec�i��95��\ñ����I��<4��xߔ`{.,5��o^�/E��VU�����^���>�\bIB���
�7�����2b���g�Nm�"����>�`�k-���H�
�/��{fnU�7H���
��E6���A~W��IP��O코(B{O�` $Ȫ'�z�=��E��[�ʡ+bD��$�o���=so�l����̡oI�a�xE�@	�A�2Z�r��J��I� ��f�H�Ț��!�`F��*���_y���o������Tb�C�>&
��s�r�L�p9��9��wD����W�3f#9�$]Z7�4]�=�x¬3ހ��+g-b$]��Y"�<������q�~~��nH9-���Vy�i��(d}�&r��j$�:�Î�NS���ܶ�Ux1�}�����`f�� ����� k�u	�eH6<�sxx?� *�m�jX5v��	�q�Ԑ'�:j�<�S��V+��\ݷ����9H��R;�	/�Y	3q$Ԓ֣6��D:͠&m 8��#iQ�}���V|h`x3��\����dE�yu(���E���OF�!k�EZ
1�	0�<-N{G���y�����܁����;u*��ߪEw�q�Y�bc���QF����+�;ObB酝L�����+ sd,?MC� Z����Qj�I@�8Q&G��I���tX���ѡ�@�C+U��
��R*miR��x�b~�K���<�0�3&�&(B~K$���W���pd^$����}sYP�
-��t1 �\���d�&)�4�s�\CW.��\ܬ�B!�~z���y�7.1��Һj����#e<?����H�Q)�X�,0q?L,fQ�3Om��F�	N�T{��Ԁ�,��b奻��e%G��� nh"�L^�J�&$��j\+��&<��l�=ca��~�?���wt�/�&x��y�i�:��L9�F�G�I�H����.��~;1�Xi��ѠH�%ˡ��/����,�W��m 7���M�}[��$ޜ��v'ǌ�?>����M�$p�� ����>7����_��Wک���w���/p�"%�^�a�C���Ǣ:�Ƥ�5I�E`�R���Z�
��޽y+-1��<��yj7��(�
}�r�B!7 <����5�oC�<t��/�&4~�E����L��T��l��\W�$���@���N���
�$�L`'�������I�z�7hK�r��'fSKv6�+�y�`���t��T�Zm��?���
���u.z2�me@p�B��*A��p���jCОA�D
��Du�L���UYq>�B}t����-��Ĩ�@v���eΚp_��X'���]��f�(P��v	����nC����d1�Չ ������G/c�`"ǘ;�k��mD��軡,��3�}ߝa�dO�����m��L�q[��C���F������P���Q��M���;|��o�"�����5�+;�y��|r$u�Ȏ�;��2��^���!��n�n�[����*�d�r��	���YDt3,7�Ow/	��0{����0J�[�^	�B1(�".��QRɏ���1�O(����W�n6�ǯ��P>�Bn���e�+%����d����b�	��H��e��A-r^2/H|W�1�	R�\�"u���9[�GC�����;��<֥��M�t	����ѠSd�u���n|�,�F��mj�҄��X_�©Q���?��e�:L%�3\���[��)��6a������ڱ�o����
�uzT���P/+b�EN��\p�G9�B�9�
��h�)�~��qcMv�)͐�XmCW���)���S�R��[2"m���;F��Os�X[�i��kAwn�����ڕ�E���Q�p̀cN�����б#88yg���*l�O��SV��/�5v��j�Ѽ/m�@��݋��!�-{@�]+��7�|iNǩ��<K�Ȉ��ٿN�|����)h�8�*%��������X`y"C�A��)��&|���$���oB;�	f���p���͐�_�}�w�[��91q�U����ea:c��i=��<I�5�:E#н^[��S]gi���Nt	܂���-o�mհ�Ӥg!�����F��Yg @ǝ�_�1A���
�h�7I�0m�����]|a� �N��B��<���Y�}I�[���~�]�6ºX �ȃ�W��-����g���hP쨵N%]=��/�µ1U0*�-ނ�=Y5u�Sɘ ��/9 ��`�Ԧ��ʵ�z�q���Z�(i�YJ�o��
s�kV���R<��!n��%ZJWxb�;�sPl0U��#|�&�:�n�<����3�M}o�|BSAX�Ū���4��X1cQhFm9
|�p����Z�M��;�ROM��9$�wy��K��΅t[ �Q������w?������ڽ����7��U�OG��T�qO���i��D\����ф��M��(v�k���]\�+h�c=�I?�/��ѯX3���%~syX�3�m�����ujl����ʸ�T�*}b��[�@��>`���R���R�C ��X�y��
ߊ<��~Ect�K��4�K}~ޭ�%�ݮI�g{,���P^�e���W���`��s�ƥm>�/63�+�ڍ�׷�P��ə~�\u��88��r�Wֵ!�(0"����:9x�K Rv3 ���E���B��0 ������3}�C`[k�\�C6��~�1% {k��Ս�g �ʷK(�F���s��^�Sw��Bb=q�z�'�-�R��"�6�u��
: 5c1�G�"u=G��]��M}v+���'J�?��ag2bI�]�:��>�J�9G��SMgU���nn�0u�*__��`h�S�0n-������e�`�!��WBs�)(�R�0�wu��0^�I�!��&$dE&o�yŭ5��ҩI�6�`oc��2��R*3ƥ�r1���e	ɣ�$�]C*�"��R�ǆ;����5��@S";?)�Yt�k�A���Ř;�U���6>h�B�͘tp�BN&=p�?�aIR��(�.�7�F� %���Za�"�/p�pDp�$���PA=�f}Α�����i%���#Q���D�GAg
�kx�r��a1Nr�QP�;����v�\�v�t����@���FQ�� �����	����:� �����6P�AO��~ŏ	]r��4\���[>����V���q���O���`��+Oj4���^t\��r?G�_����ėq��w�Ia��Ll�K�ׁӁn���okLB*P?)C�;O��R
���꒞v��q:�q͜��"u;�O�&ڱ�.�1��Ձ~��h�~�u����D5�������r۷@�5�\��S��s	|FAx��r��cC��C��i- [��?�e�OR LL���W���텤e^̓^4��-�\jcX�s��֙��G�Ms�n�K�Uk1Rqѯ����LS�8�b�<z{nA���s��x��q�	J�� H�`�(��L�,�8���7��g֏�5�7�Ѱ7���x�4�C�)˸ܖ ��7�ۨ���iTOZ6!AhQe	p�1Kt���I0�ΓT&��pi�V䪡�mƾ��_�!vwR<.��[4z�����t�J��J4��5�Y�L�Z�
Irs%A]�	i^5�٢�>$�%]�>Tm�E
���C��e2M�)f�� �cM���:�(�p��M�s5ܡ��q#�(���$�+ǆ(ҧ��fs��bUV)0�a���wW>����s�k�o:����}4�����}�R/��|�-NB%�"�A�t�ܥ�&�x!F1.�`�������;�b�9�!���e�U�����G�|�\�0˼��	&v6L!a�� �MYX6���ܰm��Ol�����`Y�}p�����s�G&���t�u�N �D�����B����kM�2�f@��E�?�S	eİ�-�LV3�@^J�j'��WU��	��O�וI�Dd��)GO<��� fk�.�V�EԈK;�~m�Hw�x��r�-���]p:⽴�ad��+��0u.���#�w\7)�č �GHdD���!K����ӿ>�[�m���8.u��A�ڰ��Yސ;m좞��!$R{���5h�9�]q��X���	��-U��jJ���c���ά��W�)�(��d���nv����}�;8�0g�&ޫ�-=������/|\F�8𹽥�������ZP\��=���բ�Q�|�_"{ˡ�jI���ƪ����m���[N���͆?~�x�]�oj���#b8����S��s�i/k����h�2�e�f�hv��z8f�]Hd�)��u����0$eQk�h�jC�:��CP�Τ��U>{�V�vj��C��&�뛦�ˤ!���_���*�I\�v�o�(O�B��g����ϰu�e\I�m��K!A!�P+S���T����!���rn�H04���8�4�����FZvDla$����]��I����
��@Yp+�B��5�R�8p<3I� ���B��KkH\j��7��V
9�FFm'��I�y&n�����t�>; 2L�TL�hH�Q�8=0�*������O��A"j���%�pN=a�E6t�?3K��M�j��܆I�*S��O)���5�ńɜ���
��<d�~��+�
�}e�2`,��(�~�Np�p��o7�՛�ř��m�i��g�O�df����
�F�a^���t�'�[��pc2�)hn�g�ٓs�z,��s㌢ן�cfĎ�t�]�V\4�}}�%}Y�/.a{z���`G֋���+�Hy�O"�t~����v{v�]A��$�g�C�6���I�d#��8;�iIIz'��E�Y�-������	'>��H��N�0k3Q���%�/eU���Ez�>vY��\��D,O�ݖl��[�eg��q�"\F�_�l�8�V#�pR�W6D0�؀�q#��8n�����Ě��`0±��_��<�T�387q>3�U�i��d#�/�9��KSt\ٛ�v�i=����*`��7I��Vy����TP ��o���f� KG�%��>��.�����+I��۷�)�:BQ$�X���ZT���DȚ���c�Ɯ@/��2��w���z�2��0��5_ �n�F�G�Q�{ޤV�� <�ի�n���	5�����e�O{�1�T�N@ì��\!��+'ok�T��/"Ț���@�����i\�>�_���]��ΐ
����ͨ�*sD�i�^V��Y�V&K��E�w����_0����I�����~�W1����cD��O�6X2����[֥|��?�0��Q�b���: �-�@0#�g�D~��1�*S�y�K��V�Z�!������j8*�f��ß�g���d�j��!��:_:@��1�m�|�sM)· �E�Z'���K����#:�5e��5�&LJrf���_�ݝd�J��nm��,��fx�.���@���?�Ťt��~�ԚF��0fl�+��}_(q�u�wd.����"�*t&V`�9�c����'��9�6]�`�_\>?�nvB!W���2��`�r��"$��k�s��c��݊U���3�컚��ݹ��Pg)�¡�#$��A,3=4�k��󆑢����@���~�(�bG�0�A2����[q7����������g}7�,�Sεk܄$pe��յSM
����g�!Ua��}s$���b�1�P'BJ˱ J���_�^4H�]=g���z7�C�V:8��"�	�ї�	ij2!���f���
��4�I�@���osrhEWͭ>�OB��2�b�<u�M���p+��s*�»G�w����a�B������0�n'x���e���t�X'8�=Jۑޡ�st���*"��@xF������g��g�����#���9=���Ej�����Fi�#�����E%}�p����W��V��pz��J��=f�nU��r_�{���o�^�[\��VI5T��h�7đ�%+��X�L�A7�	�F�>�_�4#}��F�wm=\��#5ᏹ��4̇��4=;�H�G�uk�
���p���f��}Y�z�Q���O�d�"�R�g�n���\�;�[���(�|�pm\�x��4�8LhS@�����7�8�;��r���/����{���:�S=� u&ӝ1��l��G��vwTS��s6�
)d_��>~����5��	�Q��:`l�qZ��t�,1�n[�Ѳi��S���B����fH��S,Qk���g�~P2q��Gt������W�	 ��Jc�P�J�3N�>�1�&���._�*�]8��p�M��=�E�84�� jl���үl�)�Ym�7���j�4�p��'
P||F�{�����=��7���V&Ѻ�?��Lƨa�>�����@k�SG�����Q��FB��c8K+��f�׋X:�E�qm��&��qsu��?s:�j;��/�M%1ؒ���V���dn�s�j|��8~ �� C�b~4ᒩ��S��VP��psi��̈yW�����<�U;�>���3s��D�Ǥ�������5tע��l�����Һ~9�d��[�CtP*x��C��w�O���v���QȊ�D�k$������PlL�������u�)�8�<{���.��GNk�5.��dH<e��]iH�&2�c����01<�����򯓴��-CY멢�6�n�5D�J,B'�$��=O���/���2��56�Fג0��	堥=ZFic�~0�%l��/j}��Ƅ,��7W�K�<;��z%�n�0y����Ӎ�D��͂u���6�1ğ-�K-]��D�#|��O�O2��$(�"���`�Ԡ�r=���R� ӯe�����8ǌC|ϯ̱Q�0��}� 
�Ի��:TV�-�"�7�u�;��T5��'��4o�>�7r������#���W�kU	Ә�L��Ӕ��SȄ��H�����pX�L���G�N�?lr�9Ut�o�Bt&/<o$���v�5FW�d����Xo�~��o[��q�	)�a�F*x���5T͓F� ��4�Lb�e]�2�y�e[uC%�%�G�~���$n�U2*���R�4{�R���� �ոbF����v�4���l'�s��1���0a���v~j�eS����������j~=�Uf�7�4T���%����`*������WAz�T�}��M~�<E����_G��WH=4H�+�*Pt_�Z��%A����2������ $*��	^��[u���<�S��ע g��O_��� i1B�t����O�a���_�$5�{>8���=}�4u�
N��\j����>�}<��s�E�Z�d�\8T�C�V=G'�gP��'�[箣0�s�"\К?��"��	�ⱘ�N�IB��R��$~�S�ve\t�]��/Zy�q�Ls+�WG��tV&�T�	�ނs�_��|Z�wӞ��o�0�o�
t*:�P!�պ�s�thc�A渳����;��M\8C�ziޠ��+��'�D<��9ñ���|��DC�++��=�cC��WӐt�D��[�&�1��`ɱJ��jū��}Kx��ߝ�81�B��������=��Ap��ί����� ����Sb�^�"���^4hb�S��t>���z��4�=s<�o�����K���= �;͓����di58^3����HƂ��{���n�����wDh��E�yq+Y&��S��%Ɋkυ���Eε\�5\����U��xe�̆c��!H��7�E����A���pۡ�b$x6^�����nH����hv����ce�d�?D��T�!w�7��y@};��E
H����fA���a��=�ҀK��ZC�}^�_to\>�@H��vo=�%Dy�E�̶]��b��zܠ�!�{�n�yR��u=7�O¨�;yxI�{I?C-�ޓ�R���~�G]��T��Og����րV��?���o�X~���yC������f�Q=g�u�ף�|L���<%�7/ЗA�K�bB���Y�D/�����o}��'z���Ɲ���d��S������~�4�Q�J���+�^��veb��o� yv�%��JaT�p��(Z�]�ߑ�ޭ��6�ɳ�P,^�Pq�7RtsɅ�7����)}�`��J=�`��⮝kQh����+���s��6�2&����UF+���(�,i��]����Ƽ�-#�1��0j��e���n�&M�ɛ�a�H7��ԓ�n�@$������)�)"O�l���+���kZ*4HsZ��k8�ՠ��'��?0M���C�I�u�B�њ�PU��U��4���ϊ��	ObiF2���7��a����?%���LF�,(EI4�I�9���i|xNy�`�>9{��ߨ����x��k#Q��׆\�� ��+Kp���\��\ �`��!��X�@�E�g�s�k2`"���:�Au]{�j�}��Sa�/V���P|�����c9�xE�E5Z�n�#Q��q�Y�?&d*	u�bû�.E	qZx��ʻ=zz��/b�# KP4�}��������/-͉n/P�|	�w�fiBY��N��O=Y�|�)��M�U�N���F%8L���P��۔�R�k��m�<��8	�s�:KSި��W_t�����\�6&c��Q 0��ꃧn����n 9�)�6��ƪ9��	!�9�^�B�f"��ܶFԪU�Rlz�=YpL-�k��<+����53߅}��'Dt���Ḅ�BG��5�m����l��#�\�W�(T��&�$�KMQ�J�Bb(�&�%��T]�@(��&���J����#��eX��r8hp<ݚ[�L�r^�o�c���S�|E
����$�]��a�*cq3��ЫNe�h�,^ˬ��L`U�qlt��RTht�y�J���q1O a3��JJO"���|7�
~�Ae�E�?%=:�Ϝj�%7^?v�&�w$JytM�3V|�ۅ�J�.�ţ��W���T WV8�r�����xմ�͖�d5U�i3a�9Ϛ�_H� ���1��Ơ��K�uc|<(��P_KɊj��2;к,��p�'.�H�e�p����k������[���G�r�b���⯹h7�J]�g/���G#�˘1Ho�a;P���n�%��Խ�0i��B/��q���%�W} ����P�6
�[K��4حr��'	�2�Pm��nh19_��1?R"F �vc䞋N�5����>�7�KlJ:�S"z
���?���A�!��A��֬�:I����Nл���M��O��kv�r�e���y��`qpY@�m˳tb|:U���O�C2ٵ����eDk�1��϶\_d`,�O�2� ��W/(�,�)���-��4��� T�nڏ?�4�͏뎳��Kp2�N-�'ԾBI��<���D8}��)�7P�1�E%/Hl���j�^�G�U֭p�jUP{e��ы|��V���\N����I��fH/p=l\訿�ͮ�4����E�B#�3���g i��9��2�Oa�W��{���xy{3�:�F��0��~ɼ`3���?���4*�ڶ5����^RV���6����iG� eQ���^�����ӂ�THDx�E����������C�;Q8���z�� �<?�Sn��!r�t��T���#���zͼ��B��2�u��p���m,s�Z0I:��twч	���Mdx�WD�����`u빖�_����s�~�~Z��E�� �"|?�kP��)7���Z��߿��������B@���Fq�e-�22S����<����7H�|�n�9��gS>�s�֯�Eǫ4��Dd�B�԰_s�v2��N�J;�Ov��}v/.���u�@i:iR΂�M�x"d��LQ8č��K��F�X�c�M(��@ ��3�ʐ��9+��x�4�;�_7����tڅ���qhQ-��M��ȕ�{�R�|R^�߽����[2��kmY�z�փ���30��=Ӳ-�`B\~D�E���wϰ墶�-���mjr������&�Q��ĵF��:f��4�*���E ��l�:_�ۼY�_��U�>2�~^�@�!���-�0�܄*�i��U��w��J�ڽ��a�I�6�P:s}��"�*��		�ߚ�p���R�v��m1E��oy%TA�M�d��ߚI$�LG�$�::fcN��=j���X�rIӞ�ux��ܐ�Ib��Ǵ���۫�D��Na;�sBYk)�3S�>b����	
�嵐�G�a~�󯧢���X{�k��m,����
e��gn�MN˽u�CQoh��0TՈk�x8袹z �*�t����5܎�#k7~8�k@{�ф.x0�7�$�\�����v̄�4u�g��7c�t|Y��<�#vH����b�R� aL�/Ai��L1s�����;�&�k�!��P�?z����pK�Mw##9� ��:�T2aA��ٔ2>ӷ̈́PlS�.8L�o���o����}|�d>��|:�\�Kw�܁�2���'*+}�ժ�x��/��/^^O8j��^O���ÖuE�t^�U��;�b_(ـTD�f x�M�Ք4J�.��'�j��n).~j�'��F�R�0�l���|�y�pHtYO�H	�P���P�7����x�*A[�c�UuI[~0�&����$HQ#HD�mA�f�W���\Ǟ@!uÓ��S�؞m�s�Ц�/�������Ϥ=��$xҍ��A`��-x�|@�ŀo+ә�OoM������?��g�V ��y�K�ڄ�-���b^��TёOd�
��,������^3�;�^��+I�c��.YY�<��D�er��ɷ]+�z]���L��e�^�n��B���f+�
hC�.���*�)Mbz��������Y��;�>؅����ph��.��Qqv�<ŉL[�����.�tfkP,W�%��Q+�j��H�� �(EcE [a���$$�H���Vͤ�ٻϧ��M\��b���T?a���1��^�\�Ȉ1��-f+���B
ѹ�����j��[,�,23�s�<������OS��˾��.�ʙ��Ȅ4�ڻ����'�k!�Sǲ��g��D�'+vÑ���W��Fq���� I�C�n��X���f�W��_�\�
�:�Hgin}ic���# Tܗ4	d��Ŝ�8MM���2�paM{�w����%#9�žν�Ld����E���2��5j'�l�;ȸ6����&����QC�X����CӺ`�&�㘖lcL��Gq�Rc�h;J�?Q����=���L�*L�Ҝ)��bx�v�@Mf�}>9A���/`�R�w��@<�W�4l)�F�°xyFg2I�5�J�ڱ.�i��t؆�Dwr
��I�C�^Q�ɐj喳��&���Lq��(�n���d8zݴK�P�DJ�uG���k-~Kj��D�"��fc��;��������U��d�&T{�����1��[5O�ܩ�����*z_~ُ���깖G@O|��6?��;��ry����������n��;	̮'v�3���G[�kռ�6j��>ڤ���P �^J�gD���3}�:���|I;�3r>L�u�En-(��s�J���P,\�q��bmDX��{X�Y���[��@A�=)Z��Юڡ�\���V(G�*�U ���{'�GF?њչ�{�A�B�l:1�ã��S�����;M����}R�4q4ii�wp�)HU���y}qx���`��_�-E�T��>FيQ�+.a�ތfv�SК�6�t�~V��˃��B�	��OK�eG˃�c-���՝�M�*#�6�����~ -�G<=�$�2�YZ]��s�a�S�P6PA��@h��3��4;��F��G��q� c��@�!x{��ꯟ�@���Z�c���7;�̺u��?��.�-�u��f���Tr��9�?�B�T�	r�c̬�Ƽ�h]�O���jsD�*׿��:�E�:�ߛ`I#�{�#��mk7.�z�>���9����`=�?�_����n!|K�d웕��p�>�0����B��U��W�G�3D9���Sf����]���:��F�>��V���� ����~���">�e���z*KH��ۚy����'�Y��L�(d��]	M� � ֤��D�FUU���pm� ߄��)��B���_�Ft�xJbcG�<���u-��E���Ί�ɏĖ`	�"�âz����"(�7��0��ʝ&y�4��V-�>�蒚Q�����N�Q�.>��Uu@����ԟu�t��3j�d�\�p4�%B��hoDЮǣOlډ�J�0�8k��Х�2�o�+d�^7@x
��O��'�d�]����	r�C�����滬l�3x�#�G�@!&B�+��9ooF��p��Xۥ�f�t��4��N���Y���� J6�ܴ�b�+Y!������x1�S$����g�f�]B �T� t1�Ό����'���5����L�� #���UۊjD�Fy��4"�C��[l̴�a�(n۩ϚmQP�;B�̐4�Z
]g硼���U���0���a(�W���C��P�7D��T���Dy��>���Yu�)���V�������T�����y*�H"�'T}��i�< Gٰ�_n't�����n�����J2)���̡�_쌙e�g�W^�D�x�=��^��Wq*v��*�&����R�w�f$C�+��'��;��"$��܃�������q3hZf�x(��=���H�U���55���M6f�96q�h!w�J�e?���|?���ӵ0B.�ƋJ��D����F�6kB���K������,���|(:�1��.�h�!�^�V�:�+/|pg��
��0��c-l=�[��%���R��e�]?L�Fj�k�%E���uj'�>y�↔����{�x������Ђ�.�1��A2L�bmn���!�����T�����KG�Z˜)e����'y�߻��S~%��ȏ��,@�+<{�	h=1\�n�� �L����QOL���3߭8�-�u����V��Œu�z�u�	0��A�,+4��\�8��q�ݖ�D�U4#��8�`1x7����E�{<8K�6pu���<�R�}��'4N�o�?�m�g������i�T�
8�L����?�0 i`��:��o���͐z�LԪ��P�R��~_+�u��5�x��=�2����h.��������~Q\h���%�U*���P0`p�!)���ĩ��M��a������"%ZZ�qk�ԛ�9�E9b����#����3iũ aܷ(c7�v�����A�����$�����*҃WF�T��&��X3�XQ�͇m�v����I6;z�ӳ!\�0S�����Vm�Y�3�eQdDiug|-ׅ{���RZ@��[�#��>zҶ:��L�����k�z�a�p+Ҁ
W������e��vU� +�M��nDCrn�����i��|$��@��t����YI�)�uJ_:��ō�	�,���K��0�>�߹�Ѹ
��E��%�
�ѰE����	m�r&�J�EJ޸�9�4�k���d*D�|���!�/܃�
t�?�p@�3�����
r�~$V�Y7Q���e_}��¤:�Q~��";��d�nV����Ώ�d�2�ʵ���]�D@��=��
�HT�~!/9	蘬��Aϭh�8����5�ń)��݊�Q�z�Ȥ����z��_,�j�L=�Әj��[�˝K�@*tp��e���f��⦙���|�b�`{"]��!�}���Yh'��S�-��̡r'��i.���1��Fֺ��ß)�]�1�򡒤#�1�ў"�\�;��V't��3�ei [%�/Ơ�̺b���X ����-4ܯ@��g�냺�u��@���y{�l�����[ȧ��a��@��E|H��3������)�|��=��Z7F���@鱿1踳o}��鰬��ע�/�X+��Vф�#!��/�-pJ�ZЭoʄЄ��hIj$(p}�_�
T�Prr�������qɈh#�}�[�A�^�=4�7>'�]�7���"�V}��<�s����+!4|�G�	|]��#����i~巐�w["�Ǜ�{zVOދ�$ؘ�ـ�1����d����臑ͥ�9�el�T���W�r-`�̱�U� uR⾃Yÿ�CD�n���Ɂ��������m2ݐo�2���M,rr��E��t^>Ig0~?�I�3wA2uo��z��2�G��v�R��:� ���]�
��jr.S��?�l����Gi��6�(.�*���a�&�T���ȹ�ݾ��Y���S9�olT�O�--���4i@2��9!���w��ޱˢF��%���e���f쥜U"�Ļx�Cel<�� q�qV�pA�L��(	a	��pۓЎ����Tۥ��|��d" S��`otM%��aa��.Ӯ�m}�F:����g�EOT�,� }5��{C�S���_>����#�H��q�5$�(�T�qc:��;���T熬қ��
�Y<M��#��H_��R0�oDS��:��F�)�}�:���2�yй���e�\��R%Y�(��:���Ʀd������i��e��=��7n�Z7�7�U�7����\D&��R�W'�Q�w]'*o�y�9�����#h�mT7~���Q�N�T������${M������MZ��օh�W�mӉ�/I5�n��@`��%"��1����]cJ`%E�`��(�1W��>( 1F>�"8�i�~��ɬ��S����1��B�	�4��*�u���݈�ĥ��w�/Y��Wf6��R�ũ��w���9.���g��^�q ޗ7���kW�p<[Z����-O�L�y����r�S��2��)ZD��8��`���5�`�L#zݖ��6'��!c>��9�{Cgt�C"s'|��,����W��N�t��[�v�H��Z,�"�>����OFN�\��ʔ�\a��y�+i��M�~��ƾ������v�_Ȟ%e��{�?�p�@d� �j-���<���x��i��}�B*;6x�F�2( zj5���l�c�߃U*�{"��]���.t|C�}L�?B�S1�s������(�B�E_�P�`{xAB���$S�n�uj`zD�p[�*�Wt���̗n����g ��l*�5 �g�.=~	m�G27y� ��Б����[A�&8�>Ĉ`�)����ݞ� 7:QF���f�����x4�" 2H�頻H8Ċ�7��B��
#}"gY�����F��#�۹i���ڊ�S��F�������'���S$���<�YOD�C���ҍ�`�!�d��7�#FT�QCB���\�r:I�j�+A��Yn��
EJo -���|Rlv%/����SB�%���3�gߟX끜ה��◣�ךh���`viN��a�vm��(޼�*`ci���:�I*�P�A���%��?����zLp7��0��%�����7��F�o?1�Z�2
y~!G,��P�o�1[����'�����R`��^9�B���賗����^\-P��Q
e��W92��?�ٴ���p�%�Z-�b`���.��GN�+���ػ�R}��S4ܐ��.r)L��u�<�zND%�Ge5��-@�~D���Q� |S��HQ��ky/����^Jj�ካOk�a/�h����o�ϣB���	%�O��A��@����ha�����g�i4���t�C߸_4��RLG��⸼=�
�o	먫Ƭ���YR�}`e�H����{�)����4�NO ��Byk/?�e�Ts��{ yZ%9dmx��&��o�)�Br����m(	�Ĝx7
K��L�Aߴ�l�*1������q�ٷ�v�;�����f�
��5���54)�{�����)�#}��>�B�(����n�Y�������=p�Dti�$.<1a^q�ˠ�3(�[�Z(b'z��)����Z�9���dbi���/����[<��X��t��Ѕ���� U޲(�����Z6�a�~Ҁ�A�ߴ�n���K�bj���b�<�n��SA��P���9_�����-�Io���Y�.�Յ|��I�B����{�S��[_J��t2u�n�]<���(WL���}�+�����n����9�����8�[[�<M:�)@(�`�Y���h�EB��	d|���['�H;�Hi/0��5~  ��`qف��K������CXQp���NNh-��E^�"	����C��OB\�ܮ�1�'�����Z����YBR�feA��*�d���w���5�:���#��V5���-���7lj���&%4ߦ��}���]xTACu��wB�T �	��^�vu��e��K89N��I@�S��y2\2���暸v�8r���ʧg���&��z��_�\�:�6����шZ6�P�Ѥ�CЗi�8�tF�yޖ�ʫ�+Q<=�VG�MB	�:��{�V����j���f7M�� �P2G�j1�&��f�0#�k���u��.�dh�w�"�_��LLL���dN��`^!gd�k$.),�/<}dA3j��������h%�]�e���H8+���B���j}�Cs?���>׭�.~��7��e���`{��}q�79r,T����/l���rS�z*A�Lz�2��\v;�����:��z�/	�@S>�
���r�:猀e�(�ʛ�l������_"3�v�3�:���X����d�`羏� d�Mk��n�瓂�9@5��jt��Y��‽�Iɩmp@4a��&�@p7�ϫ��d�����J���!�S��dN>���F��kv�:��jy3��o'���3�P?�������x& �HE�T�e��:(��iO�+��w9o�B]�
㩉W��| ��#��(ӫ��p��@�L���{��� ��'�HOft��@J��:/@`V{IJq���R�X��]jJ�j�����3v��憐��^h�k��<���I���c�^��x��k�Y�Π�S�@���чd�����3���,yę��5�QAI�up�Q�!r=�ы4`�ƸY���B�լ_%��vE�L9e獤�v��o���E=F�ХM2掱�&I���^�X"h����,{vJ�0�0�,��I�rC�Pa5h�n�Q�ע��r޳QJ� "���l'	h��t'b��� Wv�GOa��I������i���(��O�
��7�WT�W≷�.�r=8�L�	+��{�m ���=�K} �꺑A�_c`9<�t�x%����j�)�N�[���ԧcD݉�0���jd�y� �"$��F�v�u��e���B�I�k����������h��?��c�~��لҪ�(SdE:�d���.t�z�zh�QO=����߂�,R�1����a�T1�CNډf�^L��Z�?.�݄6*K�5	����v����i$�6�\g�������6��"BO��M�p���k	w��i^�f�P�����xf��ǐ#z�ׯyV#:^�l���% �f��HN��L+�q��ro;NQ::��`�g��b~J1��D��/Wv�KI�(�	T� ��B��s��6z�R`�H�/B�d'�1&�P�Qĥc6O{�iK~��x8EV�@瑆$�kD�4-�@]��I�6u��M؇9Kq�1-ь�c�=\�k��#�n��]܃�!���/�a��f,Piϝ�]��!e��T�^���N70h��B��Y���Gj VAgD��'m�kM�-���D�Ӌ�;���!Y����=0�E}��,���y�<#��l�P��OR
�bT����u>{,���;��|E�$��	|I���j��G�����+��I���߭�����8,��C�UQ<U��UO�I<�G����&/�"39��1�/:=`ez�ʕ:��4���mv��t�[\�9����D��8S;P�8Z!v(�^���ⷕh�4Ó��5"o�k��͝�9T������h�#��mƎ��~b{PL�ڈ���-�} ����v�f��-��Q�}l�Il$��h���N�/�E0-�\�3�����f��~�lC�_ݸw{�V��m�|�M93(_�o.�ο�گOtdZy���O2��*@�vG�����W]$lM? ;��p�1.�U{��NOl������u���N�#@e���ƾφhF@�j����4���T6p�$�@�6y�ۙ�VU��P+gM�2�RmBY�9_ze'0b���#�Ǚ�˅qP\��S���-e�M�&
�n�^C�n&�|YL��A-u��z>涎Y��ui�s�n>�JߔF ���~^;蜆J����x�A�1L���w����d��o�{��`��`
+��Hy�x���$����uz�uy汙P�&�9 �u}>������,]2�P)�'M����P�0�c6T̀jB"���u�����֠��R>�W_���zp�s�7��	y��
#��>8l3"JR��ڎ���i�Uܽ8��>N]ci@��������5Y,U�,|��5��@��^JQV�/:ثa+!�}�N��Vy��ZdQL�)S�ΐ��Mq}&8=���\n���A����e�q��1=!H��.6v0$¹�4Dl;Ye)�F䋺p��X6/J��(�)�x �w�f*�9���=��رy�̞̀v���=���[7� *�צ������j�H{�D��R�ٮ��M��V�'��{�%�T�^>+�� ���|��N��W���H
�/o2Fz|	V�����~ڔ����;I��1�{��r��;ё2����(t�՛��h��$d�P|DL��2�8)�D�L�GPT"����p�yP׭mg�I�E\3ꋞ�H0��H�E2�}��lvy<.'E�	J�D�E3�IP����W}���x�>[��v��+�o	�щ�{��Nw�mnF�I]���*&�cE�����z3�Oc�lJzЇI$S?Wzg�"��÷j�����Wd��RM��:�)U�յ\��WӖ�3�4��R�O}�����.i�ʷ4%����KL��i4]vj��W��̪�4J�]��|�Os:t��"�6��v[��ȉ��"D	>X�j���Y�[|�ŉM\�K]L/�2�HB�8�e�hZ���̿8�����#e�:��h�� /����'�z<���Fr/����h5��u҅��M� Ź�=�fyب�O{��X�r��W���(��\�{�<QN9�7��zJ؛C�g�$�>�7�(щ�/U�	*��?6 �ZJ���H��E�8>�6�WJK,����H�R�
�qt	��DL�~B_�:���u�G!��N�f� d7mb���^�Zn����/�}�^�����o�ͫq�Ӱ�\�HL0��g�+���ݟ�0��ʈu5�pRէ�P/�S*���b)���aWJI_�g"܎Z���Ik�%u��˼������<@ފU��z���%��js2�q�?T�^��4�r�B?O5����� sY4�m��GS`MD~�}�#�2���+uNAQ`r�E��xT�k���,_w��@&2	�XMcQ�U9�5,0.���r>�h!M��/`tK����xg�d�;}���bsOU����Y</ȝ[�@�͟zb|���ĢaD����q�'A�dӉ"X��B��O�*|u�����#�v%k���F��-���߈��U.*�+R}�� eJͨ��Ց�H�ȅy�E���-j��swf����A5݌���d����<���ub<�zu揣���+#K#��(��/�u����P�&��XX�ɻ")��e��.�&z�1�7���&�l�.��y*�<�������	wi��m��Q������q���7۝&\��D2�����?MS����'���ԃ g�JZ��1�^\�"Y�o�f���^"���+�F1�Dh���벁C�;1m��.����9(��`�BC:^-|��F�f���ܢ�e+C+�d]WP�R� Q��ZKl-�gJS=�zrlA��aht�6 `����]�	���-�E�C@�M�`�I�5 �Ɛ�A�H��3b�6��.�t�3�(�W����9%�he.���w��J�F���ޱ��u��	�w2G�)
�D��+qu���ncG[�1A�7��%�/���^�ĳ�FU��u��4��g��T��)䯵�jʑ��(��S�!���ڛؠ���eq�tuE@�2F,�U��|�>�O[A�+�[�>w�"ҷ���'�+_"����5/�F�r��|�VJ*е�
yϷ����ξ���Z�Wcḁf~�"�_�W	N����	�?ߤ)��3`��s���j���Z�Kb)֘X�z?�U9�X�k�� ��0�W�󿒓��B.5f�m�a|S胛�#��t�7��Mq��*	r{DD�� �y��q����/*��u�YF��1�j�δ��	��X�(�c�%��8W.&E	9�Yq6�#���E�V���+<�/��b����'o�v�h|b@���NZ| �3���>"��q�� �^D�$��v���4�إ�"�t��� ���M.�����|
���4Hr4��ﻃ ��>��H#ha����}!�_���9
��]�f�C�T�J�(�M���!��R.���_64���0Z4��_�SI�X3�ae�xp-�l�Ť½m��}�ǩ��i����"<a��KW�j���a��i)�\腲��OFO3��䙱�-���-�p��{��� ވW,QP/��U�P]-3d~���OR[ؠ���h�kd����g���c�vx8�w�$����'n��j��%؎�����^.����*�	A�������|����朻@�#���5���] ���	�"��+��:v>|�wm]�8X��k���D ���]~���
�h����꽗�-W2s��2�R����F���~�[�T������Oew0��t��,o������ �{��O��R�B�Ux��y�ѳѺ\Qks��iq4\��`���z�٫Q����Q�P|�p���\��4�պ��I.ۢ#��yE]P�y �G�v��1�)�?�Q�fj׻kPP%E�+[c�27���H�+i�qzQA��鶃�'��d�Z>,@���|��+w�(O�4�I�;�3O�vV�������s&(>�Vn��ep���r~�Z��'�E6KL�y! �(3zq�n2B���^;\L�=��2=;Y��Sdl� �i.��PB�kH��:�����{7�k�\y"�L��1о2�u����a�,S���Z^mM�5ӴS�1*s c��O�a[�,��w+t BvT���TU��a�<N��g$�7@�3�%�������J8��n���EG����5Jl�<�]5�eo���{�O�R���l�<4y��A�O�}��QN$%����(7Vx��0S��SVGpA��2��hf5�s��
�	����� h�Gpe�� �3�E��	e�"�p�wν[�$�xo$Ƌ0˪!��I�
^��'�$��.�V�<��K�z�;����Z��ǳ��Iʪ�Ӈ-m�Ǜw�"��6�Z�V������8���dMt�=;b7�~i$+k�.BZ����%���1�k<�	`�"�x�D�Ex�'L��u�$V0�?�~s_o��$9v�ϣ���W��7m�R4��_>��i��H�&������H@˜|?�^�q��l��Y�����G$�$�0�u�I[�҈Ԅ�+�ූ��m�m o^	��C	|8�?!�Θ��!d���׭y��ls���G����4�W8� �@�s�$��Bk.?�,�`�኷\/��XZr}� +Q���z���c���q�{>�Үq����Qx�A��������
��.�|4L#t���`�C��-d�L��
md��Yu깼�+���i�,p��'$wR�.2�Ur"G|�v� *ST㷅�΍��ڏ(A��@7����B���[���߳^1X��'%7��0�T��?��C��ig��.=�$c�9��x�W����j��%�	0�X�s�ʢ�ȵ�ǵ�E+��em}"���]Z��:kz�7���	�@���Z�»=ѥ=��Nt`ZM?j�+bh��<��`�ev�0�m����}���#���R{�NU�i(����]�"*��l,��Bp�ǈ��X%�����]�?(J1�1l�M����	TGq�q0�∊�w�~?��V�0:"�;ŷ�.����uA�6Mם�j8�d-$�ݺ�R<)"�G-ӕ��:B�sv2���b�]M���af:TYxP�ݭ]�yG��'wCw���8+N�l�-�fe���Ou�B�k.���qoz��/���s��~��S~��|�S�O�Y��(dG�W'���R�+��F������=mf��z�ER�P��V+P��|J��F&?ۻ?���J�2��� Cc�`">9�Ud�K�3�"I�l^�r����&�nV������<�e���k���$�>�^y���Q�5���P\Z⩔/���Rw��]��_�&z��������NLW��D��� 8��C`e
�� (�;w	r0�a�	`�x�i�1$�l�{)��lU��p����z���t�A��t��v
��b�����<��\G7&{q�<��([��Ǹ%�)�����x�k"D!G`C<�	��B���?o���
�E�<"ҧ]�Q�ׄY�s���:��!�jg6��"o�o6�y�f�cݖ��j�'�N��oáC�`�JѬ�!@ ��9����G��E<�A�d�nM��|ps>f�6�݈��{��mz/jY�w�}���G�ˆ��5J.Ey��b��ҷƑ�IE�,��P��pPƃ<)��[f��������!�0����E�S�Q�P��:L
 lB����c^�����I�л=��'#Y��'1��gC{�O�؁��bf�$���1�q���>!!�#�W$���f�b�#¹�R$(�ob��- T���j��"υ�����D���?���&���.DQRU&ۓS3@�>L�@��]�qu3��cE:k�B��p����h��3��� ���t��U�;0�m��Y��2lYѨ�R�Q�N\z�H RAa�G�K� }l�ؐ�):���r:���Q��1�Iw�H���أ-�I��C�����c�e0��4��j@���,���G�Е�է� 9׆���S�v_[��yHs��W)���Ӿ�8^�q�ơ�BG>�Xv��Z���IReT��HqL��#�P�Q��.X'<����>5���ׂ����W���+�jV��t�3Q��ϛ���+�kq�$�賰�y?_�'�ASo,�'b_:^h���>��dd�ÑS�LY�c3�����n���+O�|ho&������81~b�������DΩ3�$@]�]�H�h��%׉����x���*�:5h��)\N�o����,%?$x�j�J��W�BV�x�V`�I�9�^�7#�'���X��թ;<*9�`��>�b�sg]�W��G!�I#Vud�yDѲ2ff�W���/�d��ta�PUmX��t��m����� u�P��/q��Ⓩ����%�܍�2���{�2Q@p^i셯y\��_1��E�=�j?���֠^_vգ�XF�!劺��9����[W?��9Y�8@*:?&�0����w_Ϙ�E�E�P����]��G�/~�&��V��!8/���H�G���x6:��
9�j�w�^�TT��#>�˳�O�Oɑ0*|��������:��&W��m��0����[��LN �e^C#`\(ܬs[�0~�$�c}�2t>��V�[��̨���φ�:`�K�ߓ���T		��vI�hn�������ls�j���B���eO_���I�\5F�6�����*�?--@�p�����\Wl:���O�;��5PF���Ku����Ԓo�/ޟ�Ե�l��.�+� 奛�q.}��� �F�@������S��6�M
�a��Bl�%��۹�2�y.�nBO��4�'g�J����&�g������ �ź���q_��(��KcjyX��S�Ozqx��q�aqD�a�y 1xߥ�4�޶�?8zo_c�B�T1Pj,�F ��U�pJ�9ϭ�|O\nr����6j��E��cz;�ۂ��¼q���D���&E��FK4[2pa~��D�5�^�⏟Oǫ��yW�~G�6��.n��8�qn	/9e_��A��q�>0T�(�����,�ؼ8Y�������B��8�Q�G�l�D� �4��iy;�F�Ұ&�����+m	qF47 ] �ͭ�גY³����Ѥ�T_2ko�YT�͊�& �=x��=�jB�U����P0�Ǎ����h|K偝�W`��m���FD�w4Wg�Fr��7d��S�ׅ5Z�]8^�sh�������?�ΜD*��s1I�= �zy�v�� ��e˥{��
47� �SX�o� �8���x����
bw%q����A�Ḵ*�YF
G��ɞa�3sL����{h��"�_��'�74^�o�� �9�n�~���ai��C���
Կ��(�֎@I����b�5��'G�h��d^foa*�҉��V`���v�W�(�u:�ѫ�|_�-|u�'S�M|���]��zl��޻���Í����YF3���m�Ŷv4[@@�T������k���}x�Ӯ��JTU�ߘE,1>�O���
���.?��;r��zn'w���B,�"�-��`�$�����g�\�(�q��Q7|Q�8�C�d=�=:ξ7��qR�����Cl�ht���*ٺ"�G`�"���a���"���gA��<���R ���ք�Vi�����t��pJ[��\'	pB���"(�	�^qi������qхy!bD��U��ô��E�DJ�M�)j6b'���32'v������n'R]=�����4I����@��aj6M[K��c�h��o�-=�Y����7���`�|��Y*εj�G��ؽ+�������m��m2�(
���-���َ�JY��#����9>+t��A�!0��,%�Bu�KK�d'Q�?2���$x�}>�^�}��[�V��+XL)E�V��Z߸�wUPY��ѹB^F�S"9)[˻�k�5y)�J��ħ|�t�;�� �:�l<��m�4������_��8j�����4��!;�ќ�����2�AQ���u�aԉ�����h���uֶ����$TEs4d^�,~G�;~A�G��C�#�_')g��t}�)������Bwq�7�e�/�^T��_&Ǩ:g�C�ǿ��pr��n[��	s���+1�`�z˗�]��6A�;�1q5�Ѵ�x}z7�4W�>՗VY�!BlZ��"Va�S��}|��f_si?�iU��+|)���yf�@e��,�$J�`9�쁶�����X�̀������������2'����@�oG�Cs�Gbo�[YlJ��g�-����>�K��R���:Q�]j�������V�\�����v�=���� ��DBF��?m�\����TѨ�	Ws���H��U��^����O
�nx��˳��{�&��ͽ,A��<d}վ�����F�N������2�f��0��y��M��F���C]��#�bύY��d�^*QN���$ݲ�0�J�A:��ad[y�r97�y2��S7ʮ/�r-b���E�Ȟ��+>�Qm�:~�v!l->+�ݣr���f�"�I�=���P����Y�J�-u������e���rD{H�O�`4]���d�P�CCȢ��&f��㒭3͆��E����d�����a�޺�\��W���~�|����R���$�*1T������r�WJS.1��d[�t���v9g���=��߻�ñ�i~��(�E�"����`B2V�%"-��k����Џ�6;���`�n6{�����1����P8��7�x������syޢ��o�vJ+H��� n��ï�����ߨ�n�U����w�mG���s� �r1[^NT�߀���3�n&W�:��NM�A�f�"�}ݣ�_��B�(e@�s�C�SW�K@��=�ReҌ^����yxn�ĳc�re�t�g���E�����'(����_6���Ja�f� e��l����O��\��s�sY~xƐ��=@7�Luݱn �B&^i�^,c�a�$��\c?�y�2�{<v9���!��k��)��DY-zt#�t�|�lL[d�¸�=zlXɤ� �2p�+s����7��/��Ҧ�F�z�)��l����Jk�n�`��(��n�b�`2k���e�k~��S�IN�+A�v�a0�u��F�o��S} C�~�P�o�d�-3�F��i0�w��MO��k[Q�%�OŶ�YS("cA������+�0���1�O�iG�~�<�p9dAD�H��E{O =�x=VE�9H��Ie' ]w1���8�H����j�u�_U�=]~�)�c�#���Jp�}x7��H4׆�~o�LyM�ɋ<r���VUD��)WlE�Ɉ0z�2:�=��<h"��ׄ�E9Q��a��DWE�kV!Ҵ���+����M�!X��H8TM@��}N����̀R%�t�7�<�kO;rja1�V-jm7���h�gRk�C�+&��Ţ�4X�R��<�\�G�j
n�s��z���`r�P�s���R����H�ު�|��f��2�w,�ih�t��ٷ�&!�x(����!�1���jș]2�� L��fC��v��ؗ�~n��H���ZH�k�C��r[���R��OR��Rs�r�� L/1��@�܄n��ߞ�w?�d���r���|���r���9����n⺖Ӗ�I�%Y�v��#E�	��`�M����y��cs 
5mOg������5>�5�����@sf���+��-CpB.$o��M��kiة�u�,���E?�]��ڧIl�؛�*�.��� �a�WQ7���Л��{� �h���ݰys�8�H��(n�8a�G���V�����dh#�٭�m\��0{R�b.���D9�sK�����SU�K�i�_�f(�j��2�\`2hK2W���K�d�:��s�%ې�������m.�����%Yn���yI&�$�{R��'j�$���u�Ž��;���nr�!���7����Od�ͽ�1-�}V$[��)-���.�u4�s"��*2k)�=�v&���k��h�f�������.��X]��Ȫ6���x/�%A��v���1IEc�KY!G�?8{|v��#Z ���.�p0�8`�E>�}9��ljM�C���U9y5E$�Y�M��@���,�W��{���Ve�S��4_���k��(���6� Y��2��@�9���s�/]�%���bf�D-�S	5
�t�PMm��8��ʵ�^��a!����BA�WK�wއ�{�����%).��׉ Yn`d��+v^ڸ�/�I.w�"j�?j�N>N�T{#�͕�b<uʏՒB
�\�qًiW����
)�"�B�d>�0h����ƙC���:_6�2|PKה�g�6��N�43Ô�4#u��V�P)�,�����.=I�L0d�?���q���:�Dno������zZ�F�ĭ��A�?������~x��W�ڠf���ǧ��q�����^�I�{r`�W�T�X��[�XEhK��Q���gh��,]��9��R�av���I�xx��ғ�8�� �@��l���pp���펉��/4h.�L���{�����6��r������dRzޛS��̕5N�9����:5��Dy�5�@�#-���6��-�6�qb�	�C.I�.�HWb��/-C̎����x����5Nx���N\Tx�B�4��~hצ,�aj��?��QC,�{4W��f�
�E�HO4�(�z�ȴ�.|0ؔ��`� F�ᅯ
��rb����o�qN����3��*,����!��J��H�U����΃���k^#8��1k��I� ��7���Z{�sa�AJ��r�b�
����b[lt7��f�S~�}����^��	�Ӧ�X0:P�v�l�7�h} ��JgIg�s�n04(C�b!	�JQ��,$Ǉ��`�Z��]eY�A��Rb�����a�ohѡdԱ���8 ٻ^�a���3��m�9W��U$��
&�?��!�X>�T�{oG�E���s*+�*Y��ȅ
��������죾bID[����o��7#�1����8���,�n�G��\�RC�I_����u+�z������V��@}�z��$Q���4m-��<4T��(��/T�Ț��.̓�@塖jAo�M�M;�b+~*���u��sC���i��D5f����c��q�1D��^��7K�-����_��ad��+'6khIA�/NFӫƮ流�n��`�v�����~à?*�fl�r��c%G<�*ՙ�Eūx��f��tzt�m
��;��C��X��F �����Xʛ���R^����-n��8*�+��A�8-9�x��)�=��gʹ�r��8�����[��u�����}�%X�����VF��Ύ�}z�E�����s�#BQ�IOD�S�h���J�s*��1'r��y5@l�CBB��0�E��E
�3Ŝ @ �3E���l_0-��=C���@$��|˒��έF�~��D����j�az*��_�k��Od%!:� ��@�����q�������c��2����.{�>�b����}���|�h�u����Q3��s>_
����4�Ror.8���}��hq~ůZݩ/���̓p�U���h?��.��A����k�ʯ�RG�mqry�9)`�[�o@hJ����bB���gO�H�T���:qeo��v��?��(��MgU:�m��1�V����нNz������&�f�hR�q"òS�LJ����"GN �X�Yx�8�c5�7}G�<~�O��>��+�$�
;������/"�q�dK�s\ߊ@��x�Z�_���;�q_\fο5��M��J��}j���)��N@`� Й��ޮЕ��'�O��vo��T����?��*g�8�ྼu�_������v�	�")�E��L���o�@�k�ΨS�2K�K����/!s�C�'o�肅ﰔ柤q�Eb���R-wr$5M�4����W�I�ؒ��:6�9�mRSRZ]ƃr%�ias!�7��+�������R��E���Z�U��om�P*��q����g�������:?�,K}#(�w@c��VZ�S��@T�ϧ���c�隑հl�Dӆ+Xl���婀����Lm_�|*0d�+��yu/�M��R�^�Ȩ9�\Yy�K8,�T>v���G�����x�:D����O<��u��<�]4��#� "5��*(��IK	��K�O�^�bFWk�Q���Ný�Y�O4�ʝ��F���w m��sq��J�An����CoD�7��ʍ@5�hA�2�����͒1��m�����&Z!�ĪFLy ��Sd�<;t7Qq��%e���\��3��n��Ο/�����KEiQ��<x}�z�K�y5�v�/3�gq��D�,UV���s������K�O�#U�|ޗg���n ��_������I�� ��!eӒ徃�(�[�XR�t����~C�ʂQ�N��'�W����F(�˘�Fۦ|��=�2M�	'�%��~�������;s�t�y����(@;����=�/	��*�16���'Y�7�4�U�	���x<���o�(�1���+�.���7ڹ���n���k�*�R�=�bg��$���fX,Ht6t��G�+�͆�)���6�AhI9 ��_h�����J��XIZytķ�3U�՜{�xi���D��ܣ-:�'�˂�M;覜�.�dx������Iw�}��R�����|
l��P���)��*A�6�����B�Nzo�kQ�)<Z��P�Jl�:��R[z��]�qV˪֒W
U�"bI���=�����\��n��d񛨿	ξ��4q�5B=+܌��-���AN:Ǌ�Z�wS2S$��I�Qpg��&K�-��{cNm:��#̈�۠_��|M+��0U�e6"��A`�q=�Ϻ��g�����M��|L�ˏ�*��@?��n��y�(ͽs"�U���ڟ��D���$D��t!��kJf���Ku\�D�,�
���a�=`b�.�Wi�D	�}G)!ym�����\��g�LO�l�g�7��4EXM,#1rȿ��C☗v��|�:lJ������aN�k?�V�B�m4c�����󉐳eq�D���J^�a��u�O��F����1r^�:�4�Z����&E[�\�#p�,{��|���O�X!�A`=�5������#�H���%�:TW�����O(����\iۍ_;�u�h��m�1�t{镫��`ߪ������yٽw�+�{6��:�]!�E����
ı4r�����������US�.�\M�Z��Ђ-yH��%<�":98E�*5R�ib2X�=���Z���p[H�d3��8�sQD�t+��>�ظgg��@�H��0A��;���������l;n��?uh�4��y�}L?�&i�@&D�Wr��粥�1���ql��ҩ�Z���Z::,+��倅N��
�iDi�d7�qI���i�<��(�u)�'��>k���\׋�d*�Ղj�p�׫[9�����2>J�	v��be摵���t��4�\޾���)�I�	���=�u�(��i|O��;����ױ�~�X�Q�+Cc;�Lo���{L�X����g����Pe�+5��I���[h��h&��V��5s?�[�:De��a�W�$9�2�r��_KϪ���5��&����[�Qs�9�a���<�@�B�d�ɜkL��9T�	M;h"K)��-ǘ��_�%5��i`l��ˊ�����!/�r����o$�	�y��^�00yb�ⷱ�(r����&2,��#ږ�$��� ���l��g����9{*k�0ȴ�-��o���G�2���Ɏ�1��o1��i��<�}k�p�6j�+[o�h��f��T��Ll���e�2��K��}p/�az��4q��/�X�i�{�g������ �\�����G� 2��:P�Da&Ԧ$���N��%NKbw�mr���,e��w�)U�GL��OC��=�L�[�c�8t�����f	PM��kX���*F��4�lj�m8���vC�����8�vo|�,X�Us@�W�t��D��`b��ш~��>a�5ue�-�h��X�Q��0�x6�$�L���Lm*]<4�ϨyϦN�tቱ�K�`���}�|�ؚu"^x�~�: O���9S����V`c0W=�)ˊ�Q���#L��3�8X{fL�����w�k�O%���6�J�%9�E-���l�Z���E!>RZ��d &��Kŕax�G�9�1�ٛ�>����<��P �R�;�������V槯QuȒ(��.�}��Ǫ���/'��z�k�Cٕ`����?!8�������o��T��1b��oW'N�-�d�J���b�=NE�cWd�Fp�-���G&�:(�fɻ0R�� q�qx_�<	IY�ekhR:
��a����8�G���zib�#���}ʥ�����+�Å���6<e��ߴac����Ht��/;�w��F���x<�o\	�af�#=��J[�1�a��C|��<q��ڛ
�{�*��;�3����,i����R�G2�<�Q�	����h#p�ޛPS�o�0��m.�O���a��
���#;�T����M��?��6M���߻OpG����Ձ��݀�:0Q��r̼�tf�mqf���Atׁ�\�FY���̹B�?�Z'�6D(���kXn�}�~�Ԓ���i�Hߠ�:��b���jL��tg����p\(��?���_�l-B/h��T���R����M�+����w���>x����3_�v�Ϡ�[Iv:�6+=����@�<.N�FOXQ�IAWe���2�8�[>���\�uH�R��3%�N���1^��c�_ݦ�Ga3K�I�����^������qnr��̐F��R��v�ے_E�#�E�qNtݯ���8���*8�8&5:�F�Sя̪7�7·o��Gr>Exl���F���)U �8�*���v�hvPH5v	M��$L�6S�sye��[j.��#��Q^����o�J����d&�A����U�*c"@��-?�Yu�^�����&��	0@�E$s{���� f�tͅJ��_�1f:f�R��^ЎB�di0�Z7Sfu����y�����R�EAy��?!�Kf���ψ���F�4����`aRޓ/�Θ�z�s:�=�Q�0�24�Y<�r�$�Zs�c�C�a���é�5���8�x�`�<�$��Y�L_'� �����`?�%�Y�Cb_N_���rD�S�pb�^N!8��� <'YZa݃H�ɼ#�q��N�!+�'�c:���D�6a6���)��=���g�^��[w��3f�"Oޤ���:�"s��4j_��I��m��aɦ��N�~ز?}��t��F[���r(UBckl�ܯ]�Ż�(T' S`7�ᦲn2fEO�e��-3"��~@� HbjP$���{-�ޟ��[�d,2�/��n����X��P���6[��F�E3	vV����}���"ʧ�ܽ��wYb*G1`� Pi:HI�!��$C�S���� ��=�%s|�9��>�m����A��d<V?SU������Kx��O4ìwb-j���0�M��J���{�����zl�Ŗ�~�h������o'�%�j.I{`�e9W�bW%�ݤ,:��j�!�D_�H�J���V����*dJ�*���Gq��*q+bILI�cj�;%°h�ce��4�hډS����L��],(���.n!�P�jM�[*5Y��n��m��-'���%�6.�����1�֞���|q�V��Wb�3��<�92��qOx�1�6�&�ct`�$Wgw������X�d��W��n	��^�9�/���!��|#-+12�0�a?/P�W���jd ~�˜��L¯V$��jAL��z{������l|?)�_�ɴ�$(���2n��JWq���S���%N�0"��}f�A~���9%�z���ٟ��u�����ا�4��G�N��ZŔZ�Ҹ���!����!`Χ�*,����qed%�6��z�n����#rBN5XaU���B��{�5~��y,�� ҭVh�_G|��0�[eS���Q;�CX��3[�P�c�6�{�Sc @�l�Q-�h��=X�6�⬵�U��P0u�=�����giug�x��Y�����#�>�j&㱸�>��'V�:$#���+�̹S9�VC�j�Y	Su#|x����רW(�6�0ǭv���Ԙ;ہ����7�b}����7�l_(�?�xG�j��ɽi��B@ޫDp����S���I����T��ꝟ ��(�ɍs�����Z�������<���7O�;+�SZƘ��t�{��[.�hxL�MFh�MC=�aަ.����D��yt#fV���y�W��}|ds��S���6�@�����Ph|�x
f�z"�:&9-*YUyw�%���i�����I���foiJr�B�ޒ/b]� �@)�\��qX5?l�* �$&X���&������������zu״ܣ�h������vd�V���?	Ճ�K�¬�8  }b��&R �I����\J�X�$��q6B��oJPV�O:��K<��2��k]s�|��|���zkL�@+R
1@�螾fx;rA������0��s�|���[ѧ&��m@�3��?�Z�������k!����R�U�`;|Oh䄩�#�*�?��ҡ�c��Q�(9�-˳����Wc�S�4��O>�!�mg�ګƜ>¨n�-M)�`I"���Q �'�شd����~[x�J\��ҏ}��EM�z�ԗЪ
�s�H[36b��D�y�"��CϝBP�G-s:�I�m&C��m8��9�g�tq�C](,GA��/v��(��|��Qϓ�U��x���6-1J�����<�M8����������?B/�[�>�@4DJ���a�5g�D�v^^{��O�=�V��:�r�Kd�%�02��ޞ�f��B��c`F%����ܦ�:�t��	��!�X,�s����o*�YP����H�s�?W�<4)�Մ'�������D��L9����
\'�A���9?)��UOl���|�- _9XO���	�����JG�������R����ߤ���_��w�w3Zk2w�z����:7>y/���-j��>R������e�=���p�TJ����- �8�Q��o����9�������$5I}� �*\�oE��.��.хڗ��I�e��|aH��r2��9�*�6a��� �� PŴ�G�>]}n���O�h>�8���i��I�g0Pv\q��:,�>��9����+w�Ox�i{=)o�A�z�!+�������I��]�;`�O0�]T�����)E/���%�����,���h��M>��]���F� ���������z�$�|m�_o��,��"���xݝG�<�}�-e��h������Bf��>YY�47�N�7F��6]����
�6��'�;O?|u7P��,� �!C^���jɲO$�����t�����@�T#����C��Zv��6�?_vj���o$r��yY֨fuw-=$��@x&�E˔������	X��w>�ϙ���t@ԗW��.ȿ�TLH��q,(�ǭ0�
���f�۝�'��pgV�:/[�$�_BT��sqj\�j�H6����!k)�L{!��(F����,��[�� V�\A�<�\#��ZhȮ�.�uk�C&j�߮���\ V�.N~�3JJ(P՜���N�u�R���O�ZU��Z}q��	����&��V�pٚ����䅬&Ƀ����&з��g,��8i��z�����@3�\F94<٫�2kլ�[��t���*(z�;�8�6���Q�^m�S"��M��;�彉�����A�5�$��Qކ7^/�X/��r�k(�я�lzy�t�}S7�$H�_4��S4)6�����u��e�1��jk?�q����:� ��M�&��b;��ȵi��gm�UZ 8/4����b����@����T?��Y���'�4p����[�%pt���f�9D}Պ�wi6l��)/g��j�dh�M��J�����n�b_h��orņ��C@$�⡦q���C��Q;t�W�ݎ�}�X�8��!��|��%#�"��`#$�`�	!�������ɛ��9ʗ��t����&8�y��P �(�K$P��t�R_2���;)ƭ��~`�L�}�i+N����������'y��"�.−��R�Ҡ�ǌ�Q���/lb� f|u��~����:�o)d�"Z����bh! =8x
�Qeo�������1��)���.B1퍡� 
3]?,��?��}���Ƭ$><���Η nsژs�pm��t�d���\J���pWZ�������a�Ƶ/��\C�/V�1�� ��<�����J�xt�N�����@׵!�bˮ�����R�ՌE.%X>�gw'~����bb��JLDEq��1Z�x�9������_f���ehN�4����sl>�Ӄ���2�qH9ĕ��� E+^N�y��u�Z���X�ب��7�m��p�a�8�q����Z�����l���Wv���/t|�#_$����^�yo<�h&��sȥ�K���g�C,����MX*��Hj���'M+�3@|���+��h :�H�3N�<�՝��zy���*����)�[���`�U��rE+��dp�݊�{s�����y����8,�a	��F	�v�:j+)�� �?.h�D�H������_e)�R�?8OpV��'����h�B'�ۘ`Y��'	�'JņU�"MQ��=C!��l`.V��fb&-��)#�&8%���4*���y�G�3�1~~Y#F�sL��SIBD�����6�E�m=�Y������j�❝4��5���E!ٸm4�F��^���N�6��ܦ�w,�c�̼n7�h3��IA�
��oVD9�y�~�HEqũ�a?�6I]�ލ�>�g�Z�����B�2��e�?b$����M�V��^YM���� ]�46����8��W��;Q\�T��W���3:�OuP=�����\^w�D@޿��v�q ��$C_�u�'9[U�3�o�&�k{����0F�����0e���oWˏ�TY���9b�����0m�sK|`�1�.[R�㱥�N,"^��1��zɣ��lԢ��@�Im~swf���֠�A������zki�ݞ돧�Z��T�O��to�f�����G|S$~��z�@���t~�ں�n��r�;=���4m�n��,�~6��~[�.��rz~J�$c�
g�(E?-�fL�A�W/��,;P	����1��{ 7�3�(g�����r���Ίb�Gk����H�vO�h����q%��z��X�{ee!ޣ�_�V��te����6���6f������M�������|)�AV�J�N_�A���+!7��B�CdDc�0߼�o�������I�`�?���-�ޚ>g����4b��V������".��6�)=��]_��1��!���N���]�k�H����&�cG�&��r�M����3�k�1��(��ª��Z��]RG��s���{Ca��.{��d�WY� �(��1�mB��J\�\p��v�W��92F|�Ԃ�,W�[T�>�0���<�Ȏ�pX���(�C�(�_��6��^Ά�1QȶK� �ЁF���S�n�]�Һ�Q�sb�Q��}�P֐�*��qM�^�ɘ��EO*�>Ss�jF��#��B[?�F)�󲆎w�υ�0�7ٍ�<>�&�xG28����T��A�!{
�¡z� %~�n�������m#�y{� ���4^DϢ���)�Y�-39T��"���dB�L�J2>߾SwLoU��a�Dd�����H��`N�v���bu/=ߠ�W[^�[�q�j��%��{k+[h�TR�b;��&O�������"�pU� z��]oz'+�l��c8��[P+[^\�*"o�5r��o	茏���.�U�������� ��[;�\O�������*�~쇆*Ĭ��3ѩ":Ԥ��]3��#���V'l��=`�#��Gp����aEQ�S�A,w&��{t@H���P'��*KtBM],#�wa�ܨ�B}@�6C��KX��)�}L��]��G�h˅�ף��ɡ=i��p#�0c��;Oz��{�g*��qt�7�5k7�Y���Ś��#x�d_��h�QuL9q;?/ҩm�w)�鎗�-��q3��2��*Wx�fG�'nV �e�W��Z��C�|a��۳��7�ޫ��(��:� ���|`I�v~�CԋS `��3�#��^ս%�*�|xy���s٬�U$M_�;)�3TQ���W�������v��0�pۮU8�b�n��t�]�ՐG~h�	�r�����;ւd���Y�Ѓ@�"���C���Om`za|���*�`(�(�?�u���]!�P�/ 9��b|Qq�D�)�)��+֚hO���t�H�a�
"鎮^Y�x5	��WQXIh`��겅$O��x�͹��Xo���.�Z��S��k�2(Km�����?�=�ŝj��v5z<�Q�Ƨ	p�OҀn�"^w͋8�&�M|��a$3g��
�n@��p�,F� <n�T�4x���SƊ�L^#�q��t� c:�\DT�Q�N��6�d0�8�l@Q��[h�ό4ݫ�}cz�q�$r���8��JP.2�ە�ޙ������)��Y���}4�2Ω��̔��?��T��"!oFg��ko[r!����DWe�?XO&�Ñ�Z���<ҳ:�"j�$.�mAqp	Ϻ����{<T��� q���8~o��n�����핹�S���:���i�<��� z�N�Mۖo	��{b�C/��7�]�ְK=+�%��<@p+��������c��� 3܎�ũ(�JN��d�v�E'�vt�5ޝ� ��"e���9Ý�)��%Z;��Z����i�+�<�љ�c$�Q>�������~bX�g���<�92F�Z�F�,��N�%	&��X�ɽ�>܄I�e����--otm>a0pH��l_�-Q�0"rf��w��?�\���b���_#���<���v�@d��V7��O�a�e��������=�(�;�܂2Nc@�<�� %���i{�V�$��w� d�˱S����6t��H|�����qD]j���.�]y���|}#f_�[�}=1s^����JE��tK�!��+��<�gۏ�����g��j�ⴲ��1��n{Td���A�;o�Pv�s�������?�6u�T�[W\__.��*�Ȟ������-q�t�0��b��N�V����/��{�(�,
�j�V�S��T��?�)������n�mO�e�j2�6||�$��S3�)E������,���0�۲ޓ��[��s����-��<����z��ЅJd�[t*�E��#��Dԉ߅��=�d2:ҳJ��Ӓ3�]rЛpyX���Cvp��p�IO	R��UIY�(�u/n>u(�+FY6����VG��2��w$�o�T3PX�oAq������f'8��ώ��?�آzn=�!!�b�p�G<O���A�[�N䶝%L�rJ��h"6���2�!m��Ħ3���{3n��;���S��Vg<ۖ�I���ʊ���#M��G�RL�%D5��e$�GVF	뿗���bN\\��W�v�p� �K?&���N�ZXywA�\�#�X6�Vp�|�������0K�bJ�XR��6fso�S��,/��[�7X��W�3�+�nurB���" t�{�K�����i�.c��Ŭ���F���b���8쮳�*���,���~��|��P��
����XB�0�)�����1�|����3�J�Ͱ��8�F7(�`����-�{m���	ѿ��B��D����|�Y��?/շ�ֻ8����ծ����)A�9�M��%Tw$[e�ӡܽ4��S�H��e�]������fyRn��SF�,�X����7�*�%�����,;"������+�r�f�D9��R͋�N���(��u����4���I�Ưp{@�BP��f��<C��L����%_O�4ZH����HĢ/�g��Ҵ�r[���"�(.&2 �a�\��Qq;��a�7C�ԡ+�&��# � �����H��EoI> ���
�̐�~���/�.s��'{E]�Ƕ��<iy����^-��?m&?n���H>��]jѶ�,�s*o3�UB�������2�X�A0�g���,#YZ�Ax�҉�a��V�=)��L��.��
;5	�+ ��Mx0h�w�u��yJ���K��T��EH�hA�7���^c7�&p��%T�n���[��Tӝ�����3�9��Z��Y����/Z�=�YA��"�Ⱥ�.���2��}vG�a(���j�/��[�K�P��@�*�P9?� Y�/<.��9r���8���l&B����*rl#�x�E0�l$M��JĮML�G����cWb���G6΁�p& ��ui�g�f�!�Cv�k[����z2�7�e�cc�m�O���,}��B)n��{'�X)H���>�@.|�&NY��esD��U�%���fK�K��k�Nmx@�;�b���e�]S�/2(��P�JH����/һ��o�j���6S+r�<<<�5~2.�9>�5�%P�a��Ԩ ��-��'�x����������&ͳI�߀'�8����q�1Хb��]J���#EIhSho`��cc1n&}�0}���Ò�`�b$�N�����_�7V�^t�t�B0��yHm+����'��3���Y�V��[�ֶ�ՙO7n��c;{��:)�{Š!S"�7t��geI��p&��*gvT'.:"�\Ǉ�IނѝFk����ྎ������N�̤l _0��W`�-v�� �W���#�������-l�G»�i�s�e����G��Q�G���#��_I��?�G������/?ލh��r�2��Ռ�8�LO����Պ\��eR�d������4�&�����:b��Lf�ߣ��X�3ho��O�?ч�S��p�۷d4/�*�k$�ɴL$6�	����4�~p@��5"�ȹ|0�ջ$_�}n��3����7C��d�L}B�gE��N�;�*����;?ŷ|���L~���o���"�c��b��^�5\Z�?�H%��*~�rĜ���!��w�{vY?u���P��>���r�j̪͜��y�v��Wg(GG�K�Fh-`��U�<��n{�	 �0�s��E��I�d�k�D��S��f��.?��ǭ�H
܁P�r�d��c�Ң��*�$�ۨ�Ő�8���	��#gBG��sB��GMI.K�h���M��!N�}'� kI!�/[���c�^�b�E7�,�X�.� b�'yar]�d0u7--�~�(m�u�_r�-!��$TW��9�1�yqQԩ;��� ә�0)�WM!