��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�����3܇�g�x��to��F��Ɲ�e��5������c!�^�D��+dzb�t9P�������e@:���|�i��z�pu1�}s��J\��;����of�C�iTw��=�����H��W�t��5�I&kkm�|����q�{(ݵzP�Ů���\kBk�w޶P���-�^O!/�ef����ġ}0S�o����=b��~�N��b�V�|��@ZɄBb�R��}�����!����w�ֈn�W*��C,��G����&C��|2�i��au�ģo82�ٛ8�G,�ԖoCs����y��u ������ۥO�Zd.4��ha�h@R�rI��vz J%�vo�Ի�A��%��{9v�з����
 _1*�[Os��eگ��w�*��*����>.�����G��<��6@�^Q�K,4�A�X�<�����ن�ؐ;�8lD<��%t^������Cܮ�ƗS���Ucvf�Nv��Z��3�I��3�"F`�ĺ�aP�W��6���7<���![I��Z���C��x��X#0A��/�|b\{��7��=.j &��r�Rh��.%��O��9��*��X�R���|"��SU�ӄXpv�	�H��K$zJ� 	[I�������U�p2KcL�O+"2����v�WyP��Oư��܌��"���B��LK�ǣ7���ax2��f��
��iL,��AR�O�u���7�tC��u1��t�	���J51C���,6�:������,"��#�֪%�~]�|�� �U���3j${��Q��ۑ_�>��9'���cCi�T�R���:uso �\ ��@"i��L�͗t�&�7������O^S���梺��������ljLr�����^�>����Ť�R���lɕ��f!d��N.��f�,=�qTonp�嚈T�u��?b��m�$`Xk��O�����7����3oSAq�9-�ͯ�@X)�q�ِ�.�b�ĥka0$�P�C>A.\��A8������2?x����Sgɸ�UGDTA��	%���"ي�m6����d1�#�c��������9�(
�6	�EU�l���__��oʧ/��7	7!�H���Tּ����� C�>�)��
 �#>H� �ǣ��P��l�!�ɵG��1��Hؼ��*��Mp;�"o��] ��j*����i�����H3���G�
�e����`9��%�I��ӿ͈,�X�u���X\����n�{K���ʡ�K�O��y��FuZ�&&9���02��D���9��o�&�'-3k�*���Է��"Y�+K��Mt�� �Ѵ3PI�1��.=؊x/����Z_-r��(m���3���1s���X�}�窇νf.�I�2m�P��ֆ^����ҳW�Iļ���w�2EA<]@{~צ>�0�n�5i�9��;�G�~�@4>M}c:���`Q���mZ1}`�p ���`*�}Wo�I�`+s>���z�����P[�� �s��w�5�{�\\�e�3��������MOc��Jw !�H����0��oB���-�d^�����ir;¯Ǐ�6�3/xD������mM3��a����Q���4znx�n�k�5=���f��[L�&��@L�z��<�N�߅���+ܧ�hH�>3� �Q��s`��Ն�sW'%�T��cDǇSA���`\�q�"�A���.䐒�T+���E�}�}Ԟ-�d �����+E֗�ow���M�['u�>5��fe�N��^p��y�:a�:��䘷l/�dP��*3I�HU?�]�.���(y�H�!͡�t������eށ�i߻yN��
^���� �@��������Q�ޅz��	@"TE�]9K����,�_�E��"}fqm ���l# ���69O����6����wF�x&YY�_e�k�sŏ� ���8ĳK?���{�ú�!7�~c�-5�����C))C�-�K� �[d�;*�,��<s��ax���4ڳ�$Yc��-�-��=�Y��� GZ�5��!攄g9�Ł�<0��%N��؍��!��|I���ZS�ѭT1������΁� ���B�56�`��{�mLv|�̞��E��cT�bq�������{��c)K���/���C%�*��C^?�?�p�P�u��EBS�\�@��b;�?e��7�@�@^��t�ֺZ��Y���Yr�5:2lY��CL���'*�K�]-d+�{����$*	Yy��#n�dR$DS�B�t�ƹD��\���3NF�����Ƅ�>�%����Ľ��?hc�W�P�HPk5Ҿ�)��Jg^������`O�cZ�C��T�D�ҩ�3��t��X�����8��4�$�Wo�>�����r4H��궥畲��L���y�aY��K��ZvWBo�?���ԋ��.�C��X(��C*�Ou�R�i^�C���y|�h7S�J䏤Nz����m���Ճ��1����l�/^I�i�yJB�H��=EJUM����77���i�����������{�`	ӣ� _^��<�RS����^�xq4>��3���/��Anz�I�$�f�9g�Fc-���Al�}yWԾ�)$�V�ۑ�V5�0�|�(4��+��$ЈX)H�(ll���DӦ�9�2��`��y����혙e�N `� aK���lA7E��#��0Cv=g�<yo[oM���ȥ�%��1���1 ?4b^�5׫��dIYY&u�7C�>QζB'��j�'2��9�hͣ��G��C�`�H	��W4'����>�%����Y�R
���:
~>L��Ԉ�65��^��+����vDgP�IO��G4�9���B�闓�-8Y]v(�f�I���v6@�ι�Y�~Lu���X?���w=���li�sU��7j�uK6�^��$u����Na0��D��rǢ0A旳(�+��Af�M��jK���C�`���*�r�����]��_fI߬5ё�W�S[�ThI��5�&�^����\�0)Q�m�$1��d/S�aF!'��8��ڼO�h+�wI�H��P�Q��<�鏿⒎��M:y�_<Mw��,���KE����<9�z���Hm������t1x�	�Lg����E,.���<Bq!�.U*>�3���AR�0�[���8�G������(��9�,�w�D��K:L�����=8�ϼ����@�y��+,�۷Z	��9.Ǭ����K;'OJ��y�_���eXIIz���Bx�=���6 ���`���>,�}���)�L����f���9 ��n6� �W��nl� ��4�����\y�I%IS�P�a3���N�ᢷii����,/1\#(`p�ʿӁX$c���}§�.�M�Ї2n��s�{�w��^�ˀɜ;��uc8	��Ʒ<�p��|3��<��ۮ�Ǘ�,��d��S11�_c���U�K@x���E�?�̤z���	w֪gw� �Jr�є;ĊY0Þ��Q@y�b�鸗D��e]�E��#>��*x̡9���ٟ��gp�oKT���'^K�8!q<tp�U���i2avóXiF.�q�d�zW�@���^QzV��q��a�0'�0\�!d�w+�;�YA��;��^�k��n]��_�$R�Vl��T<w��(s#�m��ʒv0����5�4'�a^���.�t�?�a��+WYG�1So���&	F���Җ�ֽ�}U���S����'�t4���3�B|�º
�sc��5���e�/`����wz��ߛ�������b�Z*ak�dnp�+��G�w!�&�a38�M��LG�bU���k��B>H���mG�o���ؖ������/jP>�JK�t׭=A�Xɢ�}�9��L%���Aצy��"0$a��|Ӂ�m��r0d�� ����Q�;���mF��k�!:��:���!d.��9�Fv�sSh	��qǇ��Ԡb�z�6��BS����@��]~\�?����;���SY`�|�'Ny��>q���
HXz�L��第{��f3�c�O;��;���J;VW�F�.����2j		�?.��U���,{,�S�#�֑u4
�H;�{X(�U�v-�6�\�}��xu��v𨨧9PMq�vV��u�EX����sNPIprG��D/���5���XJ����s>���G|����:��Q4�����6a{&`}��v�"-='���xG�!j;`G������:'�V6���,FWr�I��x�tu�e�y���G�
%���>K�J?`�y��m���n���H�L
�Bk|Ԍ��ŎRL�mVϟ-˞,�5�����<WA�r�ӣ����)T��\n�,�b����0X�(��˘ٵGu*��/a�a�}�ɰ�0�B��56%5�*�!�a�������PI��!r�������?�U�*zo�`qR/��)B�3/K�%F�d�u���%��f��	s��80�'W�W}`,���oo�@�؍�T�^k��̺�t?�aA ���g��+���RN0��9Q�#�UB��Oy*�҈B�(�=�'�8i��Y�i^2oTy���5�06%���z�#UL���pS���g	{A�ȅ)>�tn�l�8<;*s;.>D�:�K��p�SI��=�x�x�@��d#s��B�X��p��?��{؁�vf�H~ZZ!g��z<�5 ���k��vo��9���u��vJ ��DKZ4x��Y<R��6�7^2��N�~'ō���4��[��ʜÌ-��r���@����|5��L��aR(�������g��uoa^�bF[q3��7>���>�7i_
�U�m�젽9^��Z{������Q^{�ƭ���#�zd��,A9zip������d�8���˺F:��	Ԫ�H��=lx`{��cAg|k�c�LU:���~́&�/D�'���5�Ur����C5z���
�"`�nC�읐��P����-����}���W�n'��T���]��|f���K��"�b�T�!�%"ʴ��c�p�9k��Ӿ�@uwE����q��1�z��f/�I8 ��g�c�&XW���<r�(����FX�،!�*���`L�� �� �/Dp�cN}���J�l�d��&T���b�>ʔ��������g�՟���KD���2��M��Q��%�����~��?�kCk��
=J���˸�3�o�d4����zk�V������=�5ų'ޜ&�E�ۧ+b�u��X�M���H����?%����Pͬ��'�k`���c)�_zع�G#��ۯ�'
ɄG!RQ�`��JC�=�
����*��"^�[�}�n[U�'��i�H�fw�i|�ڢQ��������l��	+P0����S�	>;�ز����s�
�@ Y5��B�Mue2d�fv ����q"����C��(V�+���m�pS�`6{C�/��
�P?NiQv߉�Ƹf�s)vg���vj4��K���vD������i�y��B�? �vq�]����Ms۾��?'�����e)�?�Y��tM�@"����3�ɺ�
9��{�=D����|��(�J#�,ߙ�5��տ�]��o/ʳ��o�����䤥��*���!_cj�m�d�����/3@�#�߶]���^��U���H�0����g�RzN���݈�lY-;}�0���#�}��l�����N|H,R�l��QR�R�K���1��y�tbD�,���P"���f���|QP��ό��xT�����O,����o��M5�. ��UT��~�x�=���5o0���W(��%��ա=���򌔓Uf����J�;��ː�H���+&����:Z�廕W�Xe����1J�W�m�M�l�+�Nw��G{���EDz{%vf�ɋ��