��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O� ` ��h�����mO���ް�2D!F�_e�4�����#!�"J'�qL��p*�uy�:<�_��"F�D�!~�E2��C����_����o-�y�� @�Y)?����܂ʱG����ʒ�W��u+����@�b�U�p��������U�f�	��5���Mt_9��2p��h�8�z�J�"�&w��������ʭh�	�v���ku��i�ݺ�8�*yp�������8�փ��LQ�5q���4g�H����w�	�Ѹ�� ų�������������熖`��l�K(ҏ6��ޢVC�i��K9J�Ҭ萕ng�Sm��_
�Os$)�ˢ7TD�j�ܪ�dx�������w�`�?�4c�]E���y���9��LS|[r}FIAN�ܵ,���#aT��ےGU��2O��ƀ��(�%Z�%���$����KsN�Ƅ�B	N��F��̌��j�AY��6e��=Y��nςG�O|��'HafG�
�
=���k�k���ydC���|�h?uP��'�t�'��v ۰-I��\��PbC=3&�n�Qi���E�n�����yJ0�.K#�V_��V�> M�lA�L�7<*#����F_+���3ĥ�Lr��qr�����ZR�=	K3����2��.����{�����<�������k���l�~�^/K���$��zj��Z��0u'��!� ���Qq5k7�\R:%�.�ȑ�#�&���u��s�en�7\ q��,W���6�N�%�rC����^�3O�Ia����f�'�r�e�BUl�O ��ʰ����Ʀ�8k��'�c��=�aa����b�J@#  �����S�K� �����;�tY�4�����l�t�9��HB��wN�-��UW����_GՑ�6=�|d���{����+e����8n%
�kp�#�M�o~�}��2���焖	-�=7��M� *H	�4�?��9��+ҥ�T�9n��	<��k:�g%C4π%�>n$<���z'�ܖm؊�ٰ���/�o���߬EN ~@g���6��k���ƮHc����qn]���i Gg�Z�;�`+l/6��٘Y�Ű��;<��U�pw�����{�R\�����R��� ��� ��ԙ���MRϦ;��E�����)���+�Y�([�u/ch�J�;9����]������0b�%���n���{˜����ݝ��{�����^���L��