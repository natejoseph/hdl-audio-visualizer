��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�"��S�&h��Ă�����M���,�0,�KH��QG���S2ʩ���8�@/1Ҿ7�F���Bؠ3-q� �l��p�dB ����\�A�W�^����}[���[��P���T�ϼr�Mb��G�d�"_U�O����m�.��3��?�X��k������6V�L�����]��%�?�v$�j@�/���@,��{D��{�����(��z�B��uS��*�L�1��,f����[��׹��8:H�m�ЅMt�����������ZZ}~S�<�OS�H��uw*����0;���L��T@ �Y�+NC��ȭ8J����Vw��̒�K���A����@:���mki��p������&$�^d>(|��`��B��tqP|%�D?���q�����Q.�d2#��{��mw7�<��V� �B��H*�s�W���x�(� ���<Rj	w����?����&���:��Z+��ܠ�Mpk�
�hŨ�f.�M7X�y�!��7�{�q&BC-��2O�+���Ḋ!4�y7)�m�=S�i���֯�� ���>�Z��xv����o���!qC�g�v&���0��&���~l�'Ʀq��J��ݍ����Mǥ)ɛ�8�����j���k*,k>/�G�� �!�Y%�4�o����7q<�����!��[%{��|��9�y��Q���G*���6�\�Y�����@O	�%�Z��JQ�r��G�N+�T���B���u��g2\�
�v��]TJ|Q��E�y�G	c�J�<	������G��Ȳ��ph&��/��c77N��~<�\x�I��vy��}hH� '��3�f	���A�Ѻ*���2 �:a*|�?ߒ�şmɐ<Q_�:�{�\N��?�'��1��,vJ�����9�����+�ZN*.�����(�%q�6M&7n>���/}��V�O��'h��T��W��3�^J-���c��y�Wկ$���y7�rz�����L
 y�,l!�̧y�t��泯�+v�}����3��uUv~ۻ�׶��x�k�p���`�X�H�W�G�A#��O�7�KR�ui\�T>a�F��ٔv�P�>��#���0�4�����Rτ63m~��J�T��ۚG߈ų�!y�x�wm���#e�}Vj'�B�����A"����8��eW�ձiLu��8��x�Z��.|)�:�`��6��9��&Ey_Ĭ���,@m�@؄�򄆁��O%���B�ktӂ׫.�����I�#�Y�'f�o�B4
�F%��2!�rv���yC!(Sܵ������H���3��ex�?jj	�C{���R.!G%Y�1ؗ8q��h�f�uT����OY�:i�Oh�yQ�ٚ�q�\(��U��6�>��T���LH_[PT�@��J4J�I��秝���+�6m���r�EߠL��(X����ˋ�.f���h��K8���I��Wht��Ţ��J�Z6*4�0&�T��=�[���>ᢽQ��P1_
�eU�y����ɽ&x��z�0V[��5�z_� ���iH� �v�G�9��`D.����P���8}7n2����6k`��)ϙ��E8�_$4�H��a�w"�CA<����p��h 
˥\�swڢ�5}s�>���Yy�3;/Q֞9���/P�'�����4/��D�}r5��hb�D��z��@��"`��y�*A�"/9��o����7^��nFN
�]���8�V�����}��f�	t}�E1�H�I�sB���_	TC-~����9���I�����v4L�9���zAD�&\�|����r��ڎ�#;RKW��D�U�J��c���c�8-���K�k���H*]J�����R�>��:��v Ս��	;z��N7�$��v��n".%��W���H��"�g�E�zB�_��7u7�R�M��M��&t~�h�(U�g�%�o27��>����:�ɌۧR��^�I;����e@���:Rf�O�^��:f�����bO��P�{����]���r�	G���W���'�68�A.IWR�F���"
��b�)��@�ݓc���4�I6�]� ��Y�v��9I�`�����}:�����u��@i���������5]/���!��M+)���S|�����)��Xr�%�r.���vN�.�<z��A�:jMp�[�,:��:�(\�j�_N�����z�K/�v��Et���?�,
t��
��? 5c1��,$X�J\\=Z��Sd��ln�y20���f ��lﳊ������/��)�"؊���9���/.yg��/mʄu�W�œ\���������ڱp3Շ�r��K�������N�gHw�-�T�R_��z�\�]PVd�m���>X���Ԭ);���I� (�m�o�i��
@aR%��o�P8�F��u�S6���U�#yВ�t����\�D_ř�ᝆ�w�í���d�<�+���ǧ��]�)pp̉�]�
���f.�F	�!.ך(��Τ�;��ky����i?P �п�}���1��Q� �Hc�Z_�_���~�qc>�7y�BH��g K�Q&n�S�߶a:�oV!���a�NY���w�z4�ֳ	��K/Y�z�/�i�>��C�
N{l&�:��*��\��߃�V&��&"�"�lh�OWŝ��D�u��$��M�.y�cw���B"B���2�4P�8ĉM��W��a�����!p�_o�w���!y V�'�GR_�M[�� [a��2�b,֎kK��EpN���b�П�c�*z���n�ρ2��.cc]|��m����h�xSa�!׏w<-��r��+
�$�.rS��ct��}���P�E�|0�G=�u���w��6��qY�W��U�\&	����ͥ0H���k�#ۚ�Wu�ٖwd�j�g5�<����� [f�Pp�P_S��1��RŞ�#��ʍ�S5����	��ߴ�9�pof����7)T�x��b�x����y�cZ����K�C::�z�Q,����?+��w������C:��e~t��M�p�U�'֠�{kѳAs�^�h:KX�`5������D�zr�/C�xƅ��:���#;H�*�m�V!�J�V��������I�e{r��%��p��RU�#Ԯ0f����?�Gt@C􈞃."D�
���)�N�av֑����}Ͷ8)q?�P�\���̚��[{�Y���9��3Mo�9���8p�
j�K�������]=�3?��Xn�e����5
5����5�-���>vݡ�'���3�w�C�֏C�Ҿ���8\�Ӆ7�0�FS�O ����ۦ�KJ/m�gÃpJ����(��Q���pf���'�2ح���/\�nC���˄��qk�a 4�W6�c^�nP�!�x��IEƤ�1�:���ɣþ����	(L���QG8C��s/eh^�]�4���߬/�l�������q���t�{M:%��l���>���q?�c�ҹ,�`5�$��Y�y�x2��PD:Sꃪ+O���:�,�W�	���_ꨲ�S��Aign ���|���E?���^9	�l���&���s���'^�l�Ă8�r�>Q�b'�ԗ<���B#���t�f���l�a ��&�P �7E�����dy�2���/�w����[:<�h����ӅZ�|?�\��Q�=�c�8�>���8R�k�lZ�&�gj$����t�O�/	C3�y�����j����=H��o\/?�l+��_��D��,�Sb!�7�#��(�(׭<�c�Ŋ��e�:
� p>.s����ǫQ1m��,�!#���I�g����--h�e	U�(
�1��$w�t6�NQU��� �;}�+7���Az�7�i��Z��Z7(;Vr'� �Gi ��LeO����4����+�^;�h#	�����o��*g�BH����r����\������S��ɷK\�b�����X�d��+L�0�;��c�U���WM���2"�����Xpo'gx��v��#~+��F�[��d@��yx�I8��;݋��Z��>HC��d�;�P�T��kF]B�ʅ�"�*�ܧ�d�п9�8��&uv�U��{p�{���D�V~�%�LE����AYʿ �][���Y��ţ��f�>���Y�O3`5S<��M�����T`�R�o[U ���sRP�#����O��èBr�I���U�^�=t��9����1b*�Y��X8e-N8�t����`��� �u�٩���f��I��+&�	��4�Z����|�aH�����
�g��]-���qgz<�L�F�"qϯ�)�a����3����?6�͍�=�T�Bx@��T�_dOD��f�2G#�Ļ�[YïBw��4`HXWc�oy�IW��`����k���b�g��|�Qa�"���`��}���s#�� ��mX��ֻ�Q:X: ߈�r�c��D�(Xu�.�m�;df:k�h�V�j=,�Rk�����)[`��X,���_��*�i;���g	j�ଲ^���N����Ok�>�����Oρ���k�kS÷D������u T!+z]�\x��Ҡ��pw�_2�p���1�m�6�1�c�ߥF�r(E��PX��3D�j;6m�����݀ժ��H��H�?�H������1��p(�Ի
˴�;l���ng� ����m��'�~��V�'m��v�,��KRB4���Z�_s3�}��,�p�a�F�ht��	*��������&-�B[�#�6*\���1u��D��┞���6���٘��$��Õ�w,��?�`?��j�� I#�[��#���얞-m����;2"��i2��:1��7�O�`������Br*�j�sczh�T+_Ր�Uw�!�E)яA�R���~�<뻨�xr�&�%W����\q�!ʒq:q��eE���J��^x>>��G�&^z�{eY�$�'Ϙ���۵ZC�B�.���g�:��=3�>�8U�.�8��-�'�v�����9�*�`���8��X�����3�<��H;�ԒF�O_�Q���5'|>��?�P�m8�9����^)�v�������)H3}]V/m��)+�S^�(Cx
��A���������W7��bh:��Y���9���JY�χ:�\��j��/�V�F�}�F��<����%�m����C&�"?*�鵤��q�>��s��TΣ��!!���.ҭ���#�S�%������nοB�����ʚ�E�-���w�� G����ь�c�N����l��[2�_���mzA�}�{+ft�&���Ru*��]6��Z�cj)�S���� i����e�S���_w�.|�T����R�+O�~�͇�vU�ɵ'8�ɴ���'��x��"�9�l�҆�-کی;���cd)���ؾkm����>=�{k��w�/��p"�B=c��z�-�8��>j�A5��, �a��wۑC��Ԛ�ʚr�+�3+�kX9R�o�A�#[I"��G�3�����	Izmz��- T���@3��-�] �rf)�(���"C�#zFy'ң���x�@R��A�4�[c�����=�
�ό��P�������HI���B[�ī�>^����M������E��+7���x�m^*Qط�t.D�wS6�`1s`eMM��$�w 0��R�!�A�KUGɉŋ����:y�E�� ��h�����v�Y��A�	�
h
�6���(xl�1⹵�����DJ���
���3^��Rj�Zʇ����n�)ra��r���̋؟�9�ƍmod1�DTz��F��(m�H<�f!Sm��v�E7ŐGw�n�s\H��k%h?>� �1A�Rt7Ï�{��A�r�G�2F:o4����
�ٛ6��Cc#�Y:[?�}9�'0bܜ�A�:a����ߟ�S�ꩁ��F��0o1�������(��j��{�k^����l�^��[��vF�!Uk�ɅI���V����}���w��:�f!����d6�!O]j2
�W!�yP�ՔrD^�%Z7�0ڛ�]�d�w���bwA�	vuhy9�2�2@1ݧ�!��r�o��_�bJ�*E����v�E�J?/���-Bɛ���9f,���h��ߙ������(��˨]b��9��9g��r�����9�
��,���1W����RS��=��aYN��R���Q6i �:J�G�ˣ
-q�@+�5E�[�[s��u(���{��(W<���%S��-�Xk�x��7�p�ɬ�R��Yc��1�����r�S�-�{�?nP&l��:�w�m��|MI��.J>�K�����'��zs��j��]���#C>\(2p�����Ȱ���q8s�
���"�*�[��V
��i\o�� MB�n��gNad����8PҰn����*"ӧ��k�qm{p��0fe8��0��cȋ�s2Q-|��&���մdrM�
�K��<��=D�hW�C�o� =��t��x��w9�jB%=�`��M`��N!�{0��#��n�
�t��a.��hv��%KsG�6bA��uTL/�M�qǓ�|�VD}<�Ny�m�Jp��֚]٦�%-/ɭ�j���uF��MknDZ����o��s�߆�#�a��&��68p��]Z��8��9Ug<�P;�K��l;���Z�T]����.ѿ"�p%%*i����.���,���/(�J����2����T�{�i��څ����;$@H<�D��.�Sb�ZPΡy��YP�g/ʒ�>�D�?i�vUö8�1�=�����3�,�%�/�8��گx�py�"l5:�z	�d��A)�Ȅ��:��Uh������`%4�uT&�.n��)���e���)�`+�(si��g�V��lP:�:��Hr�Dz�;�"xSm@�����|��J��*���j�ٯ�EV��I�()�I'�"a�o]+��^ep ���3PIl��.��$)M+q��aכ۠���Pi��]a�83��ox��1#�=��S����4�*C�8,?��b��2��==Y�-!��L̾f��"��4U���aY�8=+w��L�(;Sb�)�c�FG�4_�7Q��sqM��j�(yV55=�P��ij�=�s��EQξ�4�!]aؿܣo�#�ZF-��ϋ=F9z�m��^#q�/�hڪ����'����Oxr֖�ty`��q�p���{Q:	���A^�E΀v��*�C��Șe3a��d�r�2���"0��JN��b��PB���u������,�b�{@���W��hb�6�}�ЧJu�,����$�p�?bhUZr���h���.a��Tz6kү�(Z���5���GW�6��X��Z�P}���	���G��D�eꭸQB�t�˲z ��]@���S�O)o�9n�9�W2��10 T�Q�,��c>b4r��^�j[�]��5���<+{-�A�o�gp��1Ѻ\�b�)�/^�"L%�ڢ|���m�KT�J#�)䯀&o��h�}�ĭ�*\�:;;�ؠVx���ϴm����C]A�Q4z��{ՖRo�D����*�?��m�tH�p �������!��F��_����ō_��Q�5  ��ŵ$[b�^�IWe{0s�O���nwUC�")� ��{ל59Xzj6b��Q_�A����9�����^GR�/���Mg3&�vdVe�/��>t���(n'�z7W�铆������L6��n�>�^���^kX���L�>R+�������6[��:88�:�KG���B�G��e���?d�NA�<���W��9Qm��V�/+��;\za�8D�d�7(��l.$3�+sJP u��cV�:��hO {�$Ƣ�E�fa�P�o-	x��g&�a-��3�,i�9�Z'&�xT�ߪ�%&6(oٱ\�;1��k'��m-_�����X����`�ܛ�Z���۟S�d�B� ��ҤM��A8����bM���8�BH�J[olum�и���ݖ�;qj�5��+�2����(�w�<rm��L�Ԁڗ�^-1�J�� .[\~�/����Y�P�t3wܪ�)���h&��h�eN.�׭;�vލ�^X�C��[��%�w�v�}�"�d���YI�B�G�]E&15�̎�(N]|;ս��,�c�Ww��3vʦS�rΏ����^���0ϫK����G5�7"e���o��������P�p1|�f�/�Q2*v,��\�����ι=
�F����SzZ3ܱL7$��d�C�Y�H�����)⩓d��CDZ�A��D<ك�e�'׼�0���J�?�*�"�;���Ǫ
Rڂ)k� �,Ny�D䓭����m_�z�݄l5�m�Y�fx�D>a��[&��a�2����V�(8��,��/)��H��;�{�Aq��:pj~M�Y ����}!���GЕ����5�]n{_9v�4��������%��s�V�mR�&M�
P��޴K\H����0p���pS��';��d縗���G]X�g�eQ����k ��8�y�����z�M$L
�m���6��R�^��R�6ԙ
*�E���0�T���Ƽ�夀�*���O���a��$���=s�����.+K�Ilx�VS�xͬ���Ծ��7�eTP� n��T��+lN��U��m�fc��G ��j����o�kY�ot�س�ꀱ���T�^I��U���n��Cг���k��
8���W`|�Iwm�.X�/�{�������*�~��%�U���ֶ�&����s�u{g��*��n��6��
��Z-l	��͇�sՐ���Mt�� 
s�� O��gPy_$Z#�lq:�z�������ɋ��h|��X$5�\��W-��O^�NSUV{���Ǡ�4-%�"��8B:�R����e������B�3٠ҏQ�������`5���Ᏸ	��0�2��=:�����[��E�km��l�g��y���E�Ed�窀��-'� �"��3����Z�s��]-���}�(Uh��oH��!K�DF�����J,�=�z1��[O�bb�XМ%�`g�&�Vt�O� ��}�f�P�DQ�ל>�lif�����1��N)�T�78Z�]�K��i��[U�=B�As���e�q�OR��#W1���km8v�:�Nq.�Z�k3;y,�Uzt��Z�
���E|M��EO��~����g~�M��x=���!���8u�/����{ɴ�+��Ǳ� ��%x&�W�j�M�'��9'������H����\l'�����]�m3���"��h-�P�����:�l�k�u���0�羓6�Y��3\��O���/j*�A���Rv�&���kP�<���	�xD.�GO�=r�&#�cRnl�N�&�k���,������h�W2l����ۇ3%���&�6��Oo����%�q��^vs��������lv��v��������q�o�C>�=��5.�i��~@gĥ��������q/2>U�9a���K�*��t�ﷲ:��H�Q'ɜ��磌V�ztՀ���m����i��N�;�@�+��ǞE �e���	8�;�ܺ)�ߓF�0�'�~����?�6�Q8����/v:%�^9]�9�d��Ù�� *T]k9�ω>���Kmm��rd�NZq�$��pI���bA��m��8�1!!U��\�!��:��,C΂���_f���+��)ܔ�.b�5��#��d -��K��-��I��g��Te+m���s�;�'�	ʎ�3ld
5L�ڶ(Ýک6y���x��l�K�w��T��C�������pU������j���o�P���N&�Ж6É�<����]�Ѐz��tX��p�h+�CȨ����* ���q2�M�HmO_���Y/�l�:��֋�W�e��ٝ�
9�릓D�OگL'y���w�:�A��A�٤�B!w��"e�C��i�7�n�g�X"��'�]��=,���b���/Uw�f/D2}j�Cp�m�xS���0�gx��<bu��x��W6~h�Cx���j�//�B5��0:���cPsՈ=��� T��
Ĺy���G ;|6C��W�*�2��VU�&��f�u�1@sf�
_Ûৠ�u�U��\ڭEɁ}�
'�~* ��9�5�=A3�:��z��rKX�bi�i�ʛ��$���[�(�m	���1m�a͢Go�6��k��+�I�5ذ_�)�I�������e.�;7��Uv��JL�M��a_���Q���'�G�V8���֜�҄��'��N���v?7B�1���{'�2l<1U�@ja辽�;-;I!��[k�f�f���S��hLѸZaa&�
�'�-�M�p+H4�bh��T�.$,����b	"�d�D�5G ��Z���f��J@Z����bQ@2E���;�E�����>q�ɇ���x���p��b��k�
T�l�J"������z�����
��֚���������S������6T��{6��>1���I��vF�M�CK٠^>�C�+|5�m��Xs]��.nC����_Ƕ����
/��	>��Ƥ8���H��=�5�Jr�g�ߢ��XD|�:���sǯל{���K�}/�(�,&7j�s��8��.����� ˚H�-u�'�G�B���bQ�	T!�Ě�vRC!�����\IE�e6�f�]�v��v�]	�7��A\��yno-�\e)�zK�rG_�C��<��^��Ar�{w����f̛���QЗ,ޣS���[ʁ}ҕ߲��ϧ�B��2����-�L�~��}�^���|�I��5*�����G��Zv�|N|�zЊ���Ms��k��命��g�S�8��"Xa�)�u��m$�q��#�}��g�0,�-�.{;/��I�x�!tF|A���OQ�lj�Ԉ0*��?�U����$��q��e:���V�YãT2�`Q��2;at�ŗ�.�Ws���^_/x�\���l��H�\��8r�$b��OT_\��`�N��1�H�p��\Ci�3��l�sǲW����~����w�l�(n���p�_A�?7d��JQm|�le�!x�^pw�P�޻��/�YY@0�rq0�4.��(�FĔ�ϕ�l�Ɉ;��PiS�������o�{�t���'NНP� ��%�jx����{�ݚe�U���Ξ�O���ss
�$퐻�D�U+�'�H���D��=%Hy)��=���fhh�����^}��}�����)c>=�q�+X�2'����B�ڈ$�M�CM�'c�/���-����&_�Ķ]8բ�QxK��dt�?�u	�]k"Z���97p�����Δ"�n�r��?oQE4�mb�x����Z"���D�0�.�lc��ZPמ*�w�Z�����:��aB�E\�g<�#�[��-}�'��2��5\k��Y��Hyx�Ri�<��S#V��h�9+s��(�?�4,��j�F��}K�y��]�����yWtҍ����˖-{��6��JP� �'�My��e�&t+4��G�{�L�q�ߓGV��IKOdcEk/�~ƀ-�fF�*D*�6~�Z: ��:~E��^�������o����0������і����38�DI=�0�Y� �j����YċJ�Z*�=��i��hӝ���?c-�7\�R���U��_���
�<��M6�#q��ʞ4ϔQ��O?x5�P�8Y�3%6�8�N� H��
�*�[A)aԒm1gY�ʁ�Up��-R�y��@W�6'�`c2~M�H#�*2JT�#-�CC�8��	-g����ŊB����wX:h�ཪ@Q�[�Ĥ�|����tj;C�������M��=ך~��Qb�Y������=�<l��=��T��9?z⧦9n\S��q)��Ҧ;Z�jq�+Q83]��;��h��a>t�{9�:jކc/Ԁ�F=�A�l
jt`�)�|:�Lg�Զ��
�`<�󀛊t����W�X�s/��)^ɌH�T-�\���SͯaE89o.�M��|H"���:Ɍ1zw��d @NOϬ���zq@��Y�:W_��;��H�Q>���.����|����4����`y�jl-OH��J�,�"�Q��ޟ1��Q����~��^4�q�~]J#�Ï�*K��1��y7R'/T2�3��l�G�$ΐYc�F^�%Di�7�2 ^i�؊+�{��Y�yh]��!H�/h,�t-�YK	}i�ҳ+��N�o2@;��cNu3Y����;���/�}yak D��v�I%d�~Za�?1��j�4����54�@��0�Qxk�M0�R�S�,|u���0����N���͆M�>�����;!Ub&a}R��R��V�vb،iΪ/'@GE�5$�b�2��͑�������=*l{:�ؒ���Hl�*_�_HW��d�}Q��*����KQ��Қ�������PK��aR:aַ}��T�R)����D�{^G:�IQ)^�ª4 �+��a�Fx6Yԡu٩dP�L��m�'�;~���_����LYe[, V��Y�qn"7��s��~@�~�V�����\0N_�v���ߧ+�
Sor�uK�	�މ�W�}byG��A�b��8������jy�Ra4�\e( )�U	X�� |1�?@�{=m�X���TЃ��V�NPyv���dFT��q�|�M��RV�H��>��Ⱥ5E�D�� |%1}�^�w�%S��m���lM�a��D�_a��&6�����Si��)�q	|�l��}���(��毯{��
F��s|��x�N��7���n��еa�vh����.���,�'x8� �S�**g�t-C2hnhF������b��L!����7�D��EH�KU��u&ݮ� ���ZE�0)v�{Җgɻdb؍��ֲ�N5�
}{���yWt�q�7܉D��1��[��h����t�¶����e��mv8�*���E)x(p�`K]w�J�J����)�ǫO�;� �_�*δ��$�����/cP&��jl'�z��pw������Qn�-R"hm� �}Z����Rm�:&)v��.�5N����/���w9���Q��ܚ_�3���I��OY�~�Ν1f?�ph�5�G����' ����v�2�m�s ���|��� ��S��~���C��7B&��)��cQj��8�Zӌ60�2���+\�`7'�N����b��Ԍ�s��c��~��|�j��{Ҳ_sq����Kʪ��1�,L��&��R���R��uUa�ʍw�R��X������6U�@(�'')��9�<�3G��DW�=��2}���!k�QJ8������|�f��7��u9O�wq_3 ��⎡v��/�� +��HR�qxXj�3�dw��
V��N[�\��l�XVN�&XN�H��ծ� w�Qv���E���/N*ʇaV�4-e���n�TP���6:^����E^2�6���b�甙'E���V�Fh]�&�-'�������^�q3o��S��ZC�K}�y� F�Kt5 �Z+횺�Κr��H�-FCU�alW�I���a�?oL&����'Ip���b�cگ#N](��r��e�f}ݻ�#��"�K����؋P��9�Y
ї��9�L�)�=o��Z<j���d�����$��R%C�����tF�ɀ���L�(�f	R���
$!sh��Y��ǫeS����(g��`b��#�]�(B��e
<�_F}���E�7����������.gѨ���R
�f�K��g^�} R��d�ԅ�Q'u�ǎ��ɳg�.��-�<޷n�_r�`c�
/b|�})��-���{�*���`�������h�pΎu���O["T���9�E����+9����Ĺ,C8W�0[�B���e�����s
T&Kk*	��O����3z�l��l��=O�n���U��������o@ye�[j�O�U$��W!��I�/y+�Qy��֝8���ي���6#��,��D�Tғ9~�rXV��ur/�]�zEb�%� 	a�6�2��ֈ� �O��q��T��)�j�2���a�pˏ�-���v�-2��xYp�TG3��ܫxL��_�"a���*�!���pH:)�l� n��'{'���?���������Rj���)v�m��IQ2Ϸ{�V'�$r��>��H�V�3�}x����, ���0RE��z�8S�}�C�� ��d������1��r>���0>ť�d��9��]a��-{�����#_�0�5c�7���tE~.�'W�DI��A�A�7\ �v�:,7���)#'�!�$��v!�s'��3U�«Rzw�uez���K��y�z1�1Pb �\��hI��T!�M��a��� x��H�HwA�	a�s��7����lI�R��S��2�g|:�e���Q�]"��YS���7����Ly9���Q����;�y��a�u�h/�1H8^��	l�������J,�8��jʾ�z�m�=��ܝ>,�k8�۲���t�ǉ��̩����X�fz/U��R��:�8O3[<2�z�������[-����A	P
da�A��Ό{"�à�[<`��Xs���(��Jyk�~�)���T�(��VC�pD�:������(�c��/0����I<�]w��ͬ�t��7�q��o���������Oc[�)������ت�؆j�Ȁ�`6���bp�8$��{y��)�+ eP��7�:����p���_qd�Q��G������ .�Q��~�3<D^�!y��+@PD�t)���cN���� ϱU��8k�!����}X�j�qY4�;vy�q�ZhV~\*J�l&��7j��C	;�>�z1�˓b	���Ӆ5R�ȝʷ!ǋ��Y |���HtI:J:)��%=.+.��]�f�plj�4�9�#�/#̫��a/����]Ɵ=8n#8Tﶎ���1��M�ls$�$y�"ɜV�=�3<���㾨Š�e��x*2�K��zKZ�<�TXf�Lsg�o��4�+�^�Ԙ��O��(�XoT��w��s8c<]8Ծ�Rk��40]�'#�n/��m�Pi�E�Ry�]�����]F˘c�{
U���'�&C<���	�����S��q^&��C����#���LA<�0rYo�)��܂g��[�O~a��&�g�a6<�EpK��k�"m[�!	[n�9�L���:C[���8� Ԥ�^:J��żR|��E�^P���H����������26w�$ᗴv� �pׂJ��1;IN���\SY�=N*nX��s�۴�W	���D� ��M'Vd֬%�28'O�=)=���K޾�@���"��C��dp߅Wp~�����⯇'t_n�K0��z.�B����Y.�Ϲ(�Qr�1��-�u[b�H|��J�l��c��L-�b6��Y�OߵD 1`'_���+ԛ��v'r邆�{�tqQ<�.Quύ��d�iNE���ƫ��߶ui�Ҝ�Β�j�"i2$�v�--��ӯ�K��[zz� [�l��G��Ɲ�G����ÿ�v�R��b+�T����Bn����r��ݲE��8Ï!UH�]�B}f������|�F#Φ������Fo���i5�����PHp��㲹G��u��h9�c  =1פ�������1_������1��X��2i���S5\�UIm�{Q�7��]�vD�������NRr7$������l��B2�.=k6h��R�,��'�����gh�ww5�
J� M&�5�z7��$t>ϩ���J�6�	nT��$d��ù!�<��\��Q-�Yv�H��{��Ýn� ���� &.+��5ti/c3�8��q-�D�e�Y7~_�eRq%e ��8�߭�ԙP�"X/���.Z��a�
�X����Jx�ڂ��d2m]QU�W�R�ʢoh��=`P����h ���ŭ�g�F;�8l֟K�q}=k��*A�R�u��z\�L�*]��B�r>Mv�p��]/d�o*ኹ%W� 4ƨ�!��+~�eN�y�:e�'��d�2�&�I
r�(4Uڈ�|iB6�P���?�Zw�9���r�����mq%0PH��U���<�^Y��/Qz���,�l{I5�
�M�Њ �1n��rwVk��k'pm��`"&�ߐ48��G��;&K�N�^9C�"gxt�_����z���(˚,���┽�B��KH�"<-3������>��/ ��e�x��M@<��#(9C�̮�j�$�R�p�G���B�/X{t���m��ׄ`W��Gc�=�s�jY*�N��5Y2oV+�?�,��.�il�$��>g��*:��h���#x�F�'��B�R��p�qm��AMQ��"ԙ�Rz�ܷ�����#��9 ��ajl����?=5P�x����u�RD�6�e��N`���Q��WS !,r�x�~�����5��R��"ꭁ�[�eQ�n#W�Z�V�	=�j,�Q4��YǇ�{� �-Cֈ:����3}���I�n�L�7��YG�a�_WNțe����_5� 18|*�船%�z��z렞��ٴ'��N{Ɓ���2�~����Ѭ���.���L��b�bPO��s����X�,F�&لSb��]h�:��9���v:jC�t=�%�Z.}�R�D���d4�����c���jIt`��D�7���g-�ۤ�u��������!g��GN�gM��G�����|;z��l3�����|�<S��> �O��MC���0@����6���5T}4��	�`Air���(�Ug^7��i�eۢ��xo��������1-�i����w�D�r�mF5{��P&�L�����5���!�%�m/P���l2�9�6�Y�/Ⲁ��0~gb|Ј�#�8#Ǫ<{S�Q^MLp:��\Mo��-
$m~-T�d�;KY���atŉ�|�0;��20lr�����>c+�Ks�85��d�I3���x���!�R��[�:J��m��H!�O��Z���x1sE�Z�S��8��]�����iq,g���J*���z ����ڭT����K|�hЌ�W����������;��Z�o㰐 )q��G����J9�����H� �t�\��e�pdΓ� X3v<�����j4A�+��F�磪�Pd���q��@7��}�5X�1b����qDn���Cڀ���1nw���W���`�36���'�,����u]���)@�h.��KRƬ��i�!�=���fj�-���<@����_y ��<b�9��Q�˙SN��;��1g 
�@@Z���a��=ݜ���"l.�D��k7`�;�. +�w��4���BT����&�ؤ�U8N<^]ξP��@����rm>E�\���~W�lu�TU��A�C߈N�ٚb��#�%�*e���4�b�1����8ص��!k6۹���m��u�H�����2~c��:a�kž�~\��@������l� �ۙm �����tTPk>��ev�;�_�o0��V���N~�@�8z�)b�Γ�S/��2|��J�&�mNP�ô�3і�K:�ro��A�`�߳��>�e�j�LIմ���6����������h1��JD�T�Xv�Q^�w�s�p�U������� �W&O�1+�.��.�����r��x
�GH/��/����|M�G�'-㝇,���r�J=��$�p�n�e18���;���F�A�{���̼� ^�f��X�f�5`�4����	�k'�
��MZ~��`�_�^wE�q?� ��I�����E��<W�����������g��9[��)(�"
j)�k�������|A�1�7��������Z 
¿[N����m�S�X��;��K$��,����
�x�$h��/Ѱ�0N�����{B=R{M�7w�d��X�V���$�U��-a/�e�52<�Ƹ�]`��E��T�.�����x]�wn����%����I%y���� �,�똡���/�|�*�V~��&h���m��r�^?�.��~��ZZ|z�q��dE�a��VM.�;�y6������R�9���{�[f���
��RƹY��N��N-�,\<����́���>�����S��}��cR��."��H�������w.!0�U
�B/r�I��Pt��>�S@��|�\H��#�$kz3��+ټ����cƱ]a��;��rQ*��R��$Z��	�j�Ja-���n���c�����Z���T(z�C
��G��(�9��s���]o+��SꞟPz+��,���q��Tb�%:�q�C�aϜ�h_��%:g+��ֻ�.!'?��.���±���v��:Z�Nlw�>Q�>茋�X0�r�� U�T�Ŕَ�<҆��[6fe}w�Ua� �I�{b�छI��L=� ��?_�[�,NO�(�x��9<�H���:���8V�8x��"��o��!��p�ap=��b�XIy{�m��qq�����a�(��u����n��=%v [Tȫi���>&)�'�T�(�S��?��!�z�Nii����*m���NM�����C6�w�V(3����?( �dwYE�2������o{s�h���1	ц;k�
�H��Ͷ�6�S�%��a[��=�� �����te^��v�D�]��2��8Ә	��E���y10gд�D
�B�t!��A�(�+Z21O�MNw��uʸ��-)���ѿr�y ����(4kbZJ�>B����O��ƣ�]�a����x#�G\��{7����K�����d��b�D��=͵[(n")Z=>�ߑ�g!_rB�ȷ�wSmd�r��TK��E'ZF������j3!�Ƽh[����3cN����M1����tp�%�Qb�DS�$��L�F#>�b���?�����x���:BZ�*0�3�LV�ğH��8��� Ն�� �_���V3�����A	L�����6F%��6D���*�]+^�{cvK�<�g�a���{h��el"�lb�����2�u����R�ը!��Y
�J�3̂�G�?�F\����;�n�-�Muk=���֭j�^��sh�nj��P�-빘8acٳ!�#�Z���PR���\�$Z�,A�fl3Y�0��*���\�N����$b'&8rU���F�[4S^��f.����.�w����I%��^�A~Ҕ[Z�v��s|�Բ����J��Xm�����Z�t�*ne��H�X�r.�����(�R%IfT�,L�M���
���m��:�&��Sx��e ��Fr�Ohͷ�E"�r�G<#�U��S��f9섘W��N��:[�w�b���&�7��
?X�甊�%|B�gV�<x0�]��|юK�׫����H��7�pD��m<�,�ǖ|�o27�.{.R>�X_SSQ���^-�
@�)-���>-�r�P!�I�"2v(�1��t����W�T2�^1�J���=��M�dՃ=	���Y~��*���HX��29��Ң���a�CG���KD��ccN0+� �પ���Lv��&5R��/�Ou�چ� 
���HS��ތ�`',/�$�2o� �z-��9P�V'�2r�����1^����3ܸX�L��q���Zǐ �֯1&34s�A�Ct��4uє�(��eZB
+�J�Ըw�"�7�.�O����=�}SW�:���r����ٍ�	{��5�'��_�u� nӮx�T2],PlN䝲���ܻEl��\�-!*�
zoO�`{ʶ,�ycn��M3=%�n�" 4��s�X ��!����A��JX�)�.�$KN��l��p��9���}8�������gtH��~�'�V����R2L&ʌ��T��������ȽC��x2xmІ��b:�_�Ӹ�y5	�������@'�ϊ���PD�(��2����'SIg2���]���?���u�H_z��x���OVɇ�l�O�Gn-�(�*��Q#Uh��N�Jb����̧,��n�~��i����=4~F�n}�:*�[�o��e:ſW�ӄ6������ީA�Z��vVuA�ϐj^7�m�������;�6��b$����Wھ 4�B~ĸ�1��&-�W[��"�TL�
.�߸:Z^>�j:y��UM~н,8 �eH��6 yX"�&[c�V`��B�ʟ�Q�'���D��L���)0�*�j_=o�8ZZ�l��(l��}i?0Dm�����jla�8�	�8�c����bN��g�)c� xōC�Qx����2�\�(>J����/c12a[��RR�s�+*🱻��_I�sӴ�eI��H�SkL�[	9+Xui��Ă�eh6'��תo�L�F�C5f��5���Vd��I��H���b�VF�U�y�O���a��|� ��x�SP
�4	:_�8�����"t̭�xò���yf�M� �g���<��Q�����֚&W���U��,�}%�̈́��Xp�PPb�}U�zs��o��o�ji�>��)�ǧ�p(�x#�N.�~Q�\KS�JY;�S]D�|skr��9l��A*ʘ�-$7�����\/��!�P#�ǳ~c��;'��\x�OeZ\p��<�b�"}Ҷ؞zh�x�۷�����[��r(
2�r���mڜ8_b���`�y(���H\ƌW��Z�̬o���v�ս�Y�NY���tN�@����*�b�:	�5�zl>3U.l@��M�HW�XT��k~M?���'+P��܎M`��w��@g�[�뗾�sIq�k�7C3���N>�bw媦<�H)��q�L� �TDt����]:͝�R���&S+�$�
,�yax�S}U=����6c��{�kȀ��t�����o)�Y.ߋ"��S/4n@k��u���(�n�*A^e��3���e���X�u0�|�MSe�}���##i��d���QIo���m2�u>�8��O?n��a�X�r�䙦Y�h���~��������Hu�L�<L�yz��vqS���A4**5=�)ȹ�}|q��q|�������_=�}Gr����{}�a
������M�����6�� �%V�+�f}�S�	��.L����b�A�����4@�8�m\,�l��D�Օ[�+{L���!��)�7�2�E�\����r��t�:��)v�a<!�� g���x�i-q@ء�B�J��W�8"�d�C����F��i*ȷ��d\2��٥r�g>�)���ZY����J��yY�џ���� �����ޘ��Lb�Jy���Ot}1��E�Oq�k�֏�T�H(�×&���nՒ5�<�H����7[�iW���ŵh@;�.Q����)?W��.�?_L�I���~dSQU�1����p6*,�b�2jn_ĥ���҇8��		�-QKئ��hB�N������r��>w������@G+"O"���%!�)�h�K�n���h�ơ����~~�^4z���z��4����ڗ�^v{�:�KĬ�JYqFH��� /����6-	_�OP��2�������|�;�y��)d�ؖ�&|Ur�5>=������r��8D[w^V��?����֐��_,�G�$;�BT(E�2��1���'}Z4����%��x�#�73���_bs�`uQq���EV�#�ӎkTO8! ƙW'�����_,����C���y�Y���	��t���!G�q�+�a羋�k��:@�����XwM�;㕂��t���(LG;��#@U,P_EA�x޷��,O���ֲ8a�2�I�^�_�̴�ws��Z�`jaμ" ѱPR#phm��@�{�ҮS����@(�0/�o�{�fO�`��,����|޴����ui&�B���	���3�Ӭ���<��$ANs���	�a�b��n=f;���h��~�����C��odvM���q����|��Et6X1Tڼ�����n�tϯ`j�����֬L+K���!��������� �^Ot&}t�p�6�ŸNO4(�mk��=�ך�{�=��%c�Ҿ�o�#���F��$�i��9E^�3w�[��ݡA}uK��������zS��2Z�Ad����x7�*XN0K�%6�\q��1;��{�7
�B�{���I-Oc���b��|J��q�/���\>|����M�6�RD&u�	�+0@w���b��җ�v���>|�=�C}�F�?�vL��3E�-8�}c�N"Í��p޳L�C�2����F-�͹�^�z#.�c�)��1��(���{y���O�v��V��3(�G��\0K`����mVw��r�Թ�zMd�~��F���f=F�Zݴ��p��45ic*do/,��/�m����9[���������5��L$���:0D�cl�1����*����q�}SL�m����'@�W��2��H0ٺ�K=ªz���1�."���vխ��|B��-���Y�����+,DB%��V���a�GA2uׯ�}���Þ�-;��{���,/��a��	�9s�G��A��3�g�K��Y#��ň����}�\�hׅ��(�v͘4f�7v[��L��hei�W�u���xFʪ�f:�1$P���E�����;g.�����G����'�����1��Ă�	n��T�*����"֒�W��.��ӟy��6������տ�g��t <'���:{y�<�5c��@�.���/�2�m,�?�3�V`�y�T�B_\Ꮽ�֋�7=��1��o[�.�6x�DI�����>�ÔD+�21ϐ`��B�� ,ꮔ�`E�+�W�[���A@R�&��_V�Qx�0���	�(\;�	�:t�圗�()���h�p*~7�
�!�e��T��K���sL����O�m̏�~1<m1�hU(~�ɢ���c�	��}ۤ]{���	^$��Wh�Ӄ�β*$�乄"���͝9pƇ�ql=�5n���^�i�{≦:�A���V����<���5�'��ȗq��Ca�R��Id�-������t,������JH^R\s���Խ��Y���~,��V���=�$RvF�'-�����>���XZ�X8�E����T2D���]�����ū���ⷁ�ߌ c�i�I�@�=�������_���u �C�0�36Y�&�l�#)�.�}&�\}�O��K���"8�x�����g�[�nNf�S0�sU�8J�`�<l��Cťښ�H�����d�d�|d��t$���|�
t3�_5�l��z�j&��	A�e�!i2��a�@ ۲���>�B*��ƻ�m�T;" �g�����&#�C/$5���$j�PFf:ICjG휭l�h���� u�z�����Z� �(5��R㕘�˕��dNvP���F���2*�S'��|��3��>����m����`����Qf�E��+:�4�é�/_@�^n�ڳ��':_8��p�]D�N%�:�٦^�r�ϊ�]z����;ړ�9a�4�rt���
��L|l��������<ř�)�
<�4vz����G���a-��6#���K(�\�~�ձ�{:aY����;&���nH,9y�?0˻�pf���>X��p���y0T�A���h��J�*�⥝K�����V<j��y��̢�9m�	=S]#l�U�O�w##dL<)�S�;�bb�\��t�S��^�SM��S�t�J�=�$�R�C:9��޹,`�ؘJ$bi� �Z��u	t��\�Rʑ �am�Ҡ�kW��W�A<���Y�������D����� �J�`��|�ф�������~Z��8�QZ�zV�B%��if�e>��C�hx2q�<y�����M.�����l��e��%��B��-���riғ������?�N6 it��@�ň��F4o»L�}N.�����Xa�����0"!���E驶�7e����L����M�T��+�qb3�V�6�Ͽ�����°��T}�U(���A��0^ ���XXA�±�@���}�|�ĭj�1V&0$u1w�P_�$��(k���v�ѣ�b$�}����lȪ��y�,�O`�w���¼f�t�_�ac���Z���Ԅ��#����L��S��1zw�?�U�	�c���g�R�7'��래Cg�h;۵��|�{���!��[��ѳ\�郌���3O���Ԟ	�<��e��F����߹���	�7��Q�F�>R��9�	�O4���Gi"�wai�/��=L���/�a/���[�ζ�<W�0!�٦FM����h�
3�0ƌ�VMǡ3��<t�آ�8��$�3J��r��AV��~�K��f��`�����:3��_S�C�v{W�g�W@,�,<�Ȼ�>{͚��Ӑ��<��BRKt F�['U��9WS��FPm6KXe~뀍:�)������b���tُ�3y����>9C�Q�$;�з��R���wf�*�/�Ģz�`����-Mp4���V*�"���P>K9ab�������]��nPF�1�繅@IK��-$�����t�\�K��&�%���a��s��GBe?��ʝ	���UݾR�v��P���3wH}�ճ�ޠ�6���(����!� @{��t6���v��=�<�H��BY�
M�%κ��cd��M�F��2���v4>h���+Ǚ[���_*D��,��ع@k=%V-�l^w���Δ�o�xGW�Z&D�������dSy�rd:qJ(^�|�x�Z����L{�-B�I�3���˓<n*p�z��V9&������ O����*~������J�An��L�$n����pZ��}���˚��G�b9�H`�F�u��+�]��(*�GXZ4�&�)n�+��|�yځ��b�Ø��5F�������M���k�`M���^3h�lG8$�H���%\�0济���rN@AE�S�("�l|����S�E�8��V���Q,�'��{_����yKRgq�t0z_9.���=�M�D�J���Q��йK��=��/����W�-F�P���װ�N�H������ܔ��)D���h\haآ�X	Kw�=�گۚmt1�w"W��,vЉ��)P��-mk�h���#�ve���Mu���<�X�J`��a���;]@�}4�����E��OL����z�{z��T�T\y:9p�	`��Y���O��+?���i���L̒ҕ2o�"�ڷvJ��;��'�^�@�!cm�<&�r ��3
Qߩ�Zӣ�Ы!�
R�8����B��ɪ��$g�-���<�T}25-@*�`��t$Y0����d�p���TaDo��,���I�՘�YĈb�#{��~���Jv����&��I:�Y��@F8ݔu5r���lypЪ�t/#��J*�GL*��5_�+��vؘ��6�u�1LHn��f���=���4�^�M�����Rq���v]3�/��eѶaß��T9�T�es&k�FR�@��9�su]�j��B��CK���VWW
ή�X¾z8o�3�2u#���tr�S/��h�ħ����d'U#��Z�W"�"a����/?)���D	o'��Zέ��Ձ���x�s�5�^���۷: ��*�OX������E)��&�C����� _��`�X��P�u��b3|��r��85�m�n��;�Bs�m�`7�����/B����\��䬱@�f5�guVN��dbk���mU���#h��}�� C���L`��s�����K��*�I''��P������\u�R܇?d[3�"Yx�<_>x�7�9��:0�B��2���f"�{�����p��E ڦ�h�������K��b���T���S7s6�����A�t��_�r"�h��.3�bBn���B��s+�]q`[�RI��\&̸�W�Vp�Mz>w<	�i�vʨ���i{��Ͳ��~�ų<���Ue_W@БKh��S$Yi�r߳�Ԑ���/*m���.�G�{;�u`�����A�%���A��)>A�v5�X�����n�M]و�=�s�Acu����]�����ږ^^�^�r�!rxE0�c�y|��Σ!���J�Y\~��x��S*ֵ��7$
jPH��$��^q��g�F��N1qEM8[c��x���������&%1)�e� @���M�Y��;Q����6������02�<�歄بRr�9;���'Z�v��
�%w��V]�P�9^��"[�SA���Ѝ�K
a��,2abr�y%@(�v��Y'?10�6U.K++�S->��E��	4�~ig��RQ����]ȉ���k�Ϻh򬸾'ɭ�u<�a���ܯ�գ�Qq�V���Z�!r1��i��6}�����X�jDTF�����
|""��)J�(���9ܰ鶩��t��o(HΆ�Lq|��!��嬱��7-'���m6�x@8�'5�x����*7$Ԟ�u5y��䠽e?��˜v�#�ھn;��zH�c���`J�B��%�J�pe�\:{6��<n�:2���ұ����H��~�Y [4;9n��P��2����&��I��I��A6���8r�=��dѵ�~�	-,��#�W����^CT#��ؠ'���p`��x��@���×"���k:#1�?�Y�Da�-�g5a����P�b�Ǉ�f����)�y	���ô#�
D��*(Ϸ��B�$淬�JD����E5dv�nѾ2�㥁ҳіP��DLB7!��v?�J��n�������7d�x7[�Ữ(ڸ����G�<K�;�<ZM�[�R�����\�d��`��:�t~�a?v��R����ef�6D��IW�y�_%�d5e3�]��L[b�����(�B��t[ƣ.��<2Xޔp�ǃ�)o�i��(*��_�
����Fӎ��;͌A� �4��5�6�>+�$*j��r7W�o;4<���sg^O���F8͵u��q���'\��(���\���h�y�B�a@c�V\�����"�-���Jz�k�F�����R�go?i����t�CO`��;�����"� ad˭,�}?��VS�����C6>�|�i<2��Cn�\\iL����)�Wt���y���c�מ��A(j�3;/��Qd�6���ϫ�U�̲�4��� �srLt�����S��k��G�It]�?P�Ƈ1�)Yh9�B�3�������N��~N��l _�Ob�H�����e���D�t͂�`�Y�ߪ��k�aϑ�]�;XZ�cs6��O���<�R8 \�8sV�#,�$չ�5�Xl�}������DY4r,��Y��;E�hL��]�|�hȑ��F���<��62�{S�+��J�z�Vψ=V�\�� .H�e���A6�Lo��3�U��+7e��_6�����x$��מ2��9�S���d��ay���R�$�j=��|���;�(;�L�J�s55T��=�Z�eƩ5ѠVW1���]~����+�ߏ�%���6Sgt�\���jS�;/g�ć:�T?���|Y9+�Lv'c �J+��>��}C�~�ڵ҂v���0�4|������(%�|��K���E�.=�T�4 u�3���[yaO)�vet�����$L�M�ة'뜰�܁��N=�Z��ݻ#}WQV���Y���
gux�-��`ңJJ.�B�H�mmS{���s�&���UXUCy�[��i������V����ߗE���@� Pt�$CTbb|X��8�� �;8J���tdM�D�L�n}6FQ�zd$�rnN��H!�7����� �{l���F)*�>�Jp%�ӰcT�����)�ζ@���ƨ#�c6�Ӈk�:zaz�?lZƬ�#�s
;0i#*�;OC�"��X��(,��#��r�o%��]���B	 %������s���X�pQC��w��bq�_AEM��A��᭹Jƚ)	@��HYB�5���*<'�6�r��}����|����1�L̬s!��i�]�)�t'�0>AX��_G�#�a9>9F#j�/�,C��]�pډ?��Z��g�aLh���W��]jٽ_�P�E�RԿ8�[O7}�rh8�1VeV�J��aq�+}��ƏmŜy�kB�S�ebM����7��p��q�]��<��4�l$��b�J�����$௅�A�%��c�`���̮�B�P^�&��i!	�G'}n�	ޮ�&�Zd1H[M�#D=�csG�,���Udu���[Q�V���������ޘ��7tu��]�B1D��j��$��V.nJ�� �]��2��KVca�[=����/�SXJ��A��qA�H�-�zC�k��fG�&�����s��R�l�r&���_�E���ۯr����F���9I� ?p�������!��8��g},�T#3��w��;�9����Ǣ�Hs��d�>��j�-׮U���\E8p��I^i٧]��Hں��@Vy��ƂO���1�]�/:F������*�B ���.$	uC����Њ��� 龞'a�7L����6���a�.[�ou�Q�f6*?9#n�27	=�Љ�r׻�3O��*�O�o��ѳ�)���^�K�!�Vw��\�T��o�����j@��-?6��*�Ǿ��:j�
����W��Ñ�2� `�3<��T? �?���Һ�!s�Ru ���d)�s�kE�Bܤ�ڞ0��z<��<�^��&W[ضb��.�� �\ӿ�XËT��fn��
��xnsjYz!�B<�yu����TЕz��s�p�i�iK,|{^�����V����Zm �FO��<Bx��яq�.� ���r���cQq&A�@�*y��Z�)l"H�"�7�$��%���H�&��m/dD �H��;zz�!\������"&�����(@nP�
v��n����^������ E2M�ƿ`��c�yOkN6�a��l�l�����tx�G��"FYh��!�	s�Co�qQ�&���F</�rI�M�F��+͞��_���y��`񔸹eQ+��c%���Dnb�vB{ H���v�4ƪ_�9%�)��G?s�ŏX�4X+z�<�ێ�ϰ��詞����˷�$s���3�����=��4d���8»��x8��=��-���5�������J��E3�*D�� [j���xݶW����N�����ecX��x 4K�� &������%�<m�Qt��'��X�oU���XYG!��j���#j�IqqN�oNe��`5ÒP	1����Ϭ�7MJ�g+��f=
i��98~�D �M��z&/��Xb�e��.��a���0�}��1W%���N�ٛ�>s��A���p�ͮ�ǵ�U��`�{H%�S���_ ���N�ɵ6([Қ�sp�>�ȪǘT2�`�k3K�>����w����V�cs���O�p�q;O0�g����W�;]9�s�s���.�0���J��?�K �@ԱIQ��*�몷�'��g꿖*+���?>KH�|�ڼx��/t�ZEM���{&�H; � M0�%l+�[YB��l��3�'!�+��R����H���*YN$T{
K�#"�>+ϟYMLUf�ŏF��Mv9�s��l���3,��k��0���-{B.�P5N��n�A�I�U���N={N]'�#ã�w7�3�ԍ�$)P����@�12ׄ�_�xy�
u,������2���6�$�݂e�6�B��a���
�"�0��'����uR���v�b�X��%[�����grj=}�7�kS�0���'�z��:u��t~�I3U����,�o�C*ʧpQm(��N�8z����S�eʀ����!e�~w7�6��t�>�D	�n���?c�0	�2�5��
��(��'X�ˠSM�6��·$�2Y'1�5h�Ǆ�RN����
x��d�Fۇ?_�6��|���zb�~B�)�B�~�G�S,%|���Q'��b��A'͙bF>Kt��B��6蒏���W��^ظP�u���ɉ[��a6��U��.7����噤�Y{_��c���(fv-�0���� i,��d�A��_�3Cˡ���W����=��-j.���Qd�,��r�V/�̷'.i]��T[)-nD� B��W&��N�fʚ�yi�4�<��������E�Jv�gB�0��$1�q^S5�R<ߪ�Vw����.�%��SV ���X\�yj�ifmƧ´�D�s�Ƙ���Q�c��j��ս�7+7`I�jt����Xk����\0;W�^ю���y"EW17�?�-~�W����L+����(�6��W��n�˯�cx��o��P�<�(�G�0��-�`��vT���a��8'.���sR[ay�E�[rE�K@�s��E=���;1p{�+�b�ϦO�/��ڑ�T�p�"Єb`|&�3�X\ڵXn�cx�������������Z1���{�e�S��`���\Q����t�f����%�~��t#��h�^��a�j8bCk��! p��@R)�k��f�{}�q�����*��Ϙ�3�k���+>���-4�HF4k@����x+�.�)-a�5$q7���**�t@�s�f�n���G9|��}��6��(����������.�+�dU��UhP���p�{���MA�^�)^ݶ���}��1�}���f�*���7V%����o4�I�I���<$4���4���r�-/�e��j΋���E<2��{�ڭ�� �>���=���ރj�����5��%9K��Z�ʹ���于|*�hoB�g1'�w|6��Ah��®x�:�d<A��\��A ���wG��WGK��:$uS�B�|n>���f����#��`{�%�HH�T��!��VVf]vA��[��.C�|��8a�C�:�����C���H`�ˌ�}2A���o|H�Ճz��P�I���d3�%H�����nھN���J���;+
�w%EE<�41E�3AM���x�A2P�ʑ������*6�ᔝ�(�j�6i��ϟ+0��A�!ʚ
�����;�k� �?#r��,,��F8��)	��5�\ŭY�ۄ�h�����U����!���: �!�x�������)��r��\	m!"�**�L�81 N��=��1���u�]Rj�$JRJj;��t�,R����7qe|fe��fb#��#1%;����8 G#e3�A�f����wY��u=���m)�� �(e���Q!�]�K���w���^�.f�L��`-��x��=_
*�*�}`���"9�fJ�cʒ�+~3�W5�H.�%�BC����Ef����~��\��|�rB��z-fiʵ���%)Zq��svdn�l����}f�@����q����^�!]�Z�Q�)���K��S�syA�w/�l��7��$�����R��z*��8���S�	�&T�5�F7��h�� ����` �3:G���Vx�J~oVN~AQE��?��uSo�WshI�B,��̶Q練�<�L>�pD���5~6��*&�A�h� g<�&Ze/�\ vEV�� ��̋{���9�c���(��|J��(⨢��h�Xuw�\���k[�b���C�
߂1��X�?s:�Uøg Ke��kF��=;iG�\:�:rH���Z�TϮ3a�E_nI�Z����v�E����Mx<(�g{�zn�t��GaR|؏y���bC�Çd��$]a<�Z�# &��[n�r�~2;���
W��z�`�ev�4IPt�8Ҫ|p4��N��hNx�$/7�������<�ZS�ws=�,$C+-�tޛPE҇=�DD�se�}qV�+c��O�|y`��UXE�B�	�yW��6�V&�!��r�ށl��R��m�6�O�Ry��&�7Md ={����y�����VD��������<)Y:����) Ν����6�*�k�6Z_����TUI�o85����oқ�q;�!5�2��!�ϐ�q(>Wau�ԛ���� �.f������A�bj�t�ij��'�`���>��z�D�Z���֐j�I��n�o#�ɟ�f�
>��@��2�B�l
d?�ڪ$�3K�Jd�Ԃz���vϐ���9��l�Y(RN5�+ƫ!�n�nD`5s*t�M; ��>��� ��vN�Z�, _/�y?\��FԏC�����]d;�\O?��=%���z���d[����]�����*\���x�y]'U��/T����Bkn��_5x����B>R���Jhq^#�DC�'������!�;�P_u��/5����
xل��h��JC��>��͖���ŨuK�t#+�!�6x����땽�߅�T���D<��e�c�F��h�9��ڏFe�����	nbrs���):1sC�݉�'"��X��tb Y-�z��;e�{D��l$Y�^���w�b�n66U�3�q�=�4nb;��z1=Oo�v7B��"
��&F[��v����㽙,#��.ASg`J�������2˶ �m3��E�X"��������k��j����D<"O�C9��]�u��8f���6趖�P��>)3��cE�;0�Z�e�g�m��� �֕A���HZ�Ұz�@ژ�XV	�/�����_`-6��M]��`�"�W\d:�������v�`�����)�O��Q����Z�T����cI�
���#�qcԾ�[~ ���`�`B�t��eZɭÆ2�l� s��f�*�xf�(I1C{7� �#K������{zK�~�}�O��NR��+HոU�mִ;;��.�ڊ^�b(Fִ���9F0�Y@�d\;���� lbc-)X_t�kg¸��������b('s${(��/��baʐ��2Rj��\��dʊ��8T'1�gf�
A_`����>���G�-Ȭ?+�e�.���ט���vo���ȽtL@y�^��<m�!n���UV��#�f��������1@��㺩U�gL��.ķhS�s_t���sK�:o���߫���-�U��4��K�����!��*���E NE�l��!�?�/ ��H��?�	L��]�<	��H8w�����tVc̫ �����H���q�
�cQ�
�������e���Ozh�ê)�
���h����DĽc���Y@�Dk�� ��)��H�[���J����C�}��&TY!᪗*������^�α�k��~�ByZ�������yI(>w|�L���n�$�bܶ�|�J���#�� | �q��|����9�Nn�z�N�[�?zm���'k�k��aw�c�$ �m��E��B��Z�Ŕɩ龂�m��3�́�8�:I*�:���;17�N�:�  Zg*��E(u_DmV�>��X�ݞꓥdVa{E�E27��q�\���ݲul:�@d:�� �m~5��2��I��n-cc���͎�.2������ T^>s)�Sc-��p�D 8i��6���dD�����QO��GNe.�<�n@ME� J򛇱�i)�Cy?��󑈿�o��~�ɶA���� 
z�9�������!Q���g��"\]̓��p�o��r��T�

/ua��J�h�]��4�
V�ط�0��8��
km<��	8��������,�f{�s���gT�x�y8�Z������5=m�k�,�o��i,�'/&Π��er���o&��P�hC8����̹�xv�Hd��7�ˣk%8T�{7��{ᴹp�=pN/���?��8X�T�y�����,��pO���0�@�k�R�l��7J�]�ͭ��i�٥BHs(t
�8�n�r"�e��8:�W�68ϥ2� �&����L�z�z�O��D��f�m��ơF�`xj���=����Y-\"?��.X�{b�P�@,�K�
��.�v��61�""��4ӑH��=��	A֝���Pl �+�Jl�����}��k��ls}�I�h�
�o��vk�3V6�Ƌ�!�R+>�LK�j ��T��y��Xf������9Ggl9�L� ��`)ܲ%��L���n�c8Y���ȿ��J����t�,r�K^*��L�5;���R��d�n�#���q�=����2����Kl�a3��7����C}Sك���r;����<���z��l��oH�
R�X$�2�����a�Q�����w}��\�oQ��L�"��Ֆ�����/?~�<I&����VQf����ꒇ���� >���:�Э��G�[z�['٫��H�ő�Ξ����|oɏ9vя�6�>Ų"�|@ccG��R��O!�$��V����ڰ��zc�?�$m��݅,1��Sɴ]�:�6ex��L�Tz�'/k� &S���#H��%��Q�6F��T:ə���0}<�Ѣ�4��̋����2���"��f;�:ެMT�dqJ������Ox������bpF����z�c�Ƚ��R��9I�9;m"cl��2��١��4���qM]9��5~����F6�mƄV.g줉�*�}����t=��Ư�>�SɕC���Z$�^����4����x����2X\�ݷ��%rb	������	,4�iDmXJd�SP�P���^�����{
}^MVi���'	
�*Y�=־��OP�����c׺�#�Y{��1	�r��N9���]g�z��z5�uc1�#d��:1��0��l/m���_�4�hGE]ˉ��ۊ�(-�W�\~��+�7z����÷�#~����F�s� @���>�-���=v�p��fa��ۍo�z��O�
���S��M���UH:A����(>fb8B`�Bη�Q^*I����tz��
�f5o��.(��J~G�.��n]��y����J�z?N�G��;�u���<��['��fOŌÃ�ȋ�D���c�z��kG
C��4kmE13�{�4�	 e�I����tEY�y�V�ȑB�~��YO��Qv�M�<"�N?^������C�6I�ܐ�F>��b�
���JA8gd�Yw�ЮFS͍��T����M����K������j��Eɪ?�C3ù��+r�mȝ1͆Q	���7�����j|�8g��b�;�'o�r5��������PDk8d9;��:����5��8�<$�/�*#�?�P!z_O�Z硾�'j�m�LI�v�c�������� )��D[�P�&��%�����N�2)p�NJ_^�9Ldp�w��y�|Ճ���WK�Z��KS�˙Qǅaɵh{/���/����&��ղcף�pu"���.�mj ��"d )D �X>0�pb)�{^�yj�f��B�)\��z�꣝�Z���^�9�:�6b�]�\ɟs �\��-v�	r�JR�����ǩ�AH�lZ-!ޱ_��p���-&��1�zV+O��3G�JD����IEq�>����,���)*	5�:�x"x^�TsÍl0��:2
�T�M�]#�§���M��
hQF�2�<�^����Y2+�˰�ԋ�9U���2&��e�)�s����z�9���HR��5��@�:^��Ӎ9a˧!k�?�'�������^�a}Yl �D�sl�s����9;D�_
G_!Gش�_H����gh�
��.�M�l�!�*X���F�bc�W,ظ�ӈO�9w4�`�z��Rd�ZN}(�ċ�wn��a�8B�$��Q�6�gY=o��b��Mdϖ�pM���y��չo(��W��}�y��4�&8:���[�wDϾC�L�:�N�86��s����|d'[u�ʝ,�까�f���>���ve���\([�ta������&�A?���D�4�Ew\ME^#���-��cg\�N:/�Q� �ҽ6������(p�)��������`��:ST�]ݯ���!VD%�X ;���K_� \��cB�+[�);A���{�h�z��Y��$���?�rȥ�ǋ��ݫg��t�t��#5Ѽ�}P��X���{�A�|��x�_��^��qO!�hR�^���m֯�b��/`=� �����+���g��6�#B��bj�����7s��0��=�;������|���"�JKQ:�8�D	S���?w/�@=�	q1�I#����p��8�x$�c��M�p?U^/��Dr�寰��wC��鸁�����4]d��h��:��$G�.%��_�-d�_f+�k�����.Q��V[��z>�����v�<��gKa=�ґ��zP����LYx�):�������v�����
uWAo��6l��dh�(k�+�4�jK&3���T�Jf}����m��K��#+��ż���9�����șm��S��A'����Kjn.���7��?"�:1]<��Q���}�"Ki:v(9�*��(E_`&f���(�Te�,��F�De�u��>b#��I)�}�6���:�-S�І��:�:[�:{�`�jrY����B�O�%üԁ�g�s�q��N��Ώ���a�s��?�	�Y湤���f�"�/�Uc����`�=��_-��zb{����|g�
�[@�=)��=ݚ/��V�0�e�HC�GV-c5����Ob}���9��x�	�ZR�#M�RPf��P������s�%�7�}U������$]mq0��n�v(l4p�?�a�
����r�R>����ۦ�� �/a�B���1#uXµ2����0��� ?�bm��X�:�
�cn �������E����������{�, 0����.�Z3hܛf�52P�M�=�B&+��������"D
���a��AIv�)��n:l9�N,��2(��C+�a�������©a�2��ٶ	�J�)��B��c*9�����rw����j��LZXs��z�a�Y�=e>d��\aaE�q5n�Wdg�J���k�M� �mIu�߁������g[+!�Gm��ӈ�bi��$dT�R�Y��y�����
o�4u��O-���&�v�E��kR�^��l[du<��&@��h�Ɲ�x��ݗ�{��_�X���Rˬ�|��!u�
K�n����-���+���wא�tqZ'lS��De�T�
���X���!�$��-����/++����ܢ�
+��������9�
Հ�լ���� o��&��z���CF�Iڙ�0����*�d�ovHC�N:>�m.�1��Q��� '�#�:�p�f[ Uc��I󨐦�'�S
����El�
��J_�Oﾡa����ŗTr�.�EUmk֊��lN�I \(a�D���(@�\k���\���5IN�LF"6 ��E�چ+�+r��z��#O<�Ⱥ��<�4��k���7���"�]���+'�)&�t�X��=,���������6q�`��_y��,f#�?�ё�c>D{;�D=k&���n�_�C (��9��@�"U�1��q�p�]Rdai)���/��b�kl훺��Z-��[�?�����q�T�pr�ݗ�"Ke�6� )�8�J4r��y?	N�9�����t���002y����.���ء�I��i_��\�2`aT�>}��z��nV�]S+��V7��^s�h��#]s'�Lb��S�F�zV;�_q��i-کK�I��4Z�KjXT�fs�كpk_��Y=%y�5�2�X��n���Z�(�$��]����i�����b�����ញ(����׸���"'2��KM��x����gt.t�>��Ԩ�=��I*�� Ft@����7ړ��7�c�=��C�l}�(��[�)����Jӹ?���Ek,��:��Uis���G�mҎ�Nc��#�4��$g��T�K�Dc��z<����5��T�X���Is�.�J^��MM���z5�N�l;�g\I
B���N���GS&[�,Pz9�(��i���M�O�pэq�b$�C��W0t�J�P9Ye"S+��G�Ff+�"Txi�v��[(|��Xӵ0{��Nr,�=�~Ho���/S����~��撜���_Qd�i�x$�d,n3~������e���/��2�����<<���3�٢̈����c �l�J��+9
z\N�y�æ�p4u�I�4a�W��M��@ j��򻋔w��L�L�gT��nT؝\�!��K�TmXJ�4�٥Y;6:��B�ԙT���?����G����Q4�U~8���>��"ye2B0�?��7pf/�C�闑�aZ?��h
�<���_z��`6.m��^)��Ջ�2QTO�E��xS�#{�a��=��44�<�`�ܪ���y�QOj糸�"BVє��d^I�pSyY� �Zx`�2TP���=>f.ez`뒌��CB��@M#D���IA��iJ��L�E2�]nW�aI��}E;J�I9/�BY���_�s���D
ɖ���0 �g� �ll��A��	���w2�HQ�O��%�/B2�,=���n���]�p����������b}���q���w0" �/���ZW�4�/����JeII��7�^ʀ\d9ݼ�Z�����Uc�C<DT�J5��E����h���~�+�A�D�.�À�{UYf�X���?O���Y����� ��.�,MN�6T� ���;sA���>�Q�0\6(R�`�/j���	@ڕ&��n�����.Ȑ���F�I�o!��B��4ms�����p�ņ���[��P[O���K;�N�R�&�% ��Xi�)Ƞ`͕�駩��}�V�i�
���D-#U_#����1^�������o�=��nxܖ�vz�/������խv��
~��9Sg,\�]ׄ���ɷ�[��ѓ~�w��\�bKK����)�h�(
%���rc���*���e�Cj>v��{�Ef�����Ц����6YzBmk#)��P+U�Z`���
?5=�j0��j�������b�k��TH/��Y�g�&�*.��W���0���u�Є�/?V՜��4��uB���$�0Hw̫�[O����ڰSS#�`�d�`+�zU����$=����)����ϟ���g��-'A�F��w
;�NRDl~g�����0�E1��;P�F\���yi�v�g�3���S���㻏�"�9��:��Oղ�it�iz�oD,�јrا��$\�膧aiY��Dm��+Fn4�G���b1���T����h1�S��V�g��D^��ت���~#[���g�Z-���5ۺ���qxs�� D4�@U��`�rҲ]�����`�Jw[l��9�Z�ńY��\n~gp��s��g����#
R,lbt���[x��>r��]��W���;��t�fr�E]k<ъ���ͥ�3�4�՘`_�x vNp���J*��j���1#�+3�����'����G��9��p2���RQ��o��堖���1��W�B^6^KYE�N��࿯)�B�uzM�f�0���u,5BS�7�jR~����Ӯ8@bK�6A~n�Wvż=#yܥ���,������Ȏ�2���rYvdz w�7���fl*��{2V��D��E�A���h0*j+����!&41��hP�ؗ�3�$�Y;Pr���ڲ"�4[~1�\�k>�� 2�o�,�X���8��?D���^9-���v�w�����K�+B�l����$歸a>�ԣ�m�^L0~�R"�b�R[���9��o�*��-�o:.EQ��U�>�����7�9�OM�-���m$I�SB߾����
�YU*��;���DSی�g�+X\~�$�
�4C����`6��mU��}�A����Ā�R�Z ��F��+ߥ�C_�c�b��/D"����m �7������rCq?��!))	h���&��B �.�x��eci�Q�q!��f����Jt���AK��F��*�i��(�����	�OT0�^�4E���E����Wiu����r���ܙLDbM;�4$���0�T�+( B��Ǟ���l� �ص$gbBfx��:������GǦ@1�`*!x�H ���"`�7���F0��4��2�w3�Ԝ��u�W�;±6A�Wm���y����K}l/(�(����H-����{C�/\"Ib4^�>����T���W�e�����p��&��"�ԭ� ����C .�%X�IٲB˾+�aD��a��HG�i�7�{�Q�xh:�ǉ���=�D�F���b���G�@�kG��)��Q��u��?���������3+�|�>���@�9�7�'�I�J�	S�0�"�ɱ��|WBl�� lp:$�)ln��c�FԎ~�t�"�
���;�(�	]k¸�GY2��qN ���)m�p����d�Յ����1����eB�	2*�0��ZS�a��Z���u�-�qCs=����Ҿ�����*]�VT�~����rj�(]�Op�(K��2t�1�D�.��nŬO.z�XXʛVƆY2 ��߶�w��!�NUCb��8Њ7����/v���c֪�$�q�h��b��X��W�Ӱ�p�X_ǆ�a:9ܴ�,]4�5��E��L�:��؏s
u�H��.O_˗��{���T+uI}�-�(����$�Wz���cq�N��uC����h�N5�N^��7���_�9+`��v�I5�%�}���$�sPu�r��Z&�t>��D��>	e��W����7T�*������=�e�<6a�Tx;!�H(�E
揚��]u�+G��ޏ�F����fQI��@�^�3H'M�-*KL�0�aT���5���q�����~v��[��ٹ�����T���� Pu} D@5���r-�J�����f,QRY1=D� ����b7ٗ�ԅ�.�{��u�õ@�v��_��0]���b��:���|�L��AҲ*GMD�>1>��#�GiV��Z��W*q=�˘���Z�ۻ���"&�l0$�����d��Sf�L�1�C!;˩��#�,VV�/��v���",.۰`H�G]fh�b@�eJ�y�-�܁��z�yӾ��1(46[E�A�^}&��.����t=D�_]�7lҾ��q��F/��B�B^b-�,9k��`�iTm%#��Ǔ�l`z
��!�mo �qE���n]ثw�=���q ^4�H���1X�l��8'ɳ�7os�KCH�V)KI}v�	>���b*����:�ܹ��
�7�ur�����7f��1�2	�̬�>�لvK9U�{o�u'�^��ܜ�ulŰ.o N�:�}3�%����sW��O�[7]S�ԗ��n S�Ko{���x�Hٗ��#��� M̟������%���;A����r�*�?[{���2��߮O�5��*��!?&9=^-Œf�3��֡�`z{����%-9~��_����x��
�����俪Ͻ�Tz�_��8[RaX,9ѡt����(4\�%�a�\>�4������7�*Ƃ�� U�v.|o���zJ��Hp�PxE�Q��'���p$���;%p"���A�G�M0�$Ud*�KSK��)@�D��c�c�B
-���C	�!���r3/�tF�;式�a��N�bW�Z���=�X|sdg��YDp(|qk�V�& X��OB�' ��}g+���}�.��x
�"���%�P��$U�'�AMC
�_�/
�D�:�m@�YI�u��	w�_�<Ѐ+�I�M�!�i�ȶ�������M\!��������o�Ҵ���!��h��0��c2{
N�:���&min�@�6��������qG.;.oӍ���� �+⍖R-{�����v�A��h4c����Z�@CF���ipZ	�v�>�?��������N��xX�nA�B��y�	)D�z�Kx�:�]=g�8;��&�9�`�f�z��������q�#|Z�iIw��0]���z���.~����tt�-
�����A��Q{���@hA0����<����a�AHir|i�H^a���-kܖ�M"�X�Py��l��2[xF�Y	�j��:�n�҉ӿ�CFYD[S?�)���]�"-Y����ŵ9��cI�]P���C��RNM<�*�=�[����V{bY�)qG��ǥ�b9��S �s"�P3���0HRa���������aQ�L[<�{WaMܯr,�x��Zc�@�J�A7.�h+W�q%Ć$g��Ѓ���T���S���q��ve]V���R�8Y�Iʴ�y��(|P���0�T�[8�g~.�y�y�C�1�n}Gʻ��A7q�NQ|��=�q���]/5sMQ�+�8ˌ�~*ĥ�j\�q���z�sB�j�ʹ���4X��O��ԩa�W���'=F�_������K��pz�`�'�Ӽ;�N�PF�������;a
�Hʡ�-kV�_��a�������듓��3��NW��@.��M��Vf=��L���G��+{�[�گ��wW�ºrn>W6Yܮ�����2,I6�Z�.�C�	&���Ca��C��pҟuB�L�7��j�d{ �_��JM��-�t�������ݞd��	L����r��#NE���b��4r0�bX��6��F�l�ޫn��Nb�6�dޔ���|�74_v)�W,�5%h�<-y:}a2�<���si��;�"t&4�����e�i�1j��~�2��aT��V��X�M�	��MA�B��/������T��*���b�v��*�g�vR����@}0�})�)Ř����0rA���Vfw�󓿐��FM;ͣB!�
�y��KYl*{��pm�n�a=܅z=���'�D���0���`�Ĭ���!�չ��XjW�.�P��(�{I����4=��fI�\p>A��@܍nYZ�sS��H+mȓK]��j��F >0O�#J����ܭ^�D�yn^j�?y��~#�Vo�'���s���R��*�A�<^���nQ���3�w�$�#܏�J��i܎Lx�}�g Su�7����pK�}�o�\���Y���@H��?A�����(X*pw�݄��� /�U�#�1o[��}S�K���t'+6;UCq��%�:,��}x��<Kg?h���0���Փ�gqHRBX�q@���@���d�*�wz���Xt���\4�����$�;�H��;&�i����켥�?���@.10Jpȉ���8��)n�k�O8��J�;;��\�kQ��
<�ND �H������?���w���:mҼ�Ԉ�E����!����<qrm);|,�1���g:l�j�_�t�@�!�3]v����&,F�ź��Bdul�o�����T
�+[o�CK(py�Q��mJ+7b��"����v@�H\�������D�`I��ɡo������L�I�[!��ϖ�I�c�OE�,�c�&4�W�T<l�c'>���כ�Ҧ������6��?�y����3���ZM��,zM�Zƭ�܊&L�4HoHj
$��H!s�XQ��|Q��ޣ�J��
��R��lV�S�ܑ�(D�;�y�[�+Cao6R�]_h�=��.���9�M���\���"�Wʄ�*~�z�{k}�
&�Ҡ�{b�8�탭m���ӣY����o�*��d�%����ւ0�82�{�<n��UP���������z)�ut�ΚFo�H��,X���ɂȁ�7��\�V|���Rϰ�y�]Mr=�Ms��yjQ�&T��l�%=`��1x`����/ǽF L9 �$a�t�U�:IMˊy���A�����F�S1��=<o����a�y�pv�]}���Ӫ� ���X��OS
���ќ	qץ,��ȕ.��E��2=�lZ�%� ��`lU9M܀hTڶ4��6�<�2:�f�����W����_�gGgt��!��W������KCV:�q���E����6�����|I����j,�`M�_l��i|��ױ8���`S �峲�k=��� ���e�5S����R�����|U8���DƋ���]Q�⤉��%�8$� �W������A����1oh=��>^;
�E��ro�{F�~�'8��St��Q$OmE$3��!�l/�G����K��a/���g�������@�wP����e?�tf깵?���	ғr�o0u2��kp�A9{Ⲟ�ĝ�\�Xpq��\�QJ�v�_�C�������ؿY#��rSW�����ɢ���Eҏ���j�~��Z֧�{��2��كM�V��"�य़DcR��p �g�J��
�9w�r\��"���vr;W��V����"�GW$Rs�����Y��=B��F�+㡺p�S@~���Sd�4����0��6PVA�[�~�]n�o��F'�-
O��s��<鸹c~Y��՟zܘ)��L�!V&�q�W���*�����l��׮Q���}*�J���*$`�d��M&�~�u�З<�̟"�2���� �k���w�T��%�G�%<!��8�K>2��Qe�l�~zE&iN�ߏ�f�o����-����u�h>"J!Q
���h��4�W�3ס����矾-4j�����-����"��������/�ǊY�8,���o�]��:m���[��K�18��dG�o�:�BR>:P�sŪ�p?IBO�_��8����@�N к��vHf��ԟp�[�r�M%X�H����!j�+Fõ�*�B����!�Z袣3F @|��7]� ��ˈ�	W�g!��}X�Bfg�F�pO�R ����)�f
T�30����K�F� � =9��FGL�� �O�I �8n-oP`I�1�(�Q=i�9��ϒa>��ӮZ��8�m�Z����>(�M�s�������.0�,�p��1e��%yK��c���{�s5�3ϴ��.B��h��i�C�؏�-1��Σ����^i<3Ңb�o=��},%u�W��h �J�cx�����9�y\�*���+�Ƭ��@��dc,�"�˫VWz�p�jlʮ��AcRp��bFu3�f�+	��%fhNLW0�Jd&�Z��r~�ឪ�?'�|�	V��2qȚ���ř�j�V���RI���C�sdtRݹ�̤j�f�^�3��G��b:���BjR�Y �aQW(�]a}1]��j�	Z�O��F]O������t������RQO���F�=-�Bޅ�a��r�_D����f��gr+�9��6���_?���Ja�`F�6�%A4�j��r2q�+l�x�h����)������Df��د�J�0��L"��f�r�0_tc(��?�0���b�S2z�=6�)�_ؽ��3�NB��z���R 1R�.�'��ю���Ρ������>����Z��l;��{����0-�vb����J�4�y�3I3�ɽ#�@��}y\���X�����s�m���L�q�����bKt�GV{�\:��R�VoU���NͰ���-)je�����������cϾN9ݭ���h���K"0E�CA*N����i�F�:Y~[J8��a���Q+�tͭp��q�2���Q_(,�cQ]'�F}8�ϼ�Q�s��	K�^�ʤ�	'����؃�P�\����y�M����/ϋ����αK�O7��\a+����d�B��k������9�|.��z�%	�I�����s�g ^��_��0Ѿ��=��7Q��R�Bv��3��A����aR��b�^O�U��8�_�C��<'U6G��4�ʰ�bK�=Du�*�.��̹�+(@7�.8/�&@{2~?կ��7
\Xȯ���_�)�A���f��DUw\�Y|��۲��N�O�Z<6�7���q���r��X�)M�:d�WlV ���mT��V=���v4l��
^2:H�k���7�W�����7���?*痦	�u��n�\B�������h��j�N�Aן�]�གྷ����;���yH��
�=�#�=�D�MP�w�<��~�z�:�@������yĦ�ݼ�\?��g��QK��^�ȏ֎w��qN��¢FY�8�U�(f(�i�jV3����N/�)��W�֏��ֈ�3AI�	�C��hq�0#ٰ&��H��-TSB���eOaB@�� ����`��	F&���������C��Y:�2�����w��w<<f�4A�L�����H�E)rW�oN.���r�1�pVyJ�����*b��(GN+�}(0�,K�L
��v�Qe,�V�ZGX�� m����:�f������M&n�8�T	L��������^��vAP�/�$���?t i�*�i�H��`��f�t��١�i.u-���[%݅0)_�JVoC�4���y�U����o_���$3\�E&Zh-2'o¾�zΦ_؈�\m[��˅<�?:����R� n�� ��K|�0x�'�1;���T���(xLʭ�ɶ�Y�_o���zqɕ���~����H&�/I^L��;�܌���x͖ؤtC�9����N�0��b����xA
-E,�A�rཟ�2�zf[�al� /�4u��'ÿ����: �/����5���W�����q.�-kN���o-
�٠�oQ��ta��>�S�`��;/�xd/�Ο�]|�d	Mv:��X=蔿Ƣ!�>�R#�W�>{8噽��;���9؏���+^��y�r��Qj����U�G��K�6M�/(`��Q��A<��rR$�r�z=���7��1�#Y:M'�Y�mBj���"���(Mu����V���΄ekVFa�5��S]�K�̙���{�����:�nI�d+_H�j[6��H�z:��1�����߀kCN)ޑ*�ȳ-Ehc�����l^�Y�,��B�W�f�s8�{�.��5d�O�s�#����,Y%=*��® i
(�<&��L��m��X5�AJ����0l�G���4dy����l<�����lB�0�fIʋs��.��Ḱ�A-t��;�;H�5�����eIA;�����8EZ�6�'=�)��Gl3[��$�Q��?�d��o��w��s���ރ4�-fX�n���Z�_���=�tPn�r��s�.#�x��y�ʜ��G�
ES��m�J�����m6#]�.�>D�'+��_��:PQ��
r�i\�h̿�Ù�j����[P(=i^���uB1���Lq0��V��&ĩT�Η��B�8�F�ZD�p�K2�b���6`��am��#������ɭW
7H��m�U~$<\!A�������Ln�e
���Y�VxGt�
�{3���.*l��JUԌ��b�l��� ��C/Ҫ�����x�#%���ao3����S�H`��-�@I�_�d�wϝ�;o�,'v ��7��P�f�s#	��1*TB{�	\
)a��T�Ƀ�nr n��	vtZ�5����cجP\�����h��@>tC�E�V��!_��ܩmr�%�}��������ES;�rƎ �ɏCz��ወ��ʎ��,>��;A	cq�k��z��!j-ބJ;���`r:�J'��Z��J/q�����_I�ekH2���5O"ٌ����).�R�2�`V���{X�38B/��5Q�F��q�Gg:�^u���zш�juau���rx�wx��p�v̯���a�Ѐ�5�d0C̓��k�3������{	��� �i�d���e���ߓJ=�x5ϡE���(�Y���?�s�ù\x!�U����0������䳔Z�A��Ff.�'��x�7��pd�U�B�&�yj�5*L৉�Q:�L1G�dڃU f�~�|Z���Q�3�̉�"O�������(�$i�"�b��ݪ�J��2�=rD���fAq-�g#3�H�0S���$
���Y`[o����	�&�i��XOd����(��n,��v|v��3QT�{[�i��b[f�[0�($��1H|a�	����GT�v
��خ��� ~�@$vH�K�R*�H��8B;i3�ބ�|�A
FK!���?��d��D�3�`0��=����k���$�N�(Ψ�6�	\�q4��o������-��\)�,7m��R	����S�zi�
��@P�̚��.bt�{K���Z@w�;;Ȁ8~�0�$�/>�Z���k���l�>wΪ�!:�Ϥ���_�����@0K�e�8�^Kx?{,x5]e�5���A ���y�&+����晴�i�KX.Y��p�qg�a��d�B�ȭⓉ��`c��j5Ai�m����e�Ti��z�}E���NZJz�O;�lb�����IK�#�~�6r��py��\�HMLg��B�}gc!�c�:Rܩ��J���)ȸO,�3O����y����o�Ԕ�%��A$s���	u<�NG�� ���F�ª��y=E/ugi)ˬ��r���ugi�q@��{N������)��]������b�,�@���������S����w>��&*�����	���G+��S�%;���t��ʽ3s*�wp3�5����Ȧ�۠�`Qɤ��g�^\�p4u5��𺝠πfN�tŕ!�K)9]��s��=���+�M���dY')�����nS_wS
N(#��36Q��JL��X�q��w�Uo��i�I���`����1�6X)6�*��"B�oP������sNT��&��xY�x�N��,�Vs|L����趂�2�l��R9�{����79I,����3��@�n�>��m�<�auw�5�u�6�-~c�^������r��u
#t	Wh���*�@�w莜ۤ����=�	��eF{���bS�� 겭*��fb����s`A�,^*�g]�maDD˅٨��e��n��&6:��� �Z�4A��^&����޴ܖ�%UZ�8"��	�,�|����/�rQ�fm�_^�X��W?	
��==$tw��T'=�e�c�3n�7׏B~��6g��C(� ͐�MWEc*y	ةt�w�7�C����|NօZ�-����
n�_?�ٲ������go�Jl@�������A�N�j��p�y�w���D�.%H�K� n�l��]����kg:3��\���6&ʜ�����s��Y���;�sI��F��[h�X8yz�k��x��d�6Y�w1���6\��;ɛ��(J����;����Wj+����{?TFztU�+4�ñ�jaW���g|�z�>2mf�������t�o���+H_1r�TE���oב����_�%��*׋��K&wPz�H'
z/�.�~�mc��[�8�'�Yơq��i��-�O^�j�AR�Q+�}=@��O�O�M5^����C�s�8'��u�'IW����k�W��6y���8��Ee��g"�y�gܥ����� �Z^��4�s�q`"�ŏ�r�a��~ gc��y	�;�(�8���f�n�e��+��f28�ؚ$3w���w��;�ů7�Qiv�D��������� ��ί�]*|��V% !��#8��8��1�،t}��L���<��Rx&��@�ޓ�;pΔT����$���f8������B
���s�Շ/�ߑh����z��ON�ո��^�=�\A��lcHX����@���	�զ��#A�ꄷ�&�#!8����g���~�u�[��C�� �O6[k7* �҄h |[�3-1�����Ӏ9d��E��4վ.5k�?�Piz���V�4/�Lf���.��8o0sPIy����Wa�A��o�����c��.Կ��a����g�L�`C��q.��*ޜ�n���kc��+���Yj�+�ɹ>����l�s���x5q��=�*,�/c�W	�����'�ի,鵾�
�ZO��V5$�܀{YkU��hR��WN3�s)�(��KG�����p/���p�PFѱ�bKܔ��}��W	�h )�ct�a���<A<;^~��<Ѝ2QU(M^��l���M^�kS��=�)���E���8�\[@�Br�[��M�������� 1,��2�eED'����/t����@����6��������'�G���Zb:vO&z�W�Lr2�>>����ܔ�+0����oL"��J�E���㖳�☉.iaƳ�Cɫ}*S�i�53>������D
����� +64�Oq�I>����aց�ۖ��0?rb�c�`z����8x��MvU��� � ����8,�E��P,Z�s�F����d�H�͇�����������?�V?���ؤ��z�%�@
���$3˽˰J��H��zXߵ�/�h��e���/u������|���.]��fti�(�f�_leV=��.!{ڗ,���Y��S�P�e˪�9���':n͜�O�A�	s���B8e�$����t����O��Lk�@E7@9$$BI���g��{����ǜ� ne/F-b��x͂L���}"�=��U��v�kd��P��5P쉁��w�[S t�!�1Y�聙-��$Z=�`b��h�~W^(~���.`d�Z�����S�z��������%-�hQj��u��y����D���/<:*�^��O�3~�*^B��?�ُ�]��2E��<��W����ͱ�
~ђ�N�s���q���w ��� �Prw+C��� .��ZiI5]�ڵ羯�y�Xo/-A������ꖺ��P�G0�s/G��Pz�
N�,�j����霢���A|�l��x���y��w�K��,�˯{E9*W�o�B�E�o\�!�R#����G�Q���ݺ*�܆m��^��oMa���Ǯ��O�Ր��DH�
p\�(A;S����W9�~cA����k� �ú.�?{;�\���Ԗ���&1/ڪ�6�RǺqm��͢�{��?FÖ�ə��+� ��n�mU`#����mf�8��#g�x��9�d�v=�>C��MBrh�]���K[���]��H9q J4:��]�i�j��W�Je���wg%���a�c�l��:�}u'��U�	��Ci���Ή�g���uڌV]xP���I_�d�au`�V��7�k����$6���y�gd�%זe�]_k?*��bHR�ٓ�X/�B��(� (ŏ�t�����N����C�<�N�
��� �#Mv'���+�FD��?а�َ��#<`�{��[����6�h�E-f�O΃�`(/9�G�\��M��x�=�=�0�w��C��S�1��v���'mp\j�����@=AX\��Q�q�e>W�kr��{r�6O�q����W)���}��/e�C��fe�@�DG���}�ud:��x�R�eO�
�~���S�TӠ�����Wnh�4��o�%\�/�ö��6��q��D/�����s0�r ��� ��t���ɐل!T�^^��>��c���H���y�v/�aZ�5j8������rU�`��U����Ϸ�M���M��!���a�Y�bG�5����d3�^-{����w����4*�-W�;8!\%{�cE#�s������*r��h�l�ac{���Q�_
�_y
t�Y��cKo��� �8�FT����B崙$Ê�����`(!ڑxc�wq܊5�6��s�U�81X��ݕ�{�RS-�Q�F�jz���/����i�yz�)����c1j�V1��Td��,
@ΗT���\jm�>�H%���Pg��M�:�yuR��0-�U�o��-+��0�����Q��y����fx���Ge[a#g�!	K�Cɻ��Qؽ��ʙt~�Hg8Pa8ʇu��6B_���ҿ�'��O̮��4����s3C~�~=cV6����ߝ�B��U�o���2`zP,[0���W5(~]�J��h Ah<C#��DEl$���푸�6�A�p�MW��\�fX�;I��˗�`+$�Ĥ`�,��J����/�aH�Q��eʖ������,Ȅ���c����,߾��U��,)wTkL�6��s���Ģ�&ʳ��s�c
�77��}�ޖի_+ ܄��sfݸ����u�`�C�й�=v�8�T��%��N�5��hN��I��an��}�A�u
$p�i�¶�o��'}��k�_�wf�yp7����ó�KLS�M����x�t[#�Ԧ��Zd�4E�J>��g���!v��$�]��ȇzJ�&Q���ke���Z�*ϔ@�����IG�QiB[�xE;��TS?R&�Cn��3�N�Dv��� ��T�׶ʸD�!C�;�88y�&\/���?Qٝ��D�����غq��� :G��(�Μ�%�����(0�ϫw��ƈ��bj��=~��/FGS*�� �l��&${�|��H�|oݢZ#k1��Qa@cL�\9�/��h.q.��3d��?p`�F�[�)U/OB�E�3Ԋ���{$��� �G�2��$gK_�t5�4T�T��x�z��;Ha���*pu�~l�G	}__�$�H쟶��NB�ź����L'��7����E��_S�gu�44�����D��r�#l�����ղȧ�t�(���c1ji[���Y;������[`P�[,����/��W����(���vg�N��lַ�ɂ~\����ݥ��q�w�غ|����Ojj��z�#���{k5�AO���l�֚D1��0A��2aVe�R��l�ͽX�$�^�W1�h3��bW��O
�_�,��~�K�xh ��r��plVNf�����1G�f4����,ID�.��P�y���u�)9=�5��N}����dwD|ef�X��X`^��ʖ�*�Zu2�_b�J/�=��;�~��O`Q���		��
��}���.�jS��/���L��"'�HKy`
FI��9x� ��3[[V/Ϻ�p������g�?2�����6�i7z9%�h��2�go���(҂��_僾�BuD?�%gb״5�I-8��=#��c�^�g���8<x�^e�8���Rv
�5����m�tb�8�qH��cU�������X�䠉1vNSBA���~�����97���	f8,dJ�iRf[	�烖��NdW)��2�K�
؆�:�l�#n��/ԯ�z	)���l�&f cE:���6���7I�< F��4BI.Us[��F�7V3�9of����nբ�L��͝�$Rٟ�;����/lU�9��ET�1���}b��wdOz��'�Y�tW�_0��:5�mA㪝�ԉ.J���5\|���ӟ�d.�����?ߠf�v�%B��>5�qˏ2֞�|����L�D��l����\�B����GB����{/�D��LP�g�u�I?�)ǅ~��f��4Te;VY0c.�vcep^L�g%�x�HY� ���Z�����1.�v�����2�j*���ը:��׌�չGH~�S�U�º�e(Xt����g�X`�F	���RB
~@OgXdw��r��)�����Z�N1[k9�/E�;�D�^n���Eb<�oi�4���7 "^���J�X�Q�m��=3���v�T][�t;�fLl��g�r���K%� ��*/ �ʹ5i Ks.�r��n}��e�P]kT�I��NrM";�	K��1�𢛐�"�PEP�z�>��0�#:$�,c�z����۰?@j�n
#g�L��ۤ������m]K��/��#�g��ř�>��h�{�T�"�=��R;wl�m�H''u=v�S�F���w7�����jw��lm�OcKd�W2�{@B������(x�)��K��ܑ�*�eR
��j6=RQ�Q��!�������"/7'�m���p�n��'s߯3_]r^�Nb9m#��߷��=2����c��N�/j�yHbjS\[�1ta���x�Öc��(˓�d�N'�ƌ2I �����?R�)���I؇�#�I��촏��f�WC�UH-��sA]Q��>�F�u? l}�9W�p�flW���R��G��7��6�6��bO2�t�J�tU��I�1��Q��� �q���rbn�f�к��TO��&���M�)��<�dn�԰ ������9�ȉ��<a���S��t\C�e�Ai��Ŷ�l�]Y�Q¦���a8�}[��<ߺS$oyqHd{g����F��[��#�?�w���&8u�s�/��d v�6G|�e�qt����Q��mdP�e��b�hR�0V��څ� N��-��ve�0~w{�҇��yږ?������.�G����`|]C��&������.V���4W��P��J�Ԭ�D�s���)r���D�xI��4㭖�a���U�)��Q%:��J������,8 W�-~�A��
�Xp]+ L^���sO��t��돢,�9�-T���:�Q���k��~�I.[�����+�$�ڐ��.�cdb��-��'"�߽�
�����]�|�W瓤��C�ӈ�`�9�!�Fts>��c�R��icr��m{VV���UÂ�#���0��Ѕy�U��&�h�#p"X��� X��ϼ�jv�_1,��*C���݊6.�"�z��>�@���v�'ܷ�"�yv.q�E��1ڂG��C�c-��KN����4
��ͪx�@0�\Ǳ¤f��4v��¨$չ�2�� 7n��hH���3�V�bo A�:	=���j>~��dgn�$~�!=�r�c#"�M��E���b��'�|&:;�m8J�cd<^eĜ;�m	��.�hF���Fe�B��zA	���d���1:����}Z�.P�����b3=7ԊW���9�W��I�ǉc*�����t;:�~�����A1�D�Š�4)�[l+ಹ����x�^|	yO<d5�(�"�,�6N�+��7,�ZZ<���k�M�o@��&�^��� ��F��T���<<��mK�o���cQܪ��;��o��	&$~&���ؿD�����oJGӸ� �GηL0��D$Q��!~�޷�l�j;'���[��ͭ���5�=�Ll�z`+������l���}=-RN�c��ﲳ����Hʗ�z�V���7�dj� J:(b��Ty'FO����ok�:%��L6L&7�L�g,
3����$Q9�A�Mk�	��E����-�/�:�_����|"�m��q.�w2
����
2괅��M.��%d/�Cr��<�]���M5�3-��<�-j�Px���l���&T� �!�u��0�����	,�K64cO�x�߇��5A0�Ad��{2]H���s�+���J�y��t���6R��o둭u�(������g�t����s
�r{v"�T��v( �`�eT��Y޵�P��b������P?�uT�ˋ�ƪ�ԥ]��n�������l�E�j�1�Ǽ�Qn�j:�Q�2h��X��$8Zy��=��0����3�+Q|�ߐ��=���Tk�p_�������c������2g���,��ͨ�'܁BYS��X�|>|j��,�&�B���jL-��(�7�f"L(X�t���lc���ލ�2�^�4���lH�oM\�(��NK�dz܍�]����/0p=��]_��F�t��c���N���S�=_���S�� ���B�����{��t�7�6� ��j �a�P�+�7���	�.H~<��>X�p�X'��q��i�n0}�e�gE��r$�yW-�M�?J}����+�ɕ���xNjA{���%�m����@]�Ԝ���	��1�6��B^�d�3>O����x4�%]9���M�i �����e4�8>�lQ�����ߏ��&��|O���<��كzI"�0n"(�ν���~^�?}��X�t�a�>�l4��*Es;�j�>���������K��T���a�E�Ի�҄��FR|)�V�h�n������k�;)������1��;��!���<~����M�%�]�J.U�_
JWWj����c�3��\%ak�4".Ϳ��,9z��_�eeN`
�`�b���9��n����`��1p�A]�xl�8&@���m:�{��z�~IC[��x�c�����r�������t�X.�_-�o�K��]���F�ڳ���J }�Q�0T��0m-�j��1<�dŌ���E:jJS/!��mc�A�VK:t�UPЍ����V�ٖ���(���� k�y����v�c���#y�N6�~q� ���Z�ݪV~��EE^ⱃ��5k{*��;�ρ
Cw��)�r��Ϻ|	����EL8{��G�p�mHT��ͨ��/�gFm{���M����<�h��0�&����["��V���E`oTW�9��K��[�#�{Mr���J�v��8�#��B`w�c��y;_ހ�-�j��b%��1	^����D����8:E%�m��GF5a�C��匍!�����c2O,�6H�jb�Y����i� ��J7�8R��
���D�YHB��S�2�au ��SÀ���3̢��{��sz��Q���䆠>�fU�
�ѥ��u�0�>Y���:7�Y����nY�R_�4\קS�<�=D(�I�ّS� ֶ@���pZ㋹�3+�2�Ӱe�?d�>j��Q�\yRJZ�F7sP�,��QD�R!{e�����
P� ��'ԭV���Õ��8�	7�3���j>\��d�y���V���_"9UI�F|f�D�������SDJ��΁�"�i�9�;�k���z�(e�Ä�6��[�_c½o�?'1e��;p}�����8Q)8��w>��3o-�����U�+��{Ϋφ�3	o��"v�s���6ڂ܏J��<o�'��h���c	��N���7G��N��⽑�Cj&P�;��>!P�f��>�?������>�f��c�͠ڵ����s���|װ4*s���'bEP誇�ݟ�,2sayz�t�x|� M��X�sIn����(�M/���٣�҂-�{5�F$�@q���d�$M>xC���rC�\�l_���)uR<�!^�J�A4�G"�"QP��+�%��g�hw#E4����[6�$J�;�}�pVU���X���B�����|�V��9�x�.��/��r�f�vs�gNL�m���~sG�bI�s��y�<����C��qMҖ	���C����Q[�Nd�b��8���p^�ᕳ2�pr��-��ל*�IO�X�3�	�Ǖ}�IP���g�.f�q���7;�p˧꧎�j�d�/�,+�B��z�}SR�D���*��R�&�ڃd{�&�C�>�x,9�cx�6��\^uQ�5)D�<H��/��	>
N�����v��$Ԑn�ށr`0Z���+(�f�2#B,�6s��S*� �*���`w�ib��o��:<��a����2�����P:Գ2�h�S{d.JH��<��[��5����ޛ��B��4�?�!0�IrU���U3�
��J\XA{,%������GD�A�BxU�*���6��vW ��(Ms`*=�����U�L�ej&��8y��1�o1æw�[�{.ϭN!���(�yMI \֌�'��4C���W��"h�A&�P�A3�k�r�%�n�l����n[�C��k�3�P3��NsK-n���:��'^���f֍
��)e��3.w��N�U��C�l��\��`��,
{���Bl���zV�����}�_�!ϧ��XN�4�|�����ؠn��"`��~�5�q,�^��n��i*�~�!�����*"�[��KMS�}���z��ɏ�E��h�}�UE�Z���OO4�:csf��.�2��u~�7b�)�|�/])�JW�>{��7"I-��Z%���3z8=���/{��
FE�a�.�[�<_:���`q"t{���>�Z����#\Y����uG��8XCu�)_�!��p�����v`p_2����0�!��1\9R��$t�kz �j�
__�h�M��h��a.�y� �'�T���o������e%�S(r�uٱ���tc�Q�G�6��}9軸�Su��R��X�h����aqA�s2^��\���VC��vy�a��66g*ͤo��Ȋ��c18��pYa�'��p����UA��Vmc��^�5X�U�ɣg����fӄ%�0�OO[�����g`��(�ؿ���џ�ԋO�rp�j����LŅ�؇��w��p&7��D6�CwV�|�x��U�a��`>��g�iWr0b�)������s����X�*���?}w4
�S�MGu�Ƽ���MVo����l�Pվ�u��@%X�m~�א�&Ի�w��{�_��C�r�DU�T:�$S�ʢ����SR���M��"���QZ7�+_�eɷ�C�k�~m=v�;�ȱ�k��#/۱�ȏY���դ��fkD*�=�����x�6"
f�����RZK���p�X����?K�O��)�hQ�7(ǳ9�F����B�	����a核P#��Ly�7{��iFe�+���&:�ڔ��Z&t"H�=�9h%���xѕ �ϭ'g��=	C�d	QVv�B�\�����rV����p��h���i�J��$�#�C�ߩ���n�؃D��I������${�P��$���Dh��YC��]U(�y!���+�ﯿ��	w�L޺���yԋF�w��ןE��\�2w�IxVIt��sG�2�Q����Z�5�l���H,��('�9��Js*T�,��!��Ѵ'�a,B�녠���cJ׳�����@����`��`��)!�����6�&��.�skN��a�*-�i@(��[��V5l�7̭rs�r.ާwt<_��8|WXM��kX�#(dz2c�Fa��=M9=�H��p�[މ�5�YuQ�v��:�@Z����ѓ-�(��9E�C�0#��8=�}�t|�W[n�x:�u�\tG%�����k�R���LE��nM�m�͑G/Js
_�L��R�ڒz��a�Y���?!�����
{����d���(u���Mw*tO���_˳v����ޏA\{���~Y#��j�T�W��G!����2aC��*�^\�_��<]-���$�Z�=:׷S:kq��'�/jTm�;�kN���?�S\�/��f>�BF�'��Ft��)��wI]!�k�k�P�cu�ȊVG�J����>����o.߇a՝r@����r�ˉ�Icaxs���-eA������ 
���7�0��K{�Z��e">��(W�	�5+y�K8Fp��OB�W3��}ܴ�Ж[�S��'J��a,��kC��qP'����|ZP�s�����"~wP&1ۮ���FA{�9�զ�e����mF��inN-;�!���m)�Ck���1W+�7:�M���*���M��M�����kz�<3�@��4�[W���m�`X>��u\��6Db,�CL���(��sa�AE�>���w9�ߙ ����M0>&q>1 ��S�{^�E��J�7'�O�Y�w��x)y�i����:��bZhvս�rg�x8 k��65�6˩�٩T��G�n)^N �� ���U�
��h�4O>����=���G��9���?(M�*uA�ߋ�:z�l%=��k��!%����tJߋ���"
Ƹ���7��Ç�yosDt�����#��lT~��ۭ%�S����G�6V�d�6a|)^�^yMb�$�����ڋLV~Lw[�a��� 6�־�a���d�r�D�"]������^�]	�ҤZ,�"�mo��H�7���#�V�x�MK�/�҂��ҭ�BTM��;�Y���H���(������a��D�m۞����o�Ж��/�m�I"�7ήfmc���т��6vZ��Եr��s1���_�U��V)74-{p;|�P���2�?B��|m���'hp\��d|�ͅ��P�?Ḝ3O��$+��݌(��a�;s�>)���$x��*F��E7/T�՞�1h�RG�Ч +�oX�.J�С�S�5	�+Z�O�@�J����S��K%���b��,��'R�EQ�쁿'��^�q��?lǠR��gF9�
�Yô��*�k���Q*�5UM3���6����f�����':}���Hux��1�Uf?*ؐ�/,�!6��3>�(ՙN��1cs�Xv���z�Z�td�� :FBG*�/�W��		���cr[���j�,05 ����1����x��I;2a9�����7�[���*�5����tn/f'��E]�:��D�\BE���]� *}�bw�#�F�Cl�]	u���=�	�H&��z+��ˢL�����0A��	����|�]&�g��N@�Y`Y�ƒ[�(���|?�rs�G� U^���lF�p8c'^y���?`��<F�Hnz
��T��]d��Y��ͫze���E`?��ӝ��(f����/�f:�o���[�j<�z�+�&rѦ}>9�8�Ԉp�-G ����e.�9�v�isf��>Ʒo���KB�.�]��!5��lx�%��s�H4��"���aɃ����Q%ȤB壘nD�����p��+	�'EyCʽF��@���5��N�����͉��a��va��V=�g�����n<\�~_�9�����3������-�Z� /	�0j��t����bA���.�a'�j��k�^h>nry�4����Eee(���cA�����շ �nOr�?z�W�T�QeYL9��v�����go:Zyb�]U�\�^>�2-�Imq��	�}���i~0��cX�XCCf�"�%�g@���[��aa���$�	R�)g����d�r�?�s'���{

������nT
������x���+����{"��	�K����q��w�O!e�K�b��46GL4܋��x���p��xz�x��� ��N-��$�F�Ei�WhHC.h ]8B�*C�&^�DW�_@aj�~���@<]�8~�����9e�n`C��'Z{�U�z���֟��:�non"T���,��	6��W�h���K��8müoAI�8�"�,���|ܾH��#2ܨK�Ï=q��$��K���T�K6�<���u�,x��W��q.-uV&�|K���p��Z��Z1|M�=���(4 s�o-� �[��Q������qLZ��%���Ǒ�T�8u���k���ߜ�`��t�A 8B$����qY�׻��cW��^z����̔Yek��i��)y5�����''Q���:"8�ʏʫ��r��ߛP� c�;f�lL�Nj�ޝ!�gz���=���s�ڸsd�@1g�T�B�G��9a �.�N���<��.�S��OO���m��OUc�*{���R�d) }���m@���:��mk�_n�P��A�	���^@˹^�*]�Ӝ�y �R������d*	�
��0�Lbb� ��s]��(��)��ҩ�&��U_���Ĺ�j�I��zu,�\�%�#�XNBFk2�sc��9KBh���B�J�\��x\qR4�u�J4b�a~?z��4���X��\G�N
ޞ�Uj�����"�І�jo,�r��*H��QZx0n�߮�#�-"�C0�5�76�<x�f|�6�]���!Һ�®j�
D��䴗�fm}��̟�>]����''M�jp�w=oP�6o<�\w�0>�?9�.��^k�,A[#��e#1�Ŵ�{��) �<w.�O����|�ߐ>!7���rc�$�d��W8���Is�x�����)"���c~-e��T2�.���3��P޵إ������)ٟ��|�����v�ʉ��z�s{Gd��Nq�]ߢ��.Ͷx��xZ�"�x�)���DU��H��7w�/�Œ�?�'�� ��i{�}2���3��n�N�Wi��(�������ܔ*���M(���$Js��c~����H����EW�ŀ:���R�Q�pl�?M '��P��л+/��TWm��~�������>x�<ڕ+][d��݄�Q��YpX�+��p�d.����q5�}��)��}|�7�l��a������uQD�R�h�s�Ֆ.	JU����H��&����I%���$�NBI�����#*�s}l(���v�_E� �#%�jsH^�(5���l2�iY����\Zxn�����+_m��|���6�����@���^\߳���OWW� ��N�b����z�F�>�R�R��iW���#{�HB�J�i��(%	��L	�k�����γID�	-We��[Id�N pn���#��	=�E9wK8�r�Po�[��`�G�c ߉�ô�(�{
�lt:M"���C5���#�=̳u�����t�ǯI&�?�	/��D ���1Ӎ��F�oB,�}�`O��o�<���3Wc����X�~�ћ�|�p�Տ����%��=���W�Ӡ� ӝ9dg��N�n���U����H8%wKs�Yp�k�Q�N�6�H�4�*F�d�FR�:�7 b�˻̇,/X�z�bk�?B r���^�_C���
���� -��`׫��@S�>~��͋�C���Rl����=@�[��Yۅ�'�������z���3��q�)�Q���x%�ˑ��� 1�pJ�)wu��L�e�	�QU��gg^�q�I�B����͘��g��&r���.X��R(����3���R ��) �A�N~�~SՔ�p�2X��^�}�B�s�BK�r�\���A��H��Q)��#�$z��N� ��k�0�4�W��pk���iP�eLB�V`�6�M.�r�����y;$IF��7g���v�tl�6Ǯ���֬�؜�����	̆ ��,V��+���<W���1&�4�yr=@�3����q�~�T^1�fF��"�S?�8�ԍdC���ȿ��7Q/8gB��Z1H� )��\/G���1�Ro��0�Ol1E3�O��$:���6lΕ�aJ�)����P�	.�V���tft6&HZk�He)�?�q$���JE˚7�<�c�
��N��U9�Cq�|�ݔ��0�Q�X�r�~S)V�o�w9*
�X�T��V>��N��-�0e,lP��~�D���G��dQT�<<���}E�� 4��dX���x��3���d��5���(K~��1�QDV�v"S3d2� �>D���E�;X�%ڌ�?<�Vă?�E��6��')�7g�������j���o�����H$n.�b+)��i���4�`v��3�����}��"6x��h������e��6�hA����{W�����(F��Zsq�7z@�ꬫ&y,����(G�>t�^�_��T���j����=�&�[�����6�"�D��&�����o�����b2�7Ƴ�I�塘���BO��*�w=���A�Y�-H��0�O>�G�M��(��G>�9����^��C���H�p:���W���G���(Nt��ލ���[��R+c�
R��7���2�;^b4��#�ƽqx�u+`��YN�3�4�`<��;6EҔ:���Ī���6�j|�x�;%���\?��e�a�ЀD��Z��.�d36�,����$�_$pM�0�~�� �����2!�b��1 (3���%Hn��w�s(��g���~J�G�֫9��\3Us5q���@����H���qZ�Ý����Z��?_�8!%y���$b�;�w�1t��1�䈵�}�hg|��ḓ������A\��φ�'�ۣ�\b�z�N��kRA�f@씟�'�� Ԑb��d݀��O;��~$=9C<p��n����j���]�}h���R���d����3 ��A��b��z�	/�#t~\G;c�ٍ�Wp�5'"�4�::���tWx��a��RkrD��$�\�iړ�	��Pu�r���ԴAu�TP�Bf��w��HV�n�4��P�]{m�b��W�^C85����ܔe}��n�#�|`�����hܝ��0��W��[~����;���"˞���v���u+g� ��-�>=-o��ݥ�n|6��U�q�]������Bǭ�.��ˆ8�zJ֦yE�ae�8R��J�͎'z�`���0dz530eG�!�%FM����Ƣ��/RP�b� u5��[�2;Q�0er���$��|܏����H�c�&o�A�u��`nuX4�d�-;l.W��6h�Z�cͮ6BQ	~�'�Z4��躾?�yyb��И��GGEִb3]��+ϰ�ҍ=�SK�u�)FC�(��S��g�V~�#n.��S����kd	R6\�������iO���N.D�4PBE��i��� ."���@��^C#�r�⇤>���#�.�r�zN�v%�����o�y��� 
2�	�ЙQ�5ǵkD:si�v�[oI�*�!�����=4�i��`���9�+ڂ	��{�nP$Ty�3�r�<�<�+AS8Y�`]�F�cx� �<b`D�M+"'��D�H����v@/l����x3�lH���Zq(;��J��x��/e�id0��ɂ>�N��}s�Op�Fs]84A�r�ߪ>p����������d8��j�Vɮ��D�x���2oUs��K�|��I�U�����3��~�f?���%�����x���&�'�;>T���~��}cе�a�r�@j#�X����(3A��9a���9�
��z{���AvBB���e- ʪ�ۚ���U��.�eب�5)b���C�M����uQΡ�X�t8������������5�l���naҔx*�J�: ��[PjH3�U�9܉�bi�3�;l�C� �9	r�F^�$� H�d�s�?������?�������۹�$CX[���P���iu1�
?^2-���(�`��]���M;tL
�:Cő@�%��:)�.����$���ރ���t�ݷ񯣐6�D?5��|d�d�v9%�<a� �ms��c�t�g���i�:��&,�55��u��$?)5�0����F�?
��"�n̾�YȎ�T&�M��g_���K.u�v�Cesث�Rn���lj$n�q�%NU�؀�����{i��~r���Ag��
��/�^T����;�c��zKf���R�upe�2ܞQ�N�������}��M�v�N�������:O���~��A�,E�s��H=E�LȂ��4��`����c�a�s�;�+
1�>Wl�;X������,��%Z:�J�)4Оо��sŁPYNu�HKd�)�r���'f7�%1��Nȷ��",P�Jm���F��v8��K�+��R�6�f/K`��f|����Wk�.�F���y^����� ���f���n��#w��"D$��$8ԓ����
�K��v�t3U�>��8���4)M�Jfi*�ߌ����+!����ZI�?��Y���`n2J��On�ם��4Y�����[7����q��Yՠ$���}`,���ь��*$p�`0������f���{Q�R�'U@uW�q�s�Y��!��o.���+���~*1�w�ߧ���,������RW��c�#�(4���^��Pis�|U��"����*�]��Ӥꦨ�.�޲����
Qb֘��P����_$�%��}�A�35+��)�q�tZ���'`?̃t��r���5��.�煪2@UҮ��Q�()�&�lU9�J'a�-��z���lad�I���g/��X�T>a�6H��޸ q����VN��2߃�Fu���ո,I�}~���;VDL1<u�1̒`8���9s\�2�
���rƙ|����Qz���7-\�M8~0L�tA���x��T�Qu*�|ϻ�\O*AH���j]Q�f�mLp�0y�+���3����[�f�o�Ӷ�fo�6`S�	&'���ų�����@~8\Ж����찇�|w��}����<(8�(m,ޡ�������Y���H�������b��RGq���U�C�9�!=	�2v>���.�k��gTk�~C��W���,GԬ������i�u��]Ыr������D��v��z�f��`���7����GD�]��NH�1�nc�%b̶N�2��c����N]�$�����	�J��e	���!����ݏ��Q!:-a,k�3
�b-j��A|���z�byr���x����[�[������ �ʁ��L8?5h�AJ*In�����n�G]q����Kz�u��'Ĩ�L�f�y���1c�d�J&��z��j��!�p��@�����I��δ[��MT�W'�`(t�Re���4���9�F�v��z�'G@K������`e	�ܚ.�#�ޔRD�5Ќ�X$u.����h��0�&w:����Xݍ͡�~�*bc���*k}�\���g!��M)�`�;�����`�$_���+|�+���N.
��C�A���`�Cq�Ts��z ��_�1lE�$�e��`5���;a�U�}�my����ͮ���r�PF�Z��y��g��N�r�+yoѰ��=����f��^޺��*r�X"n��`�BBt$��Y@_?����÷#@��.���tҘ��׆�k�yQ
�$=��{��-$zm�ѓ����~Ѹ �!dM�X�����g+���>����)��K!��6!#�$˶|G�� ��'�z�uB������v�)��҆��~z�3977 �"��dD��� �bJ�s�2��8ț�a�Dŏ�Z�r����Q6޳j��$U&.��D�W�/���s8��� � ئ�c�co�����V}��\����$���y	��|�0�'��'��3�uKS	ƺ�㕨^^�B,��~}!K��bg�c�����;�Ę���Pf�<F�,b�1���;,��fA�������z;R�p�e)@R+\,J'��;�pv�fI�q6��s�"Ң3�W�Z�)Ğ�ES�o@z����}�YQX�6U@�����ȅ����G��(g�5߆s���R�y�P�h��ik���W����H!��Y���UJr���'�& H�a��&���e*X�&rJ�x{��0�Yd�EIޢgD�� �,?+@h�|V9I�����1;�$� 40�k%z��L~ Ľ`�7f9��<�S�q����>"��ς�N�i]�(Vb G���:�}�[�牆��Ҝ��T�k�6�����Ce�1/��	���拲gG�����&ظHK���ptDj�?UH+n1��/�@�G^O��q��%-΀�3ٽ�nʇ��Y��(�A�/%��q�������;pjG����%n�D~ئ�yG��'����ZYէ=Z�D������"�5��u�ASy����Η�^~6�|���r�!_!�:��h�@Uθ
���<���E�'؈ ���SK=���z,����@ޡW�<�h�HaS�F}�k�]ou A�OY��'�E�'/���F�`�<� +'\������T6��������a���־���b����>}�[����R�@�^��Z�*F���F޸#���uiZ�LK:o�Ľu+���(َ��g+�=%c��� �X��Q�ǀ��=j�X�J�o�4>
<`�	9�e�����Tf园J��B�Y}�-�;@�
޹��:>�i"��-q�G����q�i�0f��o����i1��yR[Rw@�џ�ց~���ALn�O���Э	ew�K��|n'��1~> 8�r�#��XԹ������:po1�n��s�#jh_y��N�:�+�O��+�nJ�����}x�Ja�#s�r;ms��GZ'H��g�����K܋i��0C?�u�ٝ{-����̛�OT�����^+Ǽߑ��O�z��0jb@t	�~�
[કL�ŪY֦b@�ɘ��x����_Z@�� ��z��6*�����z	:��7��%��~�Ό�lc��Bb�I�6�K
#�~_HT����.�m���Q8����"�/(G|-����$�FF�F�Io�v�Kիiu�Q�z���my���KK�@>�3� �puj����B�Y��b���1eb�\�Ƶ����R;z��sw4�R�Y�ܣ��Ş��2,�nn���3͝ⵖ���!�7���6DW۱�z��ݡ�
KG"զ)������s�^@M@%�֜U1Hd�4�T~PI@V�n��'�;(]g�s�I�xx����,Q�﬌t����3��p�H4�;ww���Eå��K�`��jw�/�ƘA��J��ݿ �k�`̙����8n�l���Z`��9��K��\ޅq��p}g�b�mK��K�s('��8#{�m|����y	A ���V��[/<`��i�i@��́���7_d��t�K;7�J����`�f}���N�U�)��Nx�]��u��N��z�:����_׹B=�0��ȬŒO�"Et�]� #�� �154�dg�&$�L��)�c�1�H"P��i��I��:�YN��	����A�ֽn��h�H��r��u��,~p|�ck��x����n$_���jD-���u���x�3I�6�Z��
��^��BҖ�)&�V�4i�͂`�׫Y�8>)*�ݑ̘���r���_���C*Ibo�-��k�zO�]Kq��;�+n2�;ԫ�pJ����ѱ2Ud`�g�J ��y�p=JSPWn�&�%L���%R��"���1\0/|��a	�>��2�9�%bA^�p����iE��T��3��٫YW���%zz�ʍ���)���+huǃs�dd�u�6H*��h��}�ә����ZJ�{��|Y}j1Z�v��$C���hb|������.�t�^94��������aV�6oUIώ-����U���zs؞?>lq�hխ}|Ґ9h��	���
�;M��n���7�A��nj�o��ig�����=��b9:���	��M�pa�oߝ~��>�H�B�������R�/���D�s�[����#۔[K��xCTV���T�̕���]�Ԗ�&i��4����O]�A�KM���W,k�-�"^��a�Sq����mC�B�,��^�s��n��$�3��g��$��	` 
@�p v�!�)�`&G��j��&��-�"�_���mP�.*��Y~��O	[�;�ZqK�6X�M�$ǰ�:\$)�s�������!bѓ��1�HD�6�&tج��l0���*��4��8]U����K�~�t#f�Ҏ���ϛa:X_��w�3ϺI5��}9Ɛ��5T�@�9��]������O(�]��<n�pk&K{t}�S���bd't�dF�Im{�,��}�~��լ�yY�U�.��|���`�_�^ ���8�G���X>.'�k�f�u�h���m+��}����Z
���;� �5��i�=��ٰ����[ڭ��4#�i�#t�ff�Px�&�����O�#������!�*�<���i�?/~)l=G��E8��bd��#��T7@[����XL:2�=c�-��SxE+}˻D"�\�a�dr#��@b�Μ��� d9Y�)E�Z͢R����p�C��2E2~[��o瑼�v~�f��Y�D`@26��#��'񾺰�%'W����p��!
J��?A�e_��̕qw8;Q����u�O{�7�	K|������^�+���n�Z�t�沅�vi�O $!�Qw���̂�#Gu���'§�3����G%:@�`�Xm�[1��l�1�cM�^θ�e/�G���>�tKl[��x!'����2�gD�+�5��s�/�+��,�;]t*v��91�{閦1����8��
�6}W�I�<Nؑ>6�]���j��4�A� �����j��~����ʹ�I~�G�Q�T�h=(�T��Pę��`Z�Ւ�c��P(-��T��(">$�sZ��/�o�O�ߎ�x�M�3Sx��k���Z|�kq��z���_�O��F�j��
�Ļ���K�����X��=å+L)l#.�Yb��4����2 ����7�m�dm;�������t'2+i��t���{�v�X��!�Ƣ6�i��Faa�ݒ�׾Yw!�^Sv�.��,�T�yzF��3���-�9 X5߽΅_6�
)-׸�i(\����$�zUM�&��ܑ+xu~�/��pǃkpS@^SX��3d?-�G���j���;ٝ�@x��2JN�KXQc缨��t]M���x-Fa�pq�7��[���
��R����rP0�N�қ�.�Юh`u&���(	M-"�_3���Y� b�[�.��ќ��{\���NӾ�R޿}%��t��Rw�D�Y奎���3a� ġՓjgl�O3EI�'q8��$�� ���3ٝ~(ڣ`��Q(I�H*��z�F��͊q*f�u�t�K����<C��B��u�?B�20�o?y����,U��>�~g��l2R���<�z𢖣_#S#��
w͏ǀ�dE�n����V�:G��`s�E��󆍆�z�t�\���-ϙ�>�)�w�wY��dՔ�������Q�J��/Dj�ܤ������j���U��Y���t/��3�J|t��Vi�RG_>Ù��7�m����:��Ԉ���A���S�(IܔJO�.?���F�u�_gw��:��a�'>Ui�  "O��u�1�?�~�`5�:����f�:3C�Q=�żh�7�1Z�ם�bKD��nW7~���� ��?�I;1�#Ͳ?ܢ�SuuR�G4�5��J �βrkd]'@���/�,,Xa�G��i�����Dd�?�a��8G�RZH7�x� q7W�{�FW�VtMY�Z�����[?�D\��~��t��s@�o9���Hsl��Z��FQ���(̽<̅�Z}��4V+	��/$@E�o~���R� `{�׼��?��RC*�g�^�d�z�� p���PF�5�15��HxH�ߡQ:����D����9wU������sGkk�Kc��7�5�|����ch_�����+�8��-���Z�k罈���̛�ם��XI^r`���ĦEY����З����d퍤B9`5��/����/�a/��m5�Ԙ�RH�����1Y�[1M#&�P�h*:��Rb:��o�\>D�D��d�g�����7�������X
��&ShKe�p�F��m�Si $�������T�����ص����?���T=�%>�N|��*��z�02����N�%g�'��%��E�2���}'���_�Y�,�,���@��X�F�ӝ����t����٬�L���gD��J���4Hȳ?}+j>0v���7��RDܔ���Q��}z�������gծ��ڽ�m�����$�	C۰�������t��2r���)��Ş�W�[$��W�QF�p�7�A70�w,}Þ���J8}�~f�y��Ό��������+��R�(K��Cd�f=�JG�4X{�rH�(�����e�)7FTl����D����[�7e�0 ʺ-�«7�0Eb9�.��gl����D�2Y�� ��@N�41��^�c?�����^ސ�%o�[s_��[�	h����8���}�:+G�r[Gl�0������*��>��|�����ɻ�7f�S�9�F���UJ�R]��X�7;>�`_�%#P
GPVǯ�*-��}��U��*�g�MV��j��g?����f�}.�2-�����b�>�-��A)���+���}ﶸ�����{���N7�8#~�ͱã��5Rjw"��<�"�>�5e'���O󝧉��b�ū�ruA,<)������:��ߛ�x�����MEzZe��\�g������)HǢ����j�0�����K�r�UU0���W#�� "��� ��)��a]��C�͵�AR䭗iMY�~��rV�����C �!�N����1��M�Ɠ5C�qQG}h��4?�m��l�¨�|W����7�%��uj��l�mz��9�c�}v�����|��
�o���C}�8����jl�Ԑ��D8W�I-���D}�g��(�SwW�45\�k�h�����u����bBW��Tpo���5�+"�ǀh�^c�7O��uDZRJ�>�����n�Ԝ���a�D^�0)u��Ӟ�q)(=�r)�h$F0B,gi~�Nr�A��K8�&�t2��;��G� ����y��l�1���Q�����>j^ވ"?4?`��LkX�s�e��!#�<;>a�)K�?#����w�90�O��5Py�Z��Vu�YI�k��mDyl�r*�R{b�&�%���؁*�����
C=Ū�[j��N���6Eh�s�����le�����W2�ek��=������YX):4�m�y���C"�p���~i�V�c�^��4
���*�~D��:�?-�S�Y�I���џ�:`�[/qpr.��mg^8CC�-��D��< ��[��r��C��g��~)�T�"u��I���$Q�����0[w��n5i	��I�, 8;�-�*R`��}_�Chs�BS�~KH��To�¼H��df��ou�������&���B0j
_/ ��>�;����4�²ʹ�L>+�@
��e_�u�ER��p�)���Q��x��́I��*Y�;������]���5 
�z. �6�de�Y�/��>����p�D��H��>�`���a��`p�r׷���p��b6�A�z!��-I�BVt�$_�1}��b��4�i=CY'p�!.b�P�/;?4s�$�ԗ��x�4F_E�qܝ�	7j��2��� ��C	=��򞄺��h�m���v1�߇�.�l��LVb������
�Gx/���!�<�{��2���+˸A�����Q�`$��
Tu��u̩>P�qY�O�����ǀ��V���`��G����YƯR��H��2s��~��A�%��dk�-��T��0 b��=��yC������G��L*6�u�Z�}Xշ�'��O��k�Z��5�ڋb�5D����kg�D��%�I���ȯF�������a��������l��+T�O���Iv\F�'�q�����7WX�� �p���~V�x}_v%7���ܻM�s����1)���Ό�(\�f�Fg��VL�ī�g����з��2APR�8�|߁WMو�d�� �GtV!b�0�݊��ZA[td���A�����gޘA�t�]�R��Wa�-<zW�E,������򋫊6�c;�%�'��)�Obf���D�ҧe0[-���f�`i1Ǻ�6�_��p���	���]���eG5x����4�o�i�A�Him���ʜ/d0Cp�?
Y���/3�����$Ӛ�{]��,�5�vqUbjfħ>�e����� +z84%Wf�&�j|�ao­^+���,��E*��;t �������Y/MX[�>U �S��2}�KU��mQ&���U*�fTzZ7��B�Iah)��§�0���C����^#:��r��v�X�Esu�(�x�s}��{�>�X��V�s?o��lC�eu����2s�_�m3�[�`�#7���Ȁ�Xz���ݳ�M���55�|p�}���ق�7�^Q@Q��t��U �o��Dk
����	VG����m�҃A�\d�}M�{n���s�d����o�C�9�0_ռ�@��'��C�.��m�Pc�\B��;(�N�[�M��G��S.]k	������Mc�ր��6�������xP�O4yzJ�����P�i�3M�G�qZ�B[�Rq�Ƥ̕�$�4���:IǦ;r�=�����r��fw�k����>��+�����E���:��wMd�͑��
f*�j*{g�������7כ���	��Z�W��ɤ��ԀF�U��\�z5�!(%�@~��t���T�r����eq���tWN��9�	Uab@w��/��Mf�8�y ��Y�" W�R�*	Ȼz/�ȑ��/j?vl�e��2�?,�j�5�i��8ܡ�R=_2��[�M)XbL{�h��Kn��v�y5�c����4/eҝ0����M�ջ|����`��:��'ٶ�4��s+O=�S[B�/��:S[��	�
\����@��R��K[�^BE�h�>�����(�W3hwZ��*D�t�*�UΙm���>������T��r5���i��*'���������8��8�d�����z��<��|J�^̋��-^��Iw{X*�\�d�6���l�սNt�-xJt�&c�0��U���h��C�5��v��L ������i!�/̵�(
�}z7,9���yA��2��6U�	/���X����D�\j���y�vS89X�V�z�Cf�،�3��xC�#i�&|��f����&v^�����ˇ�/3�z��܅֭�Ķ��"��η'8�q�M�$+�-�����0y3��b��,�� ����d��o�A.�Wo7�hg��!�`_D�v����S #�u,!���s�Cy���OgH�H��$3����0jU�JF3�c��y)�d����:l;�O��9�Ƌ�%(5�ӑ?�(�ac����-�c�R�g�7	I�N
1noj��}��0S<'�O̤5V������ʕ�w�w� 6�����w�]ksq�ك�tgF%�dw��D�}�s���ǃ�t�}R T����p����b�ΖEj�uݒi�l<��C�n�?�)M�J8a4��W
Bz�O�H..�����|�g��s�P�Y���鐾��No଱M�1����^b�����]��}p��5cr�ti�7���qF��E��c�\�}Ӓ�ʹ����'b�m%�%_�����1��
 ���3���ݤT�T$����ݼ���	�6��6�Q����6pt��;~�n��xԩ���-h�����-�u��.��*��B�t�kG�H�#p������E!�yPN
�},�6�&��3��c�������z�� ���v���U���thtm|y�if\�K�c��\�8+T��k�W�UƦw�5�1q{I!M��*.�$G����ܔGߓ�b�WOW��"�-YG��1�� L�DS��U��)��ao0���޼Z�gbQC�k 7����}�&��saπyr"�=!��ǉS��:���4�ZXV�*5�[m���E��K�x������б����ɤ�'���kL�C�$��:$y��!� ��֭���}�Ws�s��4��i��KE�w4�gv U_�[RO(�@��uH��n�a�#r�y�����2�8�W�U)�.�P�Pΐ�aޝA��m�X�B-uD���\˫�(�����d�( �WV�F;� ��(玓�f�nf�+&�1+ŝsI:�Q�I%P�P��F��sԻ�.Z��u,x2�٢V����|2zB��������[�d`�i[0>���9x�Of��^����1��Dђ�(߹aB�~
��%� �F�z��٢r	�y�ċ��@sIK��/}a��8�$��O��7��_�J\CߓK���W�S{C��r�3bif�/r�oE��"��@��S�J#Bb���`�܃�~�H�Q�R������������Z�h�Q�לJ;�6vA/�J~掝�v��VS4�U�W#�$��	���>��_K����j��D��t;U�����a�p֊X�)���7� ��w���~���Y�����Zbs�O2��9�6�@���FJ��͂��F��`��M`)V�qO_�L²�-C}�:�FЭy�
E�zr�}�1��L�ӿhJ�5����_� ��~�ˆ{`Ԫ����hB���f����_����pۖ��,7$��s��4\"#֤�M�4���Vl�<�yE�{t�ݔ�BS�u�k�'rH�- �r|)Q����kѓ�O ��Ʀ���z�����lʿe=�YF�|`ad�T�}�3��yI�ό��m��K�^�3%mt6�0�f���3c�}�]B�/�i����Pp'{�,������D����,hu��=++��j�+
�q��Ԡ�L]���_������[��Z�z�2r��"�!�&7	���c���&�L���	ĄD��>���zF�0�i'!x��k��AS�+���S;��3�+14��YZ�/A���R�P4�M�C�#��b=M��RU���E��R/Tg9"���j��e�<`����I:~]`�s�H���B����[���K������1?/���5J.�)��9|�b�EVwr��1�y�8@˰5ǬA:��P,��F�c�Z�cpZf�r�-)1a ÂA%�%B��+3��`W�z �����	nd �c^O���5�8n�f�K�*Ҵ�,��.#�0�2)

�u{�O��\ɧ ��%��(�p)�'���g�`�ɹ��_��Z���/B�a4���$s��F̄D�q��z����X!_��X����k�q��bLw��?��� ���).(�; ��3�Z����K�+�B ;��N���[��K}�/Hˉ5z�K�Õ�ڗ�9�:�tQ��.�~Ґ@�~���*uJU`g��`3ޫ�z B�G��|ĺ%G��R�^?:�HP-�TQ�y+�f{Ѥ�;|£�Z�j�`��M/���R��h2Vp�Q3ھ�O�,yq����Ԛ��%�ڳ�1V�%[��ʓ���3a1��Z5L�E�7Z��em4
�����H�T�Gb(�����~]+_���5��8ƉT���Φ/�ݴ&C�v���xo�ϣ�X=1Wq֩��^�����F��x9�^��y	���:���	�����7��|��&��5��E�$VW���t�jۢ�>���r���ܲ}�o�Mb�P�
�%��0W4)8<x3�sd�y_^����eؤrg��$����3!����Y�d�t*
�ˢ�C	�}���O�6x�}�^XG��[i�Fعϱ}�k�,f��%#��L�
�)D��C��Z�[w@`��Ry�L[>G�htҾ7]#�N��B���9�C^��`Xi�	0����)�q�L>Lcf�	��M�*$W;[�^����>�hE{�6\O��6Ж���.�Rs�Jɂ/;�$�����Z|�Kh�Q�u����)�}������ұ<����	w��Ɋ>���"�*L���x�5!
q.ݮr����(+�G�����j��5kh�������Sz-`n���ޓ���@Xխ��d��a�^0�>
��Q��8�yP�nYv�T�2�P��8�T	(�I�сz�A�V۔#]��|��8��wn=2'Qc�;���q���$C��ͺQ�[�����
�.r�X
�	V���#Ly�u�c0Š� n�jafN䝧6�3OE��WF[���V`��Y��v�6�0��qjCe]-<;=��	k#�OTr0Q�p���OVt�d�'4�j�{�x��3��"O(ٯV�=��m��B_ �,�����������W�wGh�}P��ۯ����u��⎏�@�=�U�V;�����d���s��OĮ���X29V��џ0�O��u�58�hx��{(S���aa=&t�g�)>	���0o�xs�U�p�;�,'��Ϥ��=ݭۓ9��P8Kݚ[�'�s`� �s;\�*�QU���͟���p=��Q���19�G��u&�ˀP	`�1QtOq���׉{��F��v�9qqKXs��X ����Ss<?	+�)�i��n,d��!���H��4� �z"毻�*�I��S��[ �G���B!Nw��"/��η���8�jyo���
�K����Qq�ìNuwv���X���j9��RH�����\���*֖��d�����9{�����E��ϵ�H�ߊQ�m��t���d$W"��k��r��A�K�	��	3�+Mk���42gjG�Y� r�w$'�6�+��:|O���"��it�9xf���_��x�vbU�#u̉CSi��=�%��F_[}bOw����|�x�o�']�AQtÛ�|C�y@���D&�����6��b����K�Gh8�"	7T��nw����A���{M�/�P�Oi#�V����qC�Re���/��3U:���]�zzC{BO��7O�6���5���=K����ȵ������L;�+\ Aj���{J���e�7ٮP��;$�S>7�㉿鐕Ŷ1%Ƿtu��]�M��=���w�
�H�WD�c�_%1y�s�.`���L<͆���#z���}ь�vkT�N:V�A����t�:���My�6>sZ�ؑ�~�h��o��ae������r��"d�>Ǭ9������=<��0տIq)��Kk�����O�
�~\b�+`�W�/x�q��Y�A;�s����i�C<�w��LVh#{�����0�0��ڀ'j27�p�8,ӯ�������T|_m���I��X�v�������RD�}	��ASl���� ���~n'm�v!��Q�Q��Sٟ؅ⷌ=u�^�	�@���+$�7{�3g�)�$������K)ͩ�%����E�dE��+�$�2w>����"�C!J����?��������E�O�璠����楤kƇ��a��L9qL��p;���C8e���jc�Cwn���������i��F]Ȏ���<%ʣV:��%D�ٙG ���4|�ǊɌ���%��o�j�3 G?B4޾n&�h�ݿ�r$\��,�-ے#��%���7L2r�(���.������gHz׊���5WGm{��a���s��@G��!ݖ�B�U=�8).1ZBV�6�����u�܍7B�s����6$�fDX3K'v&�Q$v؝n�A�r� ��l�Aۉћ�e��C�$@���A��g6����*6�S3���MǨ�«�%{��ɷ�Rǖ��z�ƥ�h�c����#s2���6��7�����f^i�4��H�T,$����&Ю�'�I-����D��="��
$��5��j�eb>:�x,�L�r�̅s&W[,�x�,�-�i
^����3D+�>8@f=0��3�^\n'b�g�1�,��7��5%g�ovQ*`����+��2P��o�Q� wɃ���w���:7�@��Ķ��\������=�ԄZ��
e
ڙb�ºR�r��N�-I��+*:�R���o�F��4%X�+�R�����sY�U���!���F �w��I�ՙ����I�+�{���}� �<�A�O_W`� ��	� ��5Ml|n�����?��2T/:3u����v�#�F���YvU���ܬ��6Y�hp����¥��`�U��n���z�����_8�Hb�,��a�f!�=xo����!��vl*����fW�7=��>�ܖA�w[�>���C��8~�ï���[�J�{atY`G�mK�K�t琿��(C��eo�vF[��������M?hd$~+�����<rcv�V�IQ��u6�������qa���射%ikq�Γ���#�;��7�z�M s��ތo@=���w��ks��텐<�#��LAʱHl�	�tPq���,��N;����΂�k�O<3��M�ʥ}@�]�-�
��7Y���^��a!x'�˷�!����ybO�����?��.�?]ʀ�B��~�����m��u8B!���_��o�y㿥Z���u#�'8F�o�
ݨ��r�k���t�P�˄�b͂�6�(�q+5�M�RU�(H�'Q�� }0�w�0^ډ�dע�¬
���Bãs�Z�ʲu�q�Z9a��|�^�z��u�&��lI��}��
V�]lŕr3��<m���;)���= U��x�c�RAE�:r�NP.��<R��&L͠���8��{c�I��P5�4��+��f�=D�6�"��l;\��V�Q��TU)Z��V��m�7�[��c	g�00�����:Q�J/<L4���/�$V��ئmTuT��LXº�2SZ��R��9�1�E>��%29�q��C�����\YB�.yK+8_�Hs�Z������:��`a�/��(J��s�Rj ��b�R�d=^��M�J��0{� �?�ʾHTخ�ꨓ�T��K���7�]���rz��`:�$r �}���J0+�{���EzB]ht����~x&±�>�uQ|�:�V��g�KS�ܼ�Y����M)��k�����x�Zo���Oj���u^[��G�u�ߜ+��E�2exzP�D�tt�sv�"<DMz5�����d,)o%���}�������y��4}�Dg
�FE��µrR�&��0���=9�kv�đ�?Q��hoO�6�d�4`Ɍ%���'P�<bԓ	�ـ��1D���PhBۙ��r�����E�\�*����^:.X�l�*�MY+��R����t��`!� ���g�
��=�<N:$1�z�'Sp��{�*&D��x�x��G.֛�ez�6�1��]h�Y�dU&5�ň���M	�nv/�cv�)��R2���]ƘL/��^=����i��}�8�g�|�mr�N��|��n�^�ZA�,��d��&'�u3�$M��I�O�q���sL4�GA}�Vu�Z�Jpl6B��<;��?�\sȔ�+s/���i�����( 7r��R��;Xg��R�t�|,� a�<}���C7��2��k()-?�C����c��7��B��-�W�m9���6�H(o�Rꕛ��(1ߕ��5�FYe��s���[�瞝��3G��*��r����+C����;���2KD��Q�.ҍs?t�B��\���s���}���G��_��g^k-��+y|�mv��z��d0�������U:�*	T�G'��IY`K�u�#�7��aM��)��z<��,.�^�f��BF�� :y�U��YwɢL�'mB_U�1��*�tϨ�
]�`�iD�c�8fC7�̑�~�髝�dK��`Ēl�W~���5�\�
7����$U�*׺x����	Y59�>U�,^��w��{�zn���	���@���~4W�n�(�2-�����2��˱x����l2"�2�J�m�	�T>M�b6��k�����(%[��2P-G�cl}��h/�ŉg5Nʮ;�hJT#��ޟe�t!�ʍ��^L�r9�6�ww_J��R�/=�H�	�TA��BK���*��$GXN���^��i��y󑑚�
F�D�M�+��|�����lRi��L�W$"�����
'̘�h�I��p�;�`1����}�F����2�����k���Г�����e/E]�r��7fz�XυR
~�/`	���5����S��G��6hU=0K�f�M�ݩ��h�y��<�O���dJ~���:�����%T$	�3D��Q��g��<P���u^�LQ��8���j�ri(���~
i�txǐ�"G$4��Q>���n�Du����s���t;�d"� v�%����2����gg����mj" ˑ Y-ֹl��!U�r�Z�p-撹x5Pa9��(}�C��B�a�W��������D++��wD�:��A](�_P���z��?o�~�T�=���n1�k/-'���B5���}�V
D�h���-�k#���6P"*l�IKo��{������Y�<��gs��o���jC�&R,�O���jy����ܤI��1=��O���g���ޚ���i����ɑ����x`�u�o�+.9���sth�DY����pT�n���ýk�l���'_C&(lā+��&��M\A���/V��	�f����ԯpnt E߹�(����ցP��H��і�&S�����0��a+�*����B�f�	�bZ��!s�Z؍\�*�KT�P�w-�Ώ��3(2ظ!��g���R�q��u��X�n@f��2�0��<p� G�-�t�`�V��.�R������+9�TYRY�o�w�J����fi%�D���n�gH[6�u�c�^Bl�oό���fF}S�rp�%���Jz�LIDq�2ه��~'�p �=��10�����tCG���9>.EE=�b���yy��}w�����@s�a�(��h;s�q����4d-CI�ai�u&�[�U��@h}
�)��r�h
��?Bw���m��R�D��3Q*��vw��$'���P�O�3�5���1w �"�l?��&H%nAu�\q�_����(������B�,X��"�c�?�n�ū����͗�(����[|�z��,�_���#�6cPfED�3s�J�0���{���u����m�p�*b��@.M$�3�勠�"d�0�0�:�.��������@_�S.A�R�':&}�]�|�Ġ��4�2�Q�{'��m��E����5�44���JQ�;��J��>�ff�,_ǟ�O$�EN�Z���S��Z��Ko1���M��nT-��W��Z\�(�V).%g���ϯ2ߡU��Ǹ@�6��SޭA4T�y=��rN�O���#�wr��T�꟦�5[��C>�U�f���tU�z3���u;Vx����Z��r�9���Ŗ.~�d�	���_:��ω5�;�
��ϴ�Q��(�-~ mW��.���1�����z�6:�U�EK�O��T^W8[K�zh�j�7�gΎ���_>_��.�*.n5m���ⵌ-��q	��	/l�?�z�ͽMV������d���I�3Ŀ��"�h����g�����F��?l�f�#ܲ��n�n$����DR�YXJ�r���6}�7��N��z�W�_��p�Uޙ.��cZ�#��E>���$L+CK��i] �z�Pn�_PD���u5ECvp�f�l��,=܊��T�/\-$&��c���/���?I4^������;K�޸1�~ᛸ�Lit�lXqW�P���>�h�v.�WBU>�<hpɴ'F����~�$�g�g�w�a;Q(�(�[јngޫ��3��	z�M�FI.,��6)�C�󭭯Wm\��qS�a�+d��t�3>ǔ�ο�!R����'9Q�ȥW��Bq8�	˜�U6Bcw�y�F70nLQNTddq��ks��,���ƣ��GGu�_����T3c��S�E���[6J2~J ���-�a"�ڭ�k���9� ��cҫ`d�k)[gs�$/�6�j����Z�yP芇K��<�ᑍ!��J�5/n��=�4����"u'�c����r̕�K>�eQŠ��)F���y��w�@���(�^G��+�u�'�bM��.!���g�֝C��EհL���|��3m��F�N�[����_�`f�,�|�)wf1��%j��C�L�F`T���o��n:�J ��1U���&�>5�܆Y�� Zg2 �O��~���,�����n��צ�~���;W2�]<iu�cH;��U.����Q��9��rS�LΒ�[��$�tц�\U�R+Os�W�#ܜ�Ň�F�d�����RP��eh�G�5�Qo1�;�T��<R��X-�JG�p�D�����<�0�� xn�C�P��:�pɹ��K�AtC��v��édj�0�k��|Qy�" �|%����%�A���lW֦�4�D<#1���s(�l� լ��LP���ɯҔ��B�fzH��8��j	��9^���4�B`%]&��Z71\)�C��0<~eL�C�~���2��]��(g{��}1<6���@[����nXP"��j2�Z2�v;Jz�]���*s;�$�>̯�eϭ�\Y��mi��=�]���?{&E�ʪ�rOܻix�G g�G��6:@�=��S�������hH@��!׷��?�H�4��;�����!*aN�BY��՞ZuhT؆�
���N �)��U�{��G@��e_y�o�������~�O�5'�D��Q�0���2'���C�
���>��5�S�����vq�i�r_?�7�^b���2����]����5�`��ٱ�ޮ�ch����+:�F{�^̉��aU4���\��`�ꬪ]F���j���W
�K�	A|<Dd⣷%i"˷ܤV4��Br�a�w�bS:z�c%� �N\��>����j�i��S��ZE@��3@�(��`������W��
, Vy�cӾA|Jg5�N
�^��Z�ϑ2>$��wL����S��F��v��G2݉�����v8��揆$S�m��Q�-����:����-F���Ѣ�_�^���O5��L; P��ϡ ����"�Џ_	Y�*�Ò\
M��de�vf�ȩ���,���%�f��3O97���?P�)K͒���\������8d��-���p���̑�D.;�<�-��aj��^1OLQO�89\za�Lt\y��Zכq��ldn3�fh�\� �t����}&��\l)1�T�*ee�J��j�G8ž�R\<[J
ӂ�4�dRvj�C�W|#�=P��[�|܂O$Z�Jvz��l�c��^���H���&��bj�;��D�֮/]���{7�EӠx��� �����WE��?C��:Y��6tEVC�5cK��Ǘ�*�9��s��p,Ө�zNSy�����8~e�0"�BJ���r��Y����h�Z&1[S�t@� �r����p�-S�վĞ�[bE?N\?!Bd�"=�dO�S��4�hE-���� s'@:�M:���s�@��kKU����P� �
qAg^=�	��-�Z"gV�Iﯱif��%㪗�o!�L��' �D+�V�O��D��U���l����"���\����Ц @�=I蝘I'ץ��4ޅ-���5�g���gߟ��S���~2x��>l��8�ۺm:ڜ;Q���
OB"�4}ʃs���T���]�3w>c�Y���[�*�S�Ky���y
!Jq�P�������o�V+(^C�c��'<a���X��P�n����wtic�6����__��2;�&g��ίs�H���I�qT�u���6����I��|}�i"�uiR[�\�]�"#94��rc�<��ȗ�7L"��j�OH>l析�ڧ4p��'��H�� �xCplH��&�u�b����-�4�U�&��,V=�?nШ��Ƈho�}�k��em�`���M�è;_y@|#����]�eE����}��:o �.br�#(�b�p�i�:V.V:�	[�O*�ͅ��6��	�h���mڱ�}3�<7JI�<P�p��i��䯗����N�^�F6;���H6���
��V��!Ͽ��P�;��x��Td�]ͮ�R3/��Iw���4��������Y�!�xx���L�![k�4��뙍��p.}�9d�)���T���0TU�x\.�*�G��DP��BG�# Х���Y2	�P�L��F�H�7&�ح
�@�w�P�,�&�G���B5<�:阰 ��׫b��V�y�ڒ�J�(-�ى5L]��X��T�Ӊ��a�6>'��⑌�<��1Ft��2<���AK{0l�<s���GTi�4����נB�n��Ը�^�#�Ϻ�g�J��>���9d�X0��x���豐me̆��I]T�1�>HM��k�����W�,u�)_ggj	�`�o��&��v�u���-��-B�O��������X:�_��{@�lG!q'����~&����$/ w�O��Ѯ�4$���$T]��3��B��v���G��\-D���������{"G�*��ʃA�#ȖF�g"��=?�uD$����i�am^���!���]y^[ow��� ��i�ꎡC}�� K��/ԡ�� ����K=�&��ʶ�/�ݸ����]���j�X�z�qb���bb�����쀖�Fp�b�?�{��棴���}�xe��]�p����{N�B�U=�M(���Wqc��'���E(kyxݐi9��� �q�{8"�85X�]QZa��*��8fF���"���3��뱤B���A�՚�)�N)�;�Iu�P�AJ�8rOI�v��ZN�|�I�&�"e�e帉�m���#�BN����=�&AtϡW�����~���Ǯ���Őa�p2�=�g��2��p�A(ǣx���y�>=��H�n+�7~�B��-u�P�Ec��c�ՑFLs�t�av�\�@��$��Bd�+��?.����\���������@4�?�õI�y�ٓQ^B���XE�tƤɴ� y6Ƒ�����ώ��M�e�V�x��t� �E}HX��%���O���Ջ]\:f :~��02p������ĭY�&<� ��>T!l��(���3��Kj��}�Rc����ό�-�F�������G8D��	WǙ��`��	�/�1���*�+�?�/9M�����)�·��i*��.*d\�j9��3�b�RR�==��.n�b�K�Nzߑo�;k�DQYl��>Z��j�#L��w�q��kwʭ�\2EɃ�㣷�k�n�����̊������"��=���E+~�
21*1}���/@��"���V����oNt#tsO*�1������*�6����Q�	"�/�NU��0:S�qH��݌p#l�:fg8��\1����U������X���v@B�*��j�9�x.��ӝ8 �r�1O2�
fMO���B"�W���Н�m��np�$"�衏�tq�"_5�v��e���' ux�X#G�пaJ����$T����y���Z~�p�F�(��i�'g{�0&C���ೝ�I��J&�K1~��|�֧�Ȑ��$��3CW�z��!# @3�>lꔇ9.@��1�d#���@�Z���U3cl�1Yf���Q��Rbn5E펼���d�Ml7�/�L(I�Z����q�А��דLI�8	��U�qx��c7��<��qu�S��頓�!�P�89�"a7B���N�7��׀���`�ca1NH0=��\�b���c�A�g���,E�iﲎ�"����N1_�6��Z�����4��9�{u�U�q�kw�bZ���x�|�tݜ�0���U(\8��
ٻ��c)E�O6t�M@X�9M�D���1/i���,5�� C���xW�p}u�rAt+�Op�%��hM��v{R����c����Cќ��Eg�	�Ow#t�B�M��^�ݭ:�3�K��$�
O�F�py����1�g��"�l��4K����V�c�sl����QtؾfG^���0mB��IL(.���@���U	z�B���4LY�J�%;y��5��e�7u��B.�m)��Dx��#]n�0���Dm��M?��1l��F~װ&���*u�Jf�J���Ef�L��f��ƅ�l��QL��R ��9d�˿���	ny��z�K<�ɳN�؇u�'yhxU>]�N�4��jm��%��O#�/)-_O��Xc+�)3���AZX�c�h�Eg���њ����S�T����
��"��ǍF�/^�g߬Pk2�Ȑ��J3�p�Ҥ+9��'��
�^�N^��/��or��RP�\;V�Z���>S����3�4�h?����}�O��E�ؤ͚����mW��x�����pH|��zi��T9������#V���B4EZ��f�����GF+�͚�����RG��� ���K�L+����tlOE�*Gd��èJ��UEMҋ)k=��-����	�'���\+/e��Ļ�+#�.Ou��v���b����J�-��a��0�%���F�w�}x����$H!�X�(ej�-�
+��\Q|�dFcAl|��<1�v�	$��`���A�g�3�2� "�����'��Ks8�-E3^^����_Q��+��E- ��@"?Dw')����ec�����d��b�jx��6mbu�V�����U�l
�=��\�������]:IufX�f%U<_MK��J<:N|�t6B&�Y�D���V\�R�|i>��dP r��mB�����cg���>�[N�8}��k!b�7y�/��se��=t[G�v��yS��dv��<�畝���N��\ǣ�ݓSs>������D]�"�A��%Պf��X�6T���K�+ݵ9ɞ�?�D�=	U�0�:�W�rӇ&L >�`��HȾ1�6�����o19�盤k�TA��x�r�p=`�a]���5�<+�C����S�Ղ͢m�Ґ4����B�;v�:_�]Y���k�y���a���~R�۳E&?t���}�2r���QQ���X(�� ��_ɚ�0ݐ��WfU��&�t`����gD1ٵ��
'i���k{���:?�b��&,�Mh@Rt�0�r�%VlG2�M�\g�0Pɭ� �o܉ K�~�0��ӫ�c��C����C��"��Z]�K��SH�gtq��#��b�s���I�}`j+k���IE����(i�h�A��th�]����-\y9AKW+��K;����$�8c�"&��N%�Y=|�~�w��c�K���=���hj_��h���vg�z����b��K����έݬ��hh��ct�m���)�� b���L̒\������H;>z2�C1l�Td�K��ke��_��c	��r���ק)�0],�6.��۷�7�V`���oT�s�O#��6�TD����	3K�j�u���c����p��Q��i	y ��4��r"��8���2\<1�y���Uɏ�(���x<y�cr�����.I��[��\)$QI�����b�~��#�F��{���Q����>�ass|	@{�&2w��tl�LG0C�N���D;�$%O��o����HϮ.�ÛB���`_��$wj��(�<�/6����#���������B)ec�{2��1X F����Z��E�&%���`x�� �ԦY�����RX�yvIR��#
j�R�5�4lm}�՝�;�Y��Mΐ����|������+%�;��T �����y���Uq�-�W��k��|`����4�M�A)�t�����D��QֽBD�Rv�\~��$l������1�u	��ɘT��$} J��J_��e�6)N^~���{����	y�T5(�ګz5�Tz�����'�n���`�ﬁU�i�,�ޟh�;>��Q�))��f���R'�����p ��u��N\��nڢ�-EA�r�|��ҖM���O�ܮR��8���ئ��qqM�5I���h���1W��0D�?[�hP���'U騀�e�A��v�����X��cGkIz>��w@�Su+��An;����d7��
�l���ϟ'�IxK�]�R� Q�"%��ST�'F��&t��"�0nLN_o�%��:;����յQJ��ԝ6�"��LR�s�RNF��I���v���x@�jƦ�l�Q�����?�#L����5te������-QU��	�����A���|�ٖ�ȡ���� t�|5�|��;�>���5!���x$c��K�<��<UŸ�,��f
4��0ˠkaj��W�f8/~��^����&�*�_�`]{�[v�#asS�?�3M�T3;cg2�D	�F�r���A[��V7�ݐM���%J�����o���[��s�m�� Ӯ�fW��:���/;�=�����G �^��eDV�`��\z��`��(H��η�Ƞ�A���c��nGm�%RٯJ��a�Ŋ�n�l{��1;�t�����=Ԥ�%�l{S�dr��88v�r�zƷ�~R�j�ₔ���{UU3��+��k�-* U�/3,$%�k���p��崒F
>�%ת)/�=?���V*�TD �Kbd��D6�3 �*ˇ��-ִϲ�ql�E�EĆ�J��J�r��7s�����!%��*ZQ�~dH~M��9P�)�sfz+A��pɇ,�Bܬ���:�ro\��~��uW���o�?_�ZL��,$F�!�"�k^h�E�.�>�m�H�-l)F�n��l�O����+�@7��j�yvh�|	��H�x���Y1�v&7�d����Eb���B����ލ�0ؒ����5�:�8}dñ(W�J�1M�Y�\�G�����'� ��>�J�-��/J��@�յ��i���p�>��TK� ������K� ���9�2��h��&(����tIݲcQ�B��J'v������#^�:�%�~5
tڟ�Α|k%0�q$�qkW�(N� ������G�Ǐ��r�:�Rv�R�F6�D@Q��tQe�����U�����m�˵��5b�K��m�Wc��E�UUBbYl�1��2�~p���%`����T�_@0�^�ii_�*<j��z�3�H�i(��:����c'7��f`��;�����,xVn��� r�uG@�`}� �P�kg�LܰQ|��Vg[�X ���)��n�e�)s�m���ɶ��o3���@�`��3|�s�J��]]>'ŧ�$L�?�nN����Fe_=�^$�J���6�-�C=����Z�k{B��;���-�X/�Ӣ�S�weL��A�T�}�fhz#hwI��6�}W�j�m�W�c�jj�(�j�'�xףϕ#��,���I���T`�7��zl2�o03�_��J��R,}<�B7�u��Wd�A�d��ַ*^,��:��]�n��PӐˤ���{qv%!�7eD��>P��e��<�Ѻq�UZe2��.a��]j^��;c)�����!/ι���h#�������V[�d��%��L�p9"|CRcwo��I�l0TB��i2^�m6N"�<i�!_ $�D���B
�~�a��a�@��'��m`HsǬ��k�r��DG������^�5�ՈZ��k:� 
`썚�p~�\ߢd�� *�*���O5l�s%'b�s����2B�������,�N#X���V�?^(�%�s�3|�N��@��hS��E�KB�vTa�����`�|h�Pf��uO ��j܉���MY��{�INT�2w�>�Wa
]�'���K�vxZ�3��m)!��(��N̪I:C�A��I1�f9��M��S��gݐ�G�=�%�3×���С��_3y/���D�w&x�#�x�g�ۿ�/�;���M
�Tڨ%�!�[@���TɪBK.m<x!������h�(�I�`�:�oy8�I�ُ�p���J6Q�������4f��`��dQ~��iXV��|G�!L���+��F�x%i0�}+��抅9��:\�ך��܏L�t����Dx�e�mX��{<���7j�Џ�<i�:u��?�%}�[T[s�;�{&���Ҵ�<�cؒ����Q�.(৒8�� 4 u����o������i��R��28�i�Exg�[��p���� =h){c/Ee�@�������X�iv�f��N����nJm�z��y׺�Ѣ���Dal6��D�U�BJP�aL!�\�oqLcwl�F��"iF�0`��͑�|�6}*;	}�Μ:�θ�A�-E��.�Q��ԽyA�ǺݼbRd�?Q�����1/R*��U�n����i��`G�#J�Or+�:���s�f��U���I`�j������.t�y^L�,N��Kr���i���1�N$�H yʧ++KT7V`��:�P��Z
�2��A�v&[����Op��q��HO�`񟩏��m���#q��M��h�ѫ���{=��rP�����(��"R<Ы��y�Z�f�P�����J��T�d(�^�@B�`P�S�}u��u8�=�ą��m6H�M���bw��w;�G��6����Pj̚\�=i��o����M��OKw4�,'v[�Xn� Z2� q��1}�߁x-�`2��{��u��V�w�3W��
��Uh�1i D�U%�A��d���Hd�/dq1��y���c(�D
1I�0!��0���S
6d�;X%c|D�A!���l�W,I'�d������CkZ�S��kph�Ә܋�}��xY9�{Ȑ_E3R]�vN�&>fऒ9�x3w��~]TZ��d�V"��X�%ɝ�K���.x#(2�#�[�-�~z���!�&u���g�-�P���}�P6��Ѳ�䆝H�`{ w��X����ܺF*n$���T}�M���t�۲�T�
~]�!���R"�^��Q`aON}���A��B�����I��	y�I��n���`L=]Y�s���䳌��۪0�u}=�Q���TS�M#�jI
�l���,A":�Z�F>B;^u\��@�����(|��\���\e$��ɳޗ��9ߩ���>�Ǻ�<#�T��$��]냶T���h0�]~��ݞ8�� �/U_��]�v��3㬓�8���{5����a:X:��ȕN�B�{`�B":��~X����*���n_�W����@�"�|������K]�!1(h�e���O�l#xqݎ��!��Fc{W����먘\P�z�5����Մu���<^�F�����š�,>��-�����}��=G�c���ImJ{![���?�9��q9XV�IX]��UQ$�ac��e��<��UT�|�%6�ۅ�+�~B��19�]U$����@s�0%Vo��dI+s�m�č�7	 ���t��C��c�8�D؏�.�@�[B �l6>E��-QC����wộq=l�Y7H�hn���
CI,9�UF=�|d�����XN����I;$��C����U8����ȑ~�9�"%(4У��|�	m1Tt#���mIJ�;z���yŃ�,��K��O�"Lr|X�X*O-�Ќ�so5C2҄O�
1F�k��I%�Ioݏ��	�:��E�J+�v����!W��8��
��C���x�i��\��l&X��8$�RyB��9�����"	#l8�N��~�hJ���T��A}�YGF�,�F��$��B#��w���\q�;�S1��jA���RSvzM���.|Y[�/ይ|�55\ͥ<�h� &'���{�R��j�,߰�kt/�̈K�1U�Yg��H�f��/]�_E-瑞��3�т�"җ�jԂg�02|���kR�@���p���pi�j^(���#XSIg6aqS��%qq��=�/,d��Ps�Z��q����p�������Us"��ojYO�:j Mn�$�u��]i�N��g�t�+/�������t�.�]�;�0z#���x*I�zS9������D��M�WIbފ�堋��^f �b�c&����gah���� �r��5l�n:�M�ۇg8���xN�߃�zbN�9��@����Q[%�KVV�$O���C2��P��;ɐl��Q�0���~Aқ!��?�]K,���j�|]��5�#��u'�@d
�E��t����F��uw�L��
��E#d(=��Y��>W�|�o��>-�\����]`I�o�x�r,�j��5���q,�*�אd�t�qe�!0�}&��b��SD�����wS�g�$��b�����!}�
���4�jKY-�t��IY}�3a��[(����;G��[�*�E�:���O����m���җu}�.Yd5����;��7ti�*�|��7*���QVl�J��M�F�:
���x5�ͯ�8��wN��؊�x���[�?9���I��wx;τ�sc���r�5���+�R6��2��%x��E#(8��D��Ƚ)�Tv~�ʷb}���8��-��DG�ev��a[-��<*��&Z��&��V�R	���G�����Iv�gk�Y�+�mT�P	�H�Z��6�T\6�5*X�T&�U�8G�܍�t��t'0 pr�hnJ������{R�:���'��:�LFY�����5�!�_�܀�%�iTİ9�L�������H�D曆R �uY���8�5�,�Av4.�ct-e>�{��n?���4*��&e����4^ω��j���B��T��1/����M���7ʧz�vI��j������O������Kw�z�z�z����(-�4���W6އCp�3��n����jg�͛��aq��SVm��Zl�zi3���e�	}JJ�h�A�YF�@���j���c!��vS7Hoq4�Ɛ�Υ��{G���3���I\�uz��5�-��~����:��)v4��С�Q���N��' \�!��g$�����b	r��'�ګ^|4��f����^����Z�t�}�=m<K��C�A*!�p8uK�yS�L���@�$(핛w4��̐�U�g�b�H���e�h�!��Yu?�0���j�7�������F�����q�hlۡL�g�����H����YSB,� ���Ip	`�y.�ʊH ����D�$o_���w�He�R�� �j���!Ў�׉��R���_u"���3�r� ���}��y��+��KV')hIT����Α_i5�c�a�2�7�Z-��z�Zt��Z�������:F�� >�F��`#E��0:�"�{r�^$�9~FUWN�ʍ+� g/�2S��(�g8͡G"Y�`�i�'��/� ���NR��p���駧Cqpۇ�{u��h��rǇ����!`�_ܚ��sy��SU5�C��\L´��ج!�>���r�B?�*�@��)��L ���5�����gH�V.t��ug���j[b�	f�~=C�c �$�Mn*����O-��,!=V�u7�Uѵ0)�O�o��	�9�'$G����d@h��U_"�t�#g+}1)l��>*>�&���0ܥ��{,Si��0K[_zU�m_a+��ܸ��e�{^�N�2Y�
�VeM°P��e��ge�y#Q�E}��޴�AV�h1�P��@���qAg2^��6�/t���d��#<Q�~��do�K��h����R�bT:�C��@_��33!�J�����9>����g����Gx��������x)8���`�O�@���ރ���<��T[K�(���&�|����sh�%/]���N�Q^�¢�<2U�;�H�?P��0P,3�l���uOk�392T� �Y���*��$X�E=1����H�T�%��3�"W (�5PZ����͖Xm�#��{������T���v����]	�^p���(��o�H��A;я@)��uKq�֒�)9�#{Be�V#|O�lI��d�����L���Nz^$�z�"���"��'�O�P ��}~Ж����nNu���3Cg�Z��7o)�*�-��6Na��N8�Yۑ�����w�%o��W�كq�o~̒S�x>��[]b1�Z&~�\�V���K�#B���i;����R ��wA��5.��XY�)[Q��l����'�\̓�{�B���&WB�=����-�@A ��ώ��w.��=�����A���:��h�ub��W�_^\�P(�H����c�ŋ�x~�>��#=�����D����bT���,}9��0O��#�em�� �������*�G�= {_VtP�E=�R��ݗ�UV�BdIӀ�%��r�:v|Py�����ظ��F�cS��f� ���(N^����J!��C�.��@�lFd�m|��ͤ)a\�!��G���Q��<��� ��y�Y'����?џr1�N��J^�^a]�츲	����g��3������-���ùWv[;���OU�r��k$$�N>K܌/2��it��X`�v�
1�v�-�9�a�+ђ�!����)��^����k��o��bu����>=s)~Fy�r��Qō9dh���{�%��r��`w���IJ���A��C��W�)mw�p'����/2Q;^�+W�����o��#��HOc��6��uC�(m��3ʤ��G#.�q��������﹠��Fg �S�o�&nY�N���
�@㹒�p�a�x�w�p�>C){NC1 �h�~`n-��P�]�Ո����o����*�z����5,u��%h�R��dأ��[�<�":�1����V������w�����st���V�Dk��~e_���/8��@�*�>��_1d*�;�i�`3�o��IJ�	���i,�Ŀo\�\G�i~:�w#�Z;ŉ8�I�ŕ��E���KFrïG��V�W�t���e���2-�a�a-�^/k�zy&�4��KOW�� y��}� ���!)*�e��