��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��ݷ����[h���R�@y��q�ў�BSB�3HQ��3Omި	�M73Jl�F��G�38�NǇ�[�p������$(~�5�%u=F=Z$j�����B}	Eg�~qɧծ�Ou��1�tNE106W�����g�fj�����X�jy�)K�e����8twj�%&����ë�v��X��Qe*M>M�	rG�	c�Z�Ҹu6�f8�����2�K�k����q=��3_� ������qX�W�� �;��<}����X3R�6�;(`�-~�Ҕ������	�j���w�.B����ō3��v�}\���`%,��9��>�A��!�
e��Qf��2��S>Ҏ���w&}��s0D����R��ɂ6�4�3�������`hU_��4��|��}N�ؾ[���LT
�h���z:i}�y����g�3�	%�i��e�7fߑ8D�XðĐp8L�rk�'�H%ź�g\�=��v���/o)�!�K�@�ٚl
�p��ډ�7m��������|\$���%`3�jz��P�~�{��}3�yL�vj����Y����O�`}D��Fn����$ofǥ��Q	|�ɾ2�%7��\d�E
O�r+V=)uWa�m����8]w��,f>���=ջ^�����&�s�R8��a�f�� �l��Mr⟔��ф$�!礂4a�٪KI�g>����^<�<jR�6�.3�Z�	S��ö�+�U|7������#�"��t��gWs}�VV����.���F-1���i�DT��Ĭ'��/�YOO"���e�~8���jv�\�8P%�{�Z:��.F��S/��/|�W%|�8:���,3rR'm!���_��sѕΌ�
�:ZPy�or�djT����*�VQMe("�訨��ւr_K�p���[����oE�W|,�}��3��y�w<��.$�k�eQr6��K���'��)��-TcM�А*�k����8��;1����CSW�R����{�#��	��7\�/2�ti�I�B��$��O�p�BtB��yFv���xͶ�+D�!�Ү��|�U���h��Q�|���h~�U?Xͭ6���Ĵlb����D!Q��f�[����ֲ<�:G�d��2D� �	�E1��=d������G�1�֧�����!%��kp]2ȭR�ez����e�����0vc25Gq��[���k+m%Y�	�ߑ����W�M��f>S�ۗ��x�#����2��D��o%��t=~����wy�����1�d<
��Zu u� &�5(e�����+�j}�����EQ:�@5���~>��B� ��Dt5`�V��nR��)a�#[5p��4-��7>,|n%5�KP�Fa���3�<�ѯ�%Ls�8���SKF;R�Qg\>ݍ/ݯO!=���	�����a/�R��Q���V�
i*�3��B�n^vRnE�v}�ڋ����E����T���'�Wc�#�ꑌ+زv��ُ�m"�pb����H��دE�߶�PS�����/2����F�Vj�����W'���u��{r��i5^�!�� 	����ս�(��,�l2��WIfyx�gԈ� K���.�5nP��qc3���E8I�Y�ͺ�����%#��vWBLFw�����P�΄�(��ß8�q��vT����¸�UZ�������]â��ٵ�Q�p��6��$t�Ϋ����3�Rh�ޛ�����9�H���F�$�6̼i���-���A ^�)��ȩ�rq�-����9�J%�F�I���V������?����m��+=\�]���k8s׊j;)?2%�.3����FzY �F~�٩S���㥼�\cҸ��ך����U�D�%&}+�խ�%�\��v�n��;?�_>��[!�WR�����Z�j�E2�}`�<���=����S��?�h"]��m���P�mS�O�>~)"M0��2E����J;�^�����j$���X�_x��5G8�/��Dn1c�F@ #�,_�	��o�U?B>��-�`
�&�����~�����p�͍&	Wqm�K�m��.�G	.'	x���VLҞ^��P@F����S�Ϊ�|����{��ߤ����D�]���I	fY��W���N�B�
s�V�u���&��w
�+h�i!W��>D�6�;Q���5{�R�5�%���DU���Y`y��>�P�|��g�P#/�ի&� ��`a=,Q�YUd�z�We*����9��+����pV]�G���n*�L�潚54��V@�Sm�X�vG I�,�ƐI��1��g��.CPsAJ�t-U1��_+��4	�S�BԾj��D��1|���D�ΐL螦e�r0�~�3(�UEE0��;M�����{�Y`P�ߖ�Q�5�9��'�����o��:�R��%�r�J I��G�x��Է�}�"�M����|�A������Ɋ_�J`��,ӑ�,$%���_�q$���&�P�42��a`������s���b��Ǚ�=OY����x5&�#��������BHeo��bn���\�h�����H�zG;��c���`I¿�_v���]��H��n*�qeRi^3���]����=�ռ��H���;�[���W�;��3��R`yus�H�o�.��]����k��s�aDK�������n��;W#f�s�2F��l�;y�F�C�S�c��9ĹK�q�SX c@p$\�x�9�t|��}�$�7� ̟}b�S�?��õ`$�Ї��� ���ݓ�TۦrTZ�r�j��~���A*'�y��w���B�<�o+���-k�z��uU3
����r�ʵ�Ǿ?���#�JZ��,Y���>u�=,�U�O��$}煼O>}�[	�z����X@̣k����$�2C��z"��f]���R2m�,�,0>�2,���(8����ř�ι����t(�����l�^!5�' �S������N��?D|����F���jn,Vz�t֎}�㏠�.�ن��-���;j�odq}��x[���+M�Mh�4�ʞ�r���;�0\/�lA��N�e�K�K����.���Y���J1���1�YM��Y1�R��r�ŗ���ڇ��,u?O@	��'����=�cHYCC���J�e��l}]H`!�M�O��3�Ӈg���n=?I��Q=��#T-''�x��8p��#�m�}"�^���:K�/����m�H2�khQ��L�0>wb�#y.�'?Ĝ!Ch�m��w�1s6,�V�G����DjN՘W�}�~��:d~9IM!!��?t�(��aB�|�B�(���+V7�/�G���G����� ���1)x�W��^�fd��A��q);��-���^�����$���ۨ\v�|z�r�+2Z̟��I��ug���,*~.6�P�K��X�"	$ډn��v��M�d�w>���x��ū/�F%ػ=g��YR4?���\1�3�a�;�y�6$f��Ϻ?6�5P���c3߰8z�|���X�J����~Ϫ�(���XRв�y?s����aKDQ��s�,�˸ט�gf͐�	��D���?Q��&i���b��(�����o�q�VŲ���TUsX�%������FT���Q�ލ�������X��M��8�n��q�ٖQ�?xX<-��ݹ�-{=���S)���OK?ՠd������K���E��<�[;�aSz�%�l�$�Q���K��Ftɀ��.�Ϗļ(:�.�o��?��xSS0��D|�.����-aS�+�`<g#�h�A][��j��i~�Thi)?�J�p4�\!!ň�	a��ᐖK�݂����t���݅�Rd�x%.>��(OhW���a��@e�k�Ey`�6��rF'PtU1JI4�ې);
	����H4���p�,G٫zD�^o�
}�#���Y��%�0%R�o$h���O,�BA!�6"1lC��ȭ��7�_�).U��$xx�\g�@�p[��@6l@Z�� �� ���-qP	=Q=��m�2@t*<�-���2�8TSB-��~�V�(���q����ݙz��qX��T��>q�(�9��������*̍QD�B,?^��?�S�������Yт����P���wO�����F��;�QӦ���`��=$pEzQc{��#�5��l����!�q�4���H�|�,
��u�C[��)f�<D�ʙ��"m~Ǟ�jO{�&3�iK�z�j���${�[�"�tyy�:���ǈvD���Έw��� iS�F��������(i�
�����:θ��;�R��M�vnBD�B����;4��y�0bhz&��;����|�]:�R,�e����D����^�E�C4��1ϙ�冮%*a܏��i=(k~�i�g��)NOm�s<�VH��o����2+_J��.����;C��l_|y����|K2��5���dۨsr̄�Oۀ
˔��c��e^!Ic�_�r(�	���Έz'G�ZǷIE�P�$��?��
�T�����,�=��l嵎g�bIX3��
���I�Tv��� �5�'�h`���dH��p�pK���40�r�c��+Kh��1�r&��*�4���U��p�)j��z"mP�,����	8�$=tٖG��Ik�P�`$4T���.l��H�Q90j��Ō�{ ��X�����Ty���5%���ݝ��Ā]#���UA�������r�qFm��t��5䞆�:H�W�o�f���G�P�W�d��/�O�1݊άH��٭�f:�_�ֻ�
��|����K�du>>oA]�!���QyPٙLe~?��x
��Ă�����4^��\f�K����V�4��U�y�	~�A���2  ?R����f��I�;��hŅ�Z�|Pl�{G�S�v-�ܹ���	d�ɹ�K�n|�2@B̖w�R��1���)W�cp�p}'�4&n�v�t�f6D @�)���t)��K�D�]7��Xv���'��aH�/�~M��}d�
����L{�dM���MR{g��9�4aZn�{"�aFa8N�+��/�a]��嘈UJ�bt:��3� {��? h���Xe$�\�@j��҂vj;�<��Q<i����y3��G�����TƓ�+f�9ؒ���X�EXl��$���'�;��4hf�B'f������2�����z�=e�|fQ��t���}�� ]~�4��Y�}��.� mw0��!s��G�c��(B6��[ݥ�'��?<r�'��9�s�x�z�c�N`W\�}���ܶ}G�*�5������ �/��l%Z㵈q �L�X��\��\p��S���&��F��d��l8��A\f�$5b2�\�jJH(�U�㷹i�F���~��9æ�O�߸���ho-���Z!�<h�V�sM;�ABPg�Y�\��8���6�O�T]��W����(�Vb�P��� ����}R�W�����_�� ݼ�$���t��.4�F�h8���⽹c��u�4�c���5�R�0ܑ!,����c=����z;xzoz�;K"q���Q��7а��C�>���n�`t��̲cr��04���k�bY$������$�wq	�YLHO
@O�1��%EG����@Q]e�j\4��[��|�F/���>���'�)Թo�j���a��J9T@VS��&V�د�N8�UxR{���O�m��B��Q�dM�����1���4�q�saX7B^������Jh�u��l�m�i�S��tJ���4w�%OheQ�"@�6KX�����G�
�9�Ҏ�G���s�<V�I��r����'�Ԣ����*����=�����y�lW^:?	z��"�vF���l��'n4��B�P`��}b���6^9
�<X��/��9�7��Tc�0Y{Ze�����k�حtZҸ��a��ׯ��[��RN�"�
�5�����Qx*�30����1��(�g����x�=�b۴(�.Y�l��Φ�m���ϕP�J�;��w�p.�%�*УX�^��X��-siϜ.�z�C�ƕ�T]%��i�65�b���f�4�����[�f��i�R"
�P�8��t��ҭdP*V���A�Ml�;6b�A���IZ��a)�%|#�F)zt��$wwӆ��<�@B�������Y��]u#�
��+�ܚ}Ϣ�6
��@��]� ��)�У�� ��U�p�#h��It 4ɱ�p�,b�v�z��U�Ʀ�|�4k�NDD� �31Y�Je���F���E������0:�aX��:�≙Bo �n��A����;M�#%�����c4���}���d�O��<o���
�6}D�/�6_��H��0����h�vN��`a�l2Wky�N������RS�Dv�
�R�G&#a��@7 -�=�7�BV����_�ꊴ1r)�d���)�������ErM�r���p��J0%���˳���yy7���i����A��}�Ҧj4�3S�uyzwqZ�m'�@��F`�P����@�X�6��д�kfR�b�J�2O}S�E�ۊ��ePnɠ��k:7�m1o����4� ���!����?�j��/-�3SG�v�T3��'�˫�Ƿ%�Q�et���Vo��*Ov�6�������/�Չ[�Ւ���V���!��*#Y�l�d�UU<o���l+2x�|gq�"By>O�����S�Hi��g�1�Ah�g�U��}��P9����F`G4���k���i���m6��������ёҤ����o~���wg���_~��lQ灹�N���-�ӭm��0¼k%B�
)���Xl��v�_��A�)R��,z�	 ̛��侈v�gH�������B������N��]�?F����u��T��I∜��[I�:�Q��1���Ѣ9rD�I�0�	�z�[r����J����$���Q^F��������ҨYqX�� A��щ�t��:�P��y�.�V@�3d���	�C�n�t����R�:�s�b�8�⚓�H��/�(��-�e�Zb�.��,��onP�2��W�����(�ח��E4��g+��QϨ����]S.-��m4���0�/�'���١�ڣ�iҟ�ӭAϿ|���ƽcG���HT^9�G�ʮ�ҌV|�-i�2�����ہ9b-%h��~�q� m�q,Jý�t�=��9s��1Y��A(��,T�fT���a�M(MLF�����dS^�O!�Ee���Q�]C���I0��o/#2k�ȵk�פ�P��s7F��T'�����"&7����u��,�3+[u�F����V����GV��D�H����@�*f5�,�v�2l�l�_s�2������^���+!$��f� s�Q@Ow�>��'@����'�w��q�Ȉ,fAy�=���)z���M� �O�,��
���Ot�N�d��[�υZʲ]膈'���ѽ���]Z)����4(�rߥv?��zw��$�M�0�"?;b���E0*���I#��w�G��J�N$K^��U�~X�R�zu`�ԇ�B7���N6+�	��Q�1��|ҧX�:Z�o�萐)G:��j�0d
��!�5a;�nvGQج#��v!>�g��?I�gJ`���H(�P{�T�"���C?�D��{���v��2b���7P�	F𗿼yep7!,, �޾ҹ�@�U\���[�Zc_��\��&����wB��١��:JET��L���g.��{�~gu�#ض�:Y�+�|?iI��k�$*��m)Ф^-ٓ��
���Q�?�M��c��o��n�\����O�pm�%�\[���MlY[�����K�MFjګ}g���t�g� Q���J�#0�n�n�G��k0'+�T��'���Q�+�B*�e��iSlf@�t�Ԭ?��q��iB-�칫,�iy�e��V�+�ϬE`���6}�琧�i>�U�O������qR�VQ��!�Lt6�GC�/�|=���]I��H'���w�he�O8���*3@�L�^��8��e~H�6aJ>���{�{�1$v��C��G�
4F��U)�������,%��*6� �a8��t�~��(����?�/��]A<»&=�L�š�JI 6	�.�C��Px������UB�׸\Y7��@�(�����b���OfD�n폀Q�����V��^�K�-���R�bI���=�oQ�pǗgHh9cޓC'����t��s�ˬ���¯����EUQ�\ O�����i��60v9X����ma�e�1��ي4��]VЀ:����v	h����� c�@�є��&�����d3'B<��S������{ �Yف���Y��`A���p�K`f�ݝY �蠺i��D�����A�~�v�x���+=���ft�vK��́�������'��ǂ{���� �%C��V��}�{���=�gA���E�)�SdC��7���� S1P�o�`<��eѬ*�F����\'�x���:B���Դ�G��'������X'6�|&��]����4>E���}'��=-_��Mr��M|)BKs*�I�έ)A�Hȷ��ͧ�$O�
i��+oָ�k�@�6����M*$
�t�l�c�F ��{LB/��K��6eB����zk�/I3\�Qx�@T��������9+�J��E�Ӑ,i��������?�Շ3	�.lf&���z<�_�Mu^J���`ِpHbϘ��\�N��lCպ���9��n�
L���{4�cq:¨��/������3	I�<���Z�G���ӬM|�!A��:�k�R��b��jW�bQnbB_�jDxzu�$�����t�3Qr��y5���*q��È7$�6�j�V�/T~X��2`�1���rJ��w;���D0�(�|�i��M_`�y����Ӹuw2T[���#n&�9݀��F�S�|s�@i����P��]݁�7����F�6/�b,e���#��> <Jx���x���\�}a����iֵp���c�J��ت*=��F�pd���Fu�V8��)���K!W�Yh�g9vre�ȏ~M�Lq��֧��]�xif��V�|=z�3�K�%�`A�FgG7���H���%[�R�6�oZw�D1���&1Sh(�����(q�²F�=-�]�1�%n���؆�D�W몕!�",H�m�@J ;�����@~/���)fE� F	*%[�z;k��
�E�|�bQ�K[�� �`�7=U�_ə�l/�YE��P�IA��R��B�e;�	[䡭!�}����������3�ž)	b�AHpE�Bފ7�Zi������u��`Jm@>�8k_ڧj4�*��7�s��2v%�F,9#��;՗<�" |QXKZ4c�Y�Þ���I���=�W���������S��Ǡ��f�`��k1Bu!��~��s����Bb�Qg��jR�S��$F����a$��Ka�B����,?4���'!H;�����y2�[C�}��JN��B�J���'�#�('�5(~�槱��@�7'dQ��H4ѬG���Uy��O�mJ�	��c[`RQ��N�W���g������8�E�I���Q[�	q6OV�N��C��5���z�6,�R^Y)'7���~4�&/��]؊�	��5��d:��G�6L�e;-N�Sp�oΟ}6C�l�-G:r^(����bE���h�^�@3@�t��m{��M�;�*P��h��\���gd�:M�{Uд
�S���]q�C�_?	�����%vqm��0��ё7����&W�䅱�;��G�)�q}6��4����<XF�῅���J��W­C��;7����D%���MP�/3Z,��J1�㔳8��%�>��z��!�����Ro%>e���?$7�� �S��F���)�r%2mVg��^J�iE�B�R>���a���&�s��C8���)�4�;UZ�~CQt�~����W���2,��=J�>�������U=��7���#g�1%��[`�upu�'����2��a�B�,9��箁ULݘJ��#��q�x�������/|q�[f��H��x��n:�<	' bqݱ̚2=f��$�B&ɋv0�>���LL�n�������~mu\�Fw�J�{����>+������{b��*E�6�N��L�#��)̔J��l��^IG�[r G\��kum7c%0@��@5&ڨ�AX��U�Mq���O*2�źND�e�˰�w�j4^�^�P*���A1*�|>~ȿ����L���(*��s'B�b�Y��g��ԝl����V�w��j���<`��Ü݅ p��hj2�$nq#�ZĤ_�c?��s+�Kx�;�G�i�#�vϰ��k �dA�5�������3��ρ`>�^D��!@�
����y�������R��%G�ס��19��g��k����M��)�4NA�h.}���Ex��A��^Y�UDr���;�a�Q�!�� ��U��ulfN��H�Kl�}?zo�Ƚ��Z�k��,�>_�No��Uj���V�Ƿ��M㭑���H�l"�	��O�k��C./Q�������vao��[�]�и���c�Xs.������&��V�t�C�2M�3�,H�I#e�$��6����]���?��?�e�o*�>J&I��i���ɱ���<���"�y�Յ]b���L���F㢥�K�Z�n�~�Dav�=#����������m� �:b�U�V����[dE�".	2m��y)W0<�8!���U�/v����a����[ V��������.�>�IR�W����r�a ��}P�������}���ŬN�Z��G���䝊��d��"1��	/K�L�6�#�����~�����]��IH��h<��|��9���d�+��Cum�����q��I�O�P�҅��ޯ��v����)�)�o�!)գ	C�;ͷcl������?�r;7_c;��}��XJ�yF�kuiU-�2�ݲ��VG�Ӧ�
+˾\=vT��6����{����m��c��-Qx��r*4�ƞ	(�TwIs̀OP�V>�E�mB�CbU#Y��Y
1($�ۋ}\s3v�=�����v���2���|s�����+����{s��3(�U�U�oh0E����q�n*jl�G� [���"C):ړ����x]�cZ�;@�	
�������'����`�ЍyeĪ�4��m��M#Z����KN�L���4.�5��.�\��6�/�f]7�g��el�;�o��������A��鞒T��5#q'��5GYr=�W�
�ݗ��H���	�K�n~��a��N]�/h�4�rNlna|��U�|J�||�E���\Gv����Ky������u~)Pfa*��_]�O���44	q�����Dbw����UY�U������v�:Bd>���+��������w�]I�:�o郤���ۂ�O��舘�D�p��$Ѽ!Փ;�[����v:���~X���Sĭa��o.�qc�;-�B~���2<��gw.�ߞM�hQ>j#���6�Z��jS����u���3�훴^��)ol���t��H8W��[�.h�� �\���2PCQHJI67&�??X����k�:BƣƫL�羙v�'��Ò�쳮d<�8 4�/�@�e���Fn9R���NL�K����X�jw�i�����$q�oZ9H���şZ���,gT���L�M�rO�D{���]d:%mX?�Z���P��.�ذ.*����Φ�u"�QɅ�^������)_�?�t~��i-��z47�%VO�-�F	|Kӯ���|c���Xb��o��f9/�g��|�p_���ǳ9n��D��_縐���ӫ��/ӥ�A����	���M2�.�i�0��m�M�:����:MY�T9��xq�����@	J���Y��P����N����V%�M'$�vJ7�0�2�b��2��h
?sg�H	�FZ�QV�JY�	�ʥN\�Ҏd&T�d�f{Tc��-�0;�1:F��0�MJhb�㇄���"�� �ac��;�w��L��'�G#��qZ��v��#�f���A�yI+}pDu���#ed�#�R'L�j�� �U��q�1�5���|�����RrیD7(1Βb@��x�Jj5��"�(̐��@�߼�<Fd7����ْ��!L�]t�?�I��"%z@���uAPF���l-Zv�GR�Ͳx��ͥ�h�� �|Lc�x��Zq{4��J���-M�ZVY!��PwF�߷�vF;^@%���t�|���;N;�g�D��8ݎ3J�uFj��/�-�ϚcB��吅�������/o���}��6�����"�tOA~5yhK�7O�K9*zǞ�V�7N͹v�J������S�4��ڇ#�]Bt�:�jMB�n��2�H�3� ��X�_C�OW�EْR�ٚ�4e���8o:�O�y�'��9U����R~���Sލg;"ttP H��:��YRӒ�N�t���,���2�)��y�9G��)�l�r���eMrx�k���O�?��D����x��qz~�.�%�����	����ۨ) $�h'Vy��;ZJtŠ*?X������%�3
�tE�|���q��
	pa����5u�G-��V���$v�5��L�=�9Ș�9����IVp�dQ�%F��)��|��ԩ2��;'Dë8Q�L��Gܴ%?G|�M����j|"�X�7���]��|���B��톶9�$�ۡM�>j�� KgM�AmM�(��j�Q��^P��Q�6������HQ�9�C�4�$k�Ii������n
r��G�c�2������jA��ǘ��*�((*?�/�A��eԆ�ـ]#H�:�+����Kj9᝽eZ��&F踟�3N�p��&�����x�������'�E����a�.�o�n�Qu�|�7������*Ț-�R�%��SWI\�$��r5����dN;�R�j�[�/��{</��n����>����!����eG8 ������V�Y��E�
���]&�Ru�8�{h�ođ��i^��Xlΐ�ɽ*	T�����Y��73���H~��e�ֱ#_����F�;��qe�M�7*n"<�
��#�rլ�ǱL������O�L��h\��W�x �h}�̷����E��]M��x�=�W���g���6&��4��w:pz��`�<�䤫W�S��ڠ��$����H9����*�պ���z�m�W���H:��/���BaXu�{���'���K�Ԛ��:���!���']XN"F��wm��MY��(���5`[#�ISV"D��{���I�譸K�}��:kV���9��Z�V/R�K�����B�@����Xb������M�l�ӬX�D0�T�>-W�}MȄ���/�*�ÿ��1�oFJ����l����쉌���f�i�����wR4�2���+x���V�$]$��ߨ���08�Oy@R���҈�ģ��c��xT2���9�l�F�1��B%0hz{�K��������ATH����uա/��`��Ʌ9w�0݉�S��δi+�;H��HL�F�O�y�)��t�1�ȕ���8��~n����x�h�c�`�#�Ln��W�=�b]����y�]�H�8� �":6��m
�H:\hMp&��'�������*z	r��u�/V�X	�ws�|6������?�W`��q> �H�����"_=g�=2�<�	F�m%�'2��6�&�ǵ)tY,Uļ7��Ȓ�w���\��M��yT�weQ��� �L^!����-��?z��'��l�������@�jie��&h�B^�d��=��i�q��ͬ�٫R�4kD=�N�"��[�;#FJ/�p��7xM&��f��P6�ީ��������0��	�(�6l
�����HQ!�z��Wuqš1�����R����d�z��O�Ǝ��P�(��ަ�u��E#�� y���$�4Em�D����2�-��_ڰ�7�.GC�X��r Z{���ln��0���S�9�=ՙc�U��Jm'!�6�-�Iא{
�|U�A�B����%V�+���rM({ܣ�A
��K�Daߝ)f��l�Xq�-Ũ���:�D��H~�{����O���;�$��KUu����k5��s{:ވ�Me�D�G�/t:�?a�,��eo����g�D,<����s ,���T'��2s�W^~�;���;\S�T?�ߣ�#*/
�M6<TJԢ��ȟ~�ZYuqc:5�5���ex���������f��7��[���4I��o���G14O��7����t�k����yo�8� |�8�V�_�V�,�7�4���|�.0��,�ndQhM�G�9@-�G�Aj��X�m2�_�\`W�� ȂC�`���/2���E�E)Ӕ��	kO�"�^��[ 4cҺ�pB��+��Wy�L0��dBӴ�ӈ�o�'`��u��J��}T��t�7��^$��9��gՋ7	0��9��4��mU�������qd��������[Aߘ���RS���f���~ϯ���1�/�C!-�PX5��X��F�m�<���XS��}���~���h,�FŒ�:�-��O��ׇ��ԴN��yi%EG/���I�솫�X��i�N����>�<8�{6o⥘Eϳ��TM�Bh�)�
�+}�u��`i�:�+�^��#���5�^#�m}CV��82I��r�D&�`V5��0�g,��y��u��:a�F<a�Uq�1Pke�\SA�'�k����Q�xI��2=!���>n1	��uH��|���\�t��� �d:�):gT75��t�3k�rqw>"�;���I��`Nnv;O��-�XPo��c�EBۭCT{՟�<��<��
� ~�{�/�p�w�.�oL��<�㾤��*b���l�����9>Q�2�,���"�n'��u��<Ek��&CP�Q��AU&���,ok�)[<[3�{��^6��|%����+ı��l�M�nv�q|0�,�Ճryދ�q$]�P�ނ���񉵐��קj��E�o??�m�J�0.�L`�|��v��V$kE�G���c�~/JO��kR0����~�[�����D~U.k�������0�T�j�$Qg�s��,��Y�t�1�>�".��w��0��fk��$�Q�}q ^��C���"I�d$߹f��?�<�Y��䕻�� �{U���MgH�^�j����WW�u�p/�zҫ\��CC�A�h>�p\�bk>��B�(��;Zr�;���\Y~,�d����*}d�MӊJ����,on��,��Gƍ�Z�N%[�;Z����RIee��"�!�`� ����x�^�߲�q)�}2��8��r8� #��vAk|X4N�n���٨-����3P�l��ܥ��`l�.E{/]�Y9��2��{l���=��ER�S~t3t^�Yp�|}���	r/I��ؘ�:���u���Pr���U�}��n��xq��}��/��Ж��0ѳH�������}W������h!�C11�B�9��ސ6 '�{��<:�!X���j�K� i��g��)���|��A6��޼���Y���V9K=�h;T��Z)����w��/���Pv>U�5r j�>�E�4Bt�ִ��i�F?���?��|b+A�Q��! �8�N���,qX��d2\���jI?�LP¨�{��.��Һy�w;
AG/��F�:L�K	,@N�C�H�T�rK{�ŹxsVy�y��c	��t?�Z��];^��B��.�vp섄�C59�D{��k~#3a�BP��@�����^"�g��ԡW�*��=�j�{�%��-,��������3� �-^}mv��Jk���-�)#�o/�n-@��zn;{�>*� RIdt�����.`��f��I���ѩn�vb(�X�����!
xҥ�T�BY�;��e~1ʬ[�B�$y~���{Ej��6�E�up���u霳���W�C�}bXv�}�68�8�V��3�6- *�oX 	 ��`����o7�!�ϓ�bᎂ�4��WJYoE��Q��X�A�7��ײ�H��`J=T0��J]d��G��:X-��|P����M��p�Buo�}�P�C#?��r���hp���&/��$.7 �]B�^���%�ߊ��_��%�TԷ�ӓ�/������L���\(����Ŕ��\�/�;N�p�j�#4�h?
\�WY����؁�?����0h�������|�S�XLK���'��#���v� $�a�g2h�VȵyO턉_!��b��T��2�z�����L�Y��G��r��8���������q�4�*���P'���'��3�-�]�5>�*p��1�.���wk��be�D��F�po^)�� 7�BU-$�7ge�mY�Bw�����hL�q�;��( �T��Ge���< �I���͗G��l����ܻA%�F�I�Тn ���$=ss.JHI����M�`$�1Š�E	��Yf�pR��7��v+:��
����W�j��;T͡������@,^>njW'3�TI��T�C���C���^����y K�9��heǎ%��
�A��Ը��$E�4Oi�ɽwt���p4�ҁ����\C<r��\*ݎ���m�/%Y��hu��O���4�yj�jv�LV�R�W��(λ�Q^�Vn��+�\�bD�[�6bP=v��r�`/��P16s������y/9�Ҩ�������La�@�>e{�O��\0��`���V~I��M_َ~stA7�L	l���}]I���m��Xi��V�Z.S�i��>��ޒs6L�q�f{ޤ�|z�Š�s)JՄ�X��ὖyE��;���*�7V�='�o��z���-Y��=�P'���7gaHA˕(�R5��g�z,(�5G4{�Y����i��E~�y��3RR�>�طW�S��e8��U,c����}�����oV�r��w��/�T�V|������{hj�hoiP�31��_�1����cN�}�V���^�1�*�������P4Y�\efS��W��e��*�3�$�6Г�3�7\��N�jQ ����U��A�����w?w�Q3?��2`NZn_���J��F���0��f�6l֔�z�혹�$��t�Ӌ��=��l��`�]O�e	�Da;�^� �~6��
%�cd��o�HM�F�P6a�:DC) g%?�_%�tߩP`dP�0��f�JU"�+0b��*���`�8�?�b~�d~g�JJ�|�2{$��nڎ��H�q�b�Ĩ������6���*����+�����z�p:�Dz�hf����l9��Ȉdp��X��E+{^F��*�ѦuX��@�a�/V���c�n��&eu/^���G%ф���?�l����ј(��4��r�ū��Fh�������=yaid �}�'sE�����',�*p���X�wqx�Q̨��FI�%�xS=>�43���1s�� ��-L�z�u��\;Z6�O�ْL���\��[z���*V7զ,lR��փ��ym���)lNK�џ����
!���AM)�Ҍ�4[�N�-d*�ڌ֧Z4v!�Ob̨%��8iH������+�G[��8be�jA�iU�8���;�/ٟ�퀳�F��rv�)���zO2:y28�؋��HC�*J|�'�I`|��IBx���Q��ܯ7!��T^Po@ԭw�)/��~K$G�Ӣ&�n�t��<4�tk��U����f���D4�pСD��5��h��)]rOܕ�o��憛C�x��:B5A��>��?���# ����֗/^@z��dަұ��;a09s�O�GD+�p���NO���H��F״Y��Z�h�!7�A5g�=K��������Q��v-��T��\�v㨧�M�PF�]j��gI%vWfSC2l�as^m�N��fȴK^?5UZP�L�ʤ!��K�k$��_�z�t�.�zjm !?��=r@�7����㻓d��D����,�����$2�u�2�Pݒ�,���D~�	�rG�
��e�p,@���*��Q�K��h,yN�R&��ޣ�<���77o�h���m�� |Յ���e���Y'65O����f��?�᪉��)]��Fp�"�6�8��-i1S�v�2�>�:o��v,=�؛�Hqb���򶝨�,)�����*��L����E�G��K����Tc�Z?�!Y��Ȍ?�O7�s��9;fS͆���JN�9_����Q���޳�ZR|�֦p���Z���,n6��^����t'pMg�:���Eň��2��v�N��c�8�0��Y'#�Z����E6�
f5(8<�EO$��k��Bz�pZ�V7Zt\iw������b��vD�l;����4A����g�=?ť��HW�4!�ξ�Ē�>/V��-���}s��s����$kfu!�'�*�ft�Q�M��YG��:�	�2�F����CW��،��<AG@4S���ۇM��|M+W]$8�.�4n�'�ALE�B���H��߱ڭ�R;\�_��6Dq~�x���I��}����gC�,Ag	�]��|Ob�I�r[9ݏ�ǎQ���>;�^i/Ί�Ӈ��0R��KB���D���g���F����m�X�y���4m��.�4R��/(~\��z\�_��X��m&=����!�(��TW�]�2� ���r���13�at�Zs{��A�t�D������\�Vd"�
P��y��7�D'��ߩ\�z��a$B�3S#`�y25�����M>�(*{��!��*��6��'L{����`��$,��ce�t$B WP?L�����yi{T�sn|eh�R�ņ�k�Nbou7���;�s�|��y��8&�>���F�`��k�4�U#b=�g-"��̍._JB��@cP٪�R��}�t�{�S�/����$�/5��t����yzd��}ߛ�H���=�h�T��8�H��`/2ՍJ����۶}o�$r��R-{]���r')�vfbj0D<�|K}�.}�Z/��/�RS��Sv��|������Ht^�J@A��$9a��� /g}]�W�r�����qBB��@�p�R����̠d'� %��i�.Y"�\,��D4�nAnN-d_�Tc��1��.�������\��0�P�vJ����,���>	j,`��d�CƂ�a\�����<ˆ3�x�T���y�nG2 ��2 �2}�������N���.�
�(�"E`�	{sAl�^Ԟ�dO��Eົ��>�VaX�D����,�eИ�>��P��Tp�<����L��Aև�ѩhB�-��&�P׵5��A�P��<h@�O�xi�>T�����@m�n���N�֞k#�ܸ(�F�͞,�Ə�~>s�*���7�I��I��"M�`u���>��4Pp-;U�rzLL�YZ��~��5����+Je�z���^�!�6�r�潚��~���G`��A!1�sA{ۋ��B:����Dy��[i��wc
�}Sz܅���(�Iɓ���y��%�9��dP-�q ���6��R�����D�ʹV�<�ے<�!.����AO�u��I��;х�o��Kp{)
�'���\�؜��u-�����"�|�I���+D��-
�C��U���8# I���ʀ1�|%̊7`Xܜ�h"�ױE��jis�W�n'Lh� ���pbEGc,"cZ��@%,���֥�F���S6������έ��n�kԲP0*/�N��M�	N�F�~���C�2�	G_�N����8.Z�l���9k���d�~E����X���EI��t1&����s��)K������]JӏX[�y�C�Y~��"�1�8�������؏3#�V9ra�{NMF��ǈ;�]5����b"9j����?��6�Xw��Ͻ閞q�X�S歈|�R���j���>s�B˼A�&�u��R��?��;&��/o��R��@͖�o��j��U��d:[�c�A�ˀMג�&D+�33h�.'�Y�4Ϲ�p��Gp[�����m�ٸ�Lmo��~��ثc�x�iyT�G��>���	�����q�	��dO\��Rݢ��� h�B5ڱi�Ͽ�CBkM���ie���鸗�UG�t�'�Jh	^M�rK���[$��it��{�ߚvv��k��y����`�~N*_��	_[�}bV�����]��zlQd���j�+)%�7X�*�7����K�U��O���Ywc�ڙ�����X�舸	�Ya!i�qT��:%�і�3"%��U�w��:�(��I���#5�L�|������ܿ�x��\X���}�#jG�����Ǉ�<�޽���x� -l�i����Ch�0d���򲦮u���5[Dt�Hs�/���)Չ8��ۧ���ye+�4�)7Z�c��8�����$���=���㤋I�,2k��F��V!�np;S�?W3�!IE �a��u4h�y�� �M����!�Ɵ{�LzN�{���G)���iż4ZO�	�쓾��hŉ����2W�t��DC+|�A�2���L�	'��g5Ь���h��{}e����3��l�q��t�_���]M��$�5k#$�m��]��Qa8)}؂"��}pA�FM�� a��O�
@U~O~�(��Ĩ�kitX�@��vI�V�f=��Zmޛ~�}`C�{��Mp/�̵	���`�������|h�ر���t����5�ڎrR~��3TK�@T�� �g{��< I>�O1�fBG��_��&�@���Ӓ��Y�Fui�Xھ]�4m����#��Rpߡ��/�J7z�^:[Yjǁ��`� ����,*OS��*A=+C��8�R8��/�g��ۅX'c\��%G�\�5 0�����>��� $�x��)��E˚��V�G\�=J�
��O�&Ц3�7K4���`W�RPQ_��67FX�Z�Ěb�w.ϵQGXΘ� ���}�g����.�Ѵӂ�� ���>�b�
ᯧ�$-	$�t�aIb�u�~�|��t�e�>��G���"\��6�c��Q�Y��?K�1�� ���hg�C�w����26*�{���Pe���l�XWE��/$Ua�TM@	�I��6�:=Y�^r#|,ׅ�P�������B'�������|��M�R�^�Қ�b\��+Vkxr:z�vy��}OI@����<�Z"����>�މ��wfᏉ���O��2�$G�ڹ�&!3z��9�Gڂ�L�(�gj�k�����q��w��^���ƕĦG�,}
�W��	l���\�������Z�	/ZSF��)>d��r8���q�qd�X��Y[Z��o�Ez���Y���7�f�mFg�%��r�o��=:Ã��K��:>ө�=��ߑ�T�
�Z��ֲ�I ��������S�1�*�f�}�=�ω�� 랂�/��O�A��⎰��H��l�S�;1!�3us�O�N��p�jX���|5Ԉ:I�
�y9��"�A:F[�7��ot�y;N�Ƶ��1��lJ����/?��b�Ng
�tف.:�E��%Ekb�>$�~Q5_z��-u�����%��������� ��~��<��-07�*F"��z�k�F�����ux�����_�^̎�PJ�1�Rfݿ^	�0�Rg������|QH1��D��r!��ڏ�|l�w�G�j/wGӞz����)�f�l#����n�;1�;��/�}W��'1��^�72��#h�	�N��̅g.��g$D��R{�y&#|��&kr%�@Uw�"�/��;����E����|��_�Z8L���10��B���~r��%`gR�$A2��z�i��YE���W	Y�p�)Q���=�<�tSߏWT�ȱ<�vE#����������������%�ͽ8}#)G%jҧ�|��9i�≊�:G��1��1����u$�e�t"�F�����IG�@>�<��r�n�ŭ9)On�K~Y[��=��%$V�w�t���=���[���|,x��6� ���+�rs��i%�oB��z��~m�ʃS�GMP�)#�(n���� �\���3&4�6��`!��k�Ua�F�K�����T{�쌕�������ڣw�cg��]F��ڹ�j��RI)�Pi����:u�o,͵��''6�y��҈ '���2�妔�����y��>t}�@g�����Կ���a���N�y"ٜV��@�5d,��ȼ^Ᏸ�����(��2L�I�Ź�)>�QZPSw+��9��K	+bi�Rj!�7�L�3�%mQ��u�0uMޯ��$����8���7�g��:�;�C7�y�8x�2��.�:�fHO7���8���M��En�j�L{���XTXp]аʢ�9X+�|��0��>�	"����@��ߏ��`�=
`�p�ԥ���fܾO_3�4 H]�`��ԩ���Lh�@7z��:`s�ˍ�r��W��wd�6���?�G&����4��S����t��r;��0(�w=���h�����j��ʬe��@	�ު��,�ڰ������O�V����cX����J
`ԣkY��/;�����ޒ_&\h��S�æ$�@Q�9x� g1�gcų�h�QV��Wt�@l�1��o
�7k:
�������}�A��E��#�����"GZ�dSXO[0�9Ϝ��y�c�b[�V��.)
�}�a%T؛�~\,�S�1IR_9~1@x�2���1#b�/o7�)�_ԭ�~
��鑎�K�5���-���4�Ua3^��#"0	9��z(�gG�4�Sл�f۳彪��G���,G����md�"�_��-�ZP��	=�,�������9���]�㳔�ge��[MשbM��O!E�'0����<5�
6�S��l�O���RJ�U�r����G�����ZF�����̃��J=�,��dL�y~�n�Gs����c@4�'��Oʀ�~4��ڼk���#�n��2Ce[��W{XU=BH�2����.�P$9QW'^�e�#�&Q��,fBi�x�B�	0wM J�9�;�)�;Y%�����?�~�ݺ��|�Lل��C
���y�Bs^hvׯkG��m9u��8Oy�ħ!.�M��z�3SPV����_�̽������sX������R�&R�Ɣ���v���(YI�5ΆA�)�Dy�v�Wmc�ni��:�؛W��fb�)"�>*��DZQ���;��.�����S� �ӭ��+Jɰ�#q��s (Q���*�{V񯃏�{K��DM�
�ЏԌ#�g{w���J��=g����zNF��u��@�zV�}������W����A�"ӕ�S-�x40o ��oM�`��8A�P�;Fϛ	�G����_��v[e잓񜝡�lv�%����J']�.B������	aBv����:f�Bw9����l�1�o���ҁ�@Q�P`<ޫ�=y���S��N�a�w��@�fZ!K=�>ኺ��a�8�F�Bd�1�4-���4��5g��'&�0t��չ���]͹�f��Y��(�J�9�r��IV�ʎ��{����2�dvq�	7!�P���� ʣ�kf��]�>�Ӿ�d�@iu&�v���;M�����T��ܽ%�4Ȱ���E<A&}�����T� �M��|y�&=C����j*�ʋ��Ӥx������ӓD9������68����X�Ч��D_v�!l����݅��A6|�Y<�[CtL]�F������8�ݞU7.�<�7 �i�]��Q?uX@���'1(F�ʙP�ҳ"�_k�����(��e��e
YӁ�q>F��`q�f��)������G�G� L�uD�:�9����	��(�w|OCN
��uv���d}�$[{�l��)Q�-�����!��D��:K�PC�!�+�eϘ��cT��Z`���ј/L%�Ǉ�N?gt�xE$�@ZT ��s���?:2d�<�^d�J�Yt�Bc!(����w�#;�5�+������)3�|��w����ȓe_�lx�$���z���l�֫��[�h�S?�"�1Z&�x�#���g͘�B}��4�I�q#&g�i}�tr�&W;���Q�X��]���/�A��|�!�5:Q|#�Y�/X=?����O�,#������� K���k�v�	��5z�B�h�~k�#�����t�5eK�
|`��*t�E ��ڴ/=O`�u�!;�ō�$>�Ku��`�tL�0����c�+�l�O��z3Xٛى>�҇��XDv��aI4楥<|�e�`��Z�VXlAX.=�Gsʋ��w�4z,�"���A"F0#u�`5������n��6�0���*�>$��7/��|r�}j�����/������eL
Ái�"��Qh���bk�NMw����@C�ɵ��e|��.�Qb�K�T-ע-������Uˀ�j3��n�R����l����R�ѵl`������F�?*+�h�c�\�,)O��s�d.� co��(�l�&ɤ@�K�/��ѵe3)�B'MH�Y٭^���r^�,��Ss�߁M�1�	*��^U��8j�A����*{�D�������}og)!��x{�kPSL�^r�Yg [�dd�cu���џA��%J ��	��/hS�C� �2uDk�p��n���/Z)�\f��? q�����:}�V�Vp�Y^[@�iꂛ.9n���F�<ki߂ �fg��N��� ��P�S���͉�7��u��rj�ꝫBѭf�v�8J�L?H����uw7�t��&'�8|Ã�k\)�׆�+������՝L�c2p����0���c�V�I�?H�cW�b��9́9��F��X(p鋗D0��8����;W2�⻑�ח� zϜ}N-�}�eZf '9�V�E�ȀsQ�Dd�Ȗ�K�I��r+t�H4�6@�ϔ��>R?��H��A-c��� �֕+�8�+����=��^��<ޅ�1����|#q�l(\T��:�<Iy��)[q=�H�X�H���Y��%TGe����J�sK����aP:E�_�͵c��o~LHȆ%j�hY��G�������t�a�?���B*2G��{��!�;|�T�x]�勞��ǥܦ��QJ��Ns�o��Ā�~ڙ�Tt?T�F��u��瑾��=����h+�Z�/�爏F�r����5��V�X<��;�����kRL���v�@ty���	�+��̴�J�~ƥ� ȼ�1�2�u�*�^���%$��[l�V�+s$�Ѐ��3Lڟ�����	�'OjB�\�Y��u��z��v�l���T��7���g3H^|Πƻ��� y�Pq��M�V�;�尌t��ބ�(�Ф���݂�ڢ��Ț�w���\�%ܠcF�h�A�$
�\*?�蝯�5�l��7�SE���Y��x}���e�M�Ҕd�iSk�H0��W��OOX2ҠVRjS+C��
�&U��:c��m���%r'�<�|������Uԇ^��5���c�a��&d�dZ#��e5ÿ�\���1��#n[�;��j�MW�����������(��y�;�[ c�+>ko��Nm-����������f���@?͂��?�,1�@Q��\km%�(��z����G�a�������O*z�6���e�HjH���K�NS�VƐd�
;[��FQ�Z��P�zUߙ�86~�*!P��V�?��OǍC�#�����@��	�_~�3-��c����־��#����ST�-+�����z q"���0��2�0�#�4+;�P��a]������Q�h���ʃ�$��zI�T��[�G�:��2�%o.Hq�K�W��P�WJ,�%P���:���B4��AZ�1���Ɠ����&��j�0����FW�;!�sڠ�la�Sj��-.yV27�h������-���v�w�;����b;��� ��&.��{��K)�w��ˋD3���_`�4�#��3��co�ܺ���Z���/�`⟈Q!�t�:�pĚ��X���$�6��mA�=7��;�Za������*��k:i���|�bv��h��l�;I��!_��7�e�2������]���H+��~��<��_8�׆Ps��B[l�3i1��O�S[�u��LgC�IkP�N˫�s���SNa�R�Y��0���^��ا�t{s��VY�#M��Ԯy���?��i���	*jդ�bX��u++ ��T��b1�T�٩�|�!М�HtsJ�˸�1$���<O�MS�V�س��\,�ːeܷ=gT��fo�;��ҝ��ǁDhb���8�ui.��k� �.���{�^r��Sŷz�p}n%d�M����;0 \��un3��n�i�ج[�����V��\�1�79�-Ç�b,�\g�.��@JK��KBzbC<<P�m��|n��gs�S=���ܨ9�	��eV��`��ĵv�)5�0xӡ��WXs�G����|��<�4Jz���5�[��2�В��{C�aZ�I;*��Ü̕!��~WI�#�Ew�[ս�Idq�2��۷���(6.hIV�����=K���P.��#X��Bm�{�����]��.�p�{�l����۫j��'��oH���R��ט�d�5݀���}oh0���>���(��ۣ��2��A���
��nq 4V�yq�-k�篲�
s��9US�)8a^�%�$�>7�5|�eJ(�\L-�+��m���O�{vn��-%<���k�;�J�4y�,�y5�x�T0��W�D���W=��|��wV�������x���w���}b����i�`z�.�İch�Q��Y���R[��| ,l4��2��7�7]��D�қ�w��l�Z�ق ���B�f0�;��T�026�������9�ݫU�9+���@y����rԚ�r'�Ҝ�;$�)$��(K�+���pH�HǄ���hE�.}��=S&Q��)�n�Bݱm�16�8��UT�`W2�����@_��sO��'!ۭH���"���a�����+Z���94Y���0AB<�0a/�#&' O�<95>�i�{oY�R�3n��b�)�݂��D�-���	�
y9� e�r�D63m7�
� +�Q�(���������r����8B�5��/q��D�N�NAtx�� ��K��Q�M��gU�O�'�z�bSy��D?�߯����)O ����9���5��� �+��I�6��a�ER��f!�N��[�����Z[ ��/y4I�-o.xB��٭?��0�*�V�X�.�hg,ԈT�I9��:�2R¢g�c�����y�B`��ZE�plf����V�s �р�N���V۞��sҕj�L�r�����/^W;�r'l9ǻ�Rh�6]F�G<�Q��?���Eܚr�]} +��^�.��>}��׃Nl�&��;��i 3LR��i���	x"Z�2�T��7"s�l�f��К-��8�)�K�a�D��"�q��|!��]����Ŭ�E��V��uF�6�=B�Nu��^W,������"[�Fa=�E���wEN�����IwET�<$� ��-��h��1�B����H��)d�t�`W����̘Q��0�aP�돢�@F���r�b����z������K���ÿ���-� ���y},2����+^{��=�(�M��<���a\L��芛�Tf��:�e����A�T��s��~���g{U��[����w6M���S������xz�&$����79G�E�D��^2�l'C�W�̿q7q:ml�kŊ�;r���{Ww8:`]^��$����X�i�X+�-{��r%UQ��D����Urr�.�H';�%�����O�:��y�OP�}��ۣ�Cd�hs�<%��閔uX
�+V��j����6���i�8S�jX�-�,�`��Q��Zh}Mc��%K�b>��ǟ�5�f�B�}��'#����/��Y�
�J��t�(0*v�8��E�r��|%��z��ZQl.G�J���E;�"��I9N�b�5���ܪ�Ns�_��0�5���|{�p�2��T��8�X-7�����p��(H���sa;[�xXd�Y��g�����Q���^6>ZCg�R��06�l݆��}���e�vߙ	�)�y�y3:(�W�@x��ְ8v�
���,6��{�V<�,`�8�%6=��-~�ZÂ�����Z��ݏ@Ι�ܔ]�QM$�ݻA����'���Ø'��h�\�ÎCT�_u�|�8v�9d���^_a-����A��t���C���j��:�$�TUM�JWhoX�t���h|����z?�[�sY��!���K5H$���J�^˪��y�iD�.��F��63�h���g!�;��3ݍ����<s�D���9�Rê���ӑ����/ۻK%�#6 "����!���v���өGx�Ԯ0c��g�~��&rQ�+���0���S`c
]b��R��I�r��?���[���x�q����#��9m�Si��`s��&4��o@��(.�þ+�;K�:�ٲ	���`ܿU;!�g�T�ЛXpg�;	�4�hM�}����?.1�-v�������#���������[��Щo+��44E�"NDQщ��D���F���:�(��ʬ{��S���)��Z����٠q���T-P�d8�Ni��wL(W��R��S�=(�~6�ʥG-zXޟ'�M�=WDI	���ݲ�H�O[�Jv�/Y�R����������s�9�9O��	@f󤌭��Dw��ʆ|M�R�����>�	�Y�pwo?�bX�"2d�a6Čge����qB����:��.#w�!O�3vv�yK�ޱ���^��WtSj�����2t"�W�	>=���p8V'�tr�9	cv�D���nݱ�R¾����G��kW��G����ʹ�����Rv��)�ׇ��螌2o';��>댄��9v0��9�<�K(�.����{��q�?����Y>O���������t���}�R��IӞ��&��C���^Q!DM�I֍k���ʬ=�~ĪOD��r&�)!0F|t�R���ׇ�pz�e��a!FMKr5�<2�u)�*v���ђ�~����	l�;�c�!�߻�!Fw�)	z�M�?v�<lۣFWtۢw�tp�oE�a�䇣D��~��t;��1>(�#�ӌ碮z��Cnq�j&�gHs��m<+��1���ַ���5�aTɜ�"m�S�(?�%⏗� ������/�̵b�^��)$&J꽘N�~(��T	�v+ae��܋ f����ߋB�?��?�H��]ٹ�,Ff".�ł�Z}�!������kj������R7�m�pO�/�S˭�)�):��[�3ǖ���VE��&b�Q�5�)������e�%�0i����=rQ�N)L>���?U����L�q{���-��3�QC�^�1ܓ�<^�q3��q�&��>Jx����2O���:��1����*Ѝ�J���D�V**�e���{Â�"&��P��"ۊ���Y��f�Q����8L`�s#�
M���O�E.LI�[�-���>!Q���o���A�����#�hs|��
�����a�[k)]�b�A}Tx�w�|a�%���h�$��1�i�Ƨ��q��>��m�=�vH�C �Q���g��2�rL�12>h1��f��J���O+I&X��U�@�8�����j#$�x}|�@�(7n��>��>�U�LEgDq�k@�.���jM�y���w����d�i��H���ڥ �O�v�8��EƢ��AJL	�lV���G4�V���m�z���0�}8��p�i�R��K���)�-3^�s7�~����-�0H�ŶL�k��=t4w�.j�P^�aaLcFn���V��	l�X�Բ*��Li��
��$�Mb��m�}*���fTw� *<�O��X��F	/�ך^ ���+y��<��h��C��*�[��nq5	C٥�Q�?�i�n��^�C���"i���B��6,�?�����{�V���T������s@����=���~�5C��A�<�)ę�*�́�y�yn�W` ��81��@��FI��xO��Jq䖃ld��,���W,�|�[ �͘{��l�AUz� ����f�L����yK07k�T��v��~�M}�?R�R޿<��%�6jga�s��D��׮���'@,�#؎1�]��l�@�M0��Xp/㽯�%��1���I���'�j�<�n1���\�'A�}W�Cd�f󵜩�u���!�4=/y�)������Ӵl���[�,�MzT���|(=E�{{�~���r��i*,�sC����Z&z��5�r4��M)�=��R0p�p���4�l1@�'� ��å*�D�J2c��:q��#�z�qk����-gU��4)�{�@���iY8��I_b��F���e~��W��%�2oO���@r�CUǺ��Vݙ0�{.��������iAZ��5�,���+"�p5<V6�&��sm��i�<�y���Bo!RҗХJg�v���|l�P�C+E0�W�9ܩ}�F�%t���s`=�i���i��J�ۋ�d0��Ft�_ɴ��)���JamHoNc���gN�Mr�>�Z�[���Uf|�W�Rb��R�)��J���8Y��<!��īz(^Y�KH�E�m�"�f��V%��
�m%��Hۨ�� %�=`i'M3�p-0<Y i[�"��Q���(����@��̥v���M�kلX诓�zI����
�g ���X?z��j����'_.yh���,���]��Y�R°B���3�8~x� 9��/yQf����oˀ
df��F���^q\�w����B�ӷ
K!��iQR;��-���kE)�J1\�z��g|�٘�Ož�zk��J<Ŀ*
0ˣ巄����Ab��n�{�?����Ȧ���~*�JN�~>��~3oN0�J�%d������?��L�h�p�M��s!b7A��蠠�ZW��*3 �����1�_����Q|�Rn�'���yxY/��
⊣�Q���z�n�4���*�u�7������}�"S���@���}8���H�A����jUpK#8�r� �ө7��az7��T��Q��E�*���j ���?��c��@	�Ow�R1^H�D��f�T>�$��^y�O���������")4�֣�*93�j3�"��	��x_�ՖpT�!K��Xz$jUd�P_��_��2[;�9! Ɠ잧I�������=O[�i�4qZUnM�e uO8�9@�T���R�Kk_�OC�$=�[..��ݲ�Rh�r��0�d �@�7I�܁Umo*h�W&Q
.�V��i"�^[We	G����������[�>��j)��[�����h���ɐ&���QNί�����B^�庀�8�X��'K�� R����%�B!�V���5t3�:r�>)d��o!���W:LXz<���a6����.b_��_�U$}��E~BZP�9
~*oL����t���?�a���FY��V-x�;2����5�׼<o�}��4��z��H���{Djs�߂���)�i�O�&?�0<9��l�@�)��A�J%|�l�@��$Ae�+y��p�a��v/׸t ;�`�c%��e��M�KU/�d�c�f^�B�m͗?d��a��+���� -6�\��-~�Y]1-x��s�#�uz4<�a*�t|��a�dG��:5�ە!��=�~*�_�\:2G�{S2���O�Y��/s;X�m�3�&��`{a�C�AIx�m��V����V}5C�	g�ﶓ���^`5�N[/�([綇�/��z�S]_�-�.��4��p E��v͂ż�c'�jz�s�k+g|!%	p����&����ïzS��lE(�3��
U|��'�)!���I1١��0� �0k��Y$�6~�X"�l��^�(�<S�d�ݸs�g�!�Q�t+SOnB�OU��i�(�E�UڶM��ߋKB�8zE�K%��vu)������5_�|vTT1��q	�8^���7��rc��{M[�/��U�p^�����+4T���V|U�"wB]rN�%���X~�A��0סl�ʻ�*��$�{�o��z��g�f�x�s�B���׽����B#��\�L����|[[�CV8�a)���<���g�Į�T�	�O�j�^o��D��z���K�&��ח.4�CP��N��bVD��sM.�L{#�)i<%� η���C�Yl������}��)��0�5֘Lwlu�,��Ho(%5��O��e!!/+�~  hX�/�ە	]9��gY��S�(9��ڵmΉ���n����U͡�w\{�1��� ?�E�|��q�ĊV4'-̟#� � )ي��?Ļӈ5��t��!�%�/<F�>p�s���c�*�Á+��{��kd�L|/�9w�>��v�����V�ܩ`c.�P��J���,~�%k�d/*r�NnQcj+;�����l��R�x���)�fht4��'���.��a.e�J�xX�R�j�(�H;@�y �,��Bž�qD�DW1.C"i8ٗ��V� {P.��a��I[�F[�'�e*_$��V�����u�%�����:#Ī=@%��/