��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O� ` ��h�܂$@�{�>�*�[ӻ-����s�|@�z9�W��`���S�4���ն|��p���v�xm��W!�N�c!O�X̟��R��b�d���P0k��R��Q��\
�K~���VV�[�pZ���.��������I�$�y[�bEaK������C�Ћ*�}I��eKp���^jL	2A?p\���3�p]�qà�M���T����Z������S���,2�Pv�IMi��'`�x]�����;T�m�p�*x�:���'��x5/�U�+����c�����F�zkP��Fj=�;/��d9�a�Fdsd��dg�"�w=�m�b����i���7֓B뙶F�D((���� 7j#�f9�:Ӣ��dW,ë:��GB��>+<��t%��cO��(o�k퇡�j�[�]yI�=/�y�O��9��C{M�ѫ���\��\(�(�y�ez����a.f-���	0�0�gs&��!��b�C�h$��E���<����:�-0tvW������e2�T(�w���"�H̎�����#C�� Y���9��Ģ]�6m���k;�a?�\�wߡ�I�f�pذ�~����X�N��F?z���{z����XF�����b-1�� f�,��K����	������pJWCC����Y�!)�&�!=�V�������I�NB�;'	�mg��H(t
G؏��-`���3a�E{�.���}w1���>eĘ�L{����-���{��_')3=i����Ep�x��� ��T�,v�jaŕt9m�ѷ}�LyR�����9��-s�A�W����!zr~o�f�y3�	BI���K]:&�r�E�f���q����H�A��j��`�_&L����E�
M�,����+P��hRG���=T�\L��Yc���e#g?����.�И���5�7�ٸ�G��/��}����|Q�2JYc������Sm$N��Q�����YEE>�̽�Ĝb@̭fJ1�(�%##J4ec�K累�z��ET���R�I�l2F��I)p�%+�&�<�=(U��.�!��ʕ&�'�{������S��<�c�7��d�����U�3/(����J׷��r�hp6��w�[�hHz�SW�}�=��^MC���X_�N�D$�����͋��{��Ɵ:]3�ҿ6�W��n�C���;l׌v�׼�(=	�3��"NMӋ����%�Z��
9b��mo���L��F�r1�_�r��;^>Fخ8�R�($�>*-`v������c|���(�2G�e��BM�jks�'��U�'��}�.��s+ߛ\�6]6�: ���~L�;�Nol�#�jhkѣ�,+�:E؀W�5G�y@�#V���������vWy�9�0�j"�_�g���?]퓣�+�{�ݢ�ی�dW?Ԫ���l�2�4�&~�HM>�Yr�.������,����~l�d:�1�J.x��#E~m��v