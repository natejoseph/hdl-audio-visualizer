��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C��Oҷ�$�S�u��B=R0R�E����X{W�yh�)Y���ȷ[��Y94Z�|�cLP��!��U��se��\���?��C���k �:5\�,��I��l��:H���C����#RH�t"�qͿ�ǆJ���F�J��↫���������_��g0��?�/w��Y�?'�R���ئ�m�T��jmdK7O�0���\?�m5&ě�	��];��v*m_�#Z�M�{��f��ٜ��ʬ �&�5(�^=�V����kf�|Y��H��Lz�w��kD�4����4P_����ΐ�l�cS���x�W�pl���[��n9�{�dUp�2�߭b���G�~���A��?c�i!T�4Zd�$��'���.�v��g�y琳���9{i?�-[g����/V��M�=6=��Jc�&����%�)���Y�a�i`[��ȋ�R��a��O�a�߶I���}�_�6�� +IT�)��74��:��@�l��j�V�%�~0N���3ߛ�2ޖu\�KOj0����xO�I:��93q�5(�PS��lzNXJY��ϓ1մ�f\u�>V�/�)���vڄ�����3d�+��d�E��Ӫ�^+pQN�!`���b��8������[���a,+�����0�r$&Hr�g*Q�Af��7��zR���7�J#%f���E1�����-i)�'����S�I����jW�ȹk+�����7v��Kb�Ecޟ3�'����ZX��r(c�e-��
�&���zŧ����`��B���g��ϟ]�Ec8?�xd��=f�!"su�_3g�Ė�ٳ�u�ɉA���"��-M�{�Hz?L;�{�L��)`�[��ݰ��<����]Č``��1�]Ku�����Φ��29�1�z������uf$Pv�2��~�(߇�h�:�ש�J\��:����:�'
Ӿ�h�B5���	4�o?�q�W2�kwA��=n&� �ofY,�h�:TM�+�+�39 �M��]Ģ觿 �{r�O�O��a��Z2Ҹj�vV�<Cz@��N��m0l���c`A�6�PH�	2�;�w��Ha2�1�֫�!��5`�ӈt�:U�p��p3�f�	c�0�2�js(�����TQ�l(@�̠cq'Xd7�-��i��Wm�w��-l��Z��v�r��ӯ��a^G�m�b
�
s7��*w�j�a�8b�!���b��P�3.q��VR�/]�U���.1A&�ҫ%yhAo���~cI�VOc)�| 9VNY��ŜK�%���A��E*�z��y���ӴD�Wy؃�l-|���
⃆(�r�D:�//��:�I���_a���ٱ�wU*�&�ې��EK����xA 麢�/�Y�t��3�I�ԦWg��ϫ,�z}%��[I��V�*�HyM+v,�L]�� ��X����p���A��@�J���Q�9Z^�gB�ޒ5����&���b����f��4���*����?u �-?r�N���?�_������g��w�]�\ j�y�O9o��Ɯ��N�M�MNbw4�<��e�|��Krc#wn��q'���0� `˧lك�?��A�I����
/��f5�x#���El���mt%�x��|�F���O�D�(���>*��Z���l�����M�'�φ�3Y p}&)f$� �|����������F�"����;�z�P��4�W��C���0]%b�U.8���58-:a`�]f��r>����S&���^�gɀ3�%���vR��	Y&��R���:X\Ul���b.��}�M����p��b�;�'M���ء� �!#���,�����&9=m��$�����>j���U��9�!�J���X��[�J=�}�&`H\��7Bi�7�]+EUZ�9���/m������y���^r��8[.����`6{A+�����%S��=1,�9qG=�_ze���9��-�9���?�-�<�y���c ڂ$9(D�ZIp�����<���gk\
�^���4o�n�����mc�vA=2�>c����Y�%��䢕M��ȓ�P"�$'H�F����x�#*�K��TRn����~<��F�<���U"�@&Q��:n).�Óq��ǧ3��z��]Eo�+t ;�[�
�֓{E�����p��s�j�"v|�V�i�H�|��:���;K0���<������h�cY'��-u6��9w¶WyӁU��}P^U�����#d�$h$�Ȳ�BS��/�%-FŬ��%9��[��xPq� �<;qkU���6��CR��ԱO�����������T��Ev����8	~�����氇o�oJ��Qѱ��g��|�s��x�eI� �]J�i�+�!t�`���' ��v_�+�6�g̒��Q>� �����Է�r@ׄ���^\�u�M�0ZW�;��_]]����a,x��|�$�̩:��e!��	�mi�TV�q�߃j�e�h�%*��)h�V�����8O��khShϦ�o��N���W���oD/������0�0�+_LJ�c<��g��>��L�4����Q�#�2��9s_�ke|L�'�!+ O>E
/�!#�$�R�l�+�5	_��:�$,���Hwa�9+Y��v�PjN�����Z3�Z����㙡������Z	70�L�*��N�1H��lC�FE�C�ov+II����]-'��~���j��O���D�\��>EƳhq� B��t�X���G��b�W9uJ@D�"h#�@���{o1������z�H"��r��&j�wvy"����YS��s��*¬j��!�o�7�{���T)
���I.�Եޟ p׃hj �l#p�����*��=���ne˒9|��+��[a_W��	�eF��2��I�l��Bl��dT�s�����e�t[�k!���jQ��CTF�(��+�ƹJ��J,ᾝe��zޏX,F(�䭢���b��)��7���ց�O������ j��8�aS�b3�%���q]a���8R|z:���^�#H��YǄ��NR������x��
�A�t��T�W�@��Dx���L��ND.���e��/$�"�Q�CW�3lU�s����0�Ւ]F2�$[@�D���OԱ���uce�/�E�̀��2��#���d�|�����;{����L����j�g�FAX�I�	=1I"��:��@@������T�i���M4�\��q�N콏�q�2%��U6��h��Ta����q7�Ũ��!�W�%+�d���(���H�sS!H���/|5�Q�=o�����/�mQ޹'��<�"��;9�EF�F��\յ��+9gQUܟ��	J�� ·��±b[1XH=W�\�߆��뤭�A\!�%ыe�r���L��	�Wʂ��׻6�倆�n�_����Y����U��tw��~�5�@�z)?��W�#��-��	��Ҙ�W��3��;��{UP��F��Jm�ƍ��/hvE�BEpSƊ�L���₱5�B����v{�C�"�B���3��o m�w3����Y�cxҎ~���T]�5��p	�*@	�a �ۛA�GG���$5�$5��f�b��	���+vx�PT��.��Q���'�D�ϝ���UX�;�(-�aO���ۭ{�bnM�a�(Y����^[�ƾӂS'h.�7N��`��׌�����Ƃ�	�Bڭ�}/��.�[o�甒�9�����#x�����v�� �/0��p�EfTp;Ea�R*�t��ht�%�e���#p�0O���Mm�[Y.�?̧��F(�������Y���^�����GԄ1��+U����<�Tx�����{%m,��c�}���K��Ru�q`�=g� �m'�o�����43���ժ {Eտ��i����|M{���� ь��l9���v�afM���j�}G��y�1��pl�L�x<]Ǌ�JG]L���T��H��2�2+���������R�z�7���.-�$����|�)�)�R#c��G����5����sS�|Y����X���n��2F	[2��u��G�y�F;�p��@�-k�}崔����B�tc�oTP�N�������Ws��]��
��	mP��\"�S]Ph�:�1�*~bE�巋J`��t`�_�B<_(����WA������@3��o=���D��L,��ٶ�����\�	s�@�ѼeߕB����@�[�Ց��
K�6���gm�J].`!��C�_�fu�r��`��2,h�q!��S�0��v��|�d��mQH��4�w�̂��g�i���g��
�c�mb��ڋ�����Ks���I �}�$B���w��P��{\2(=i���[�ѭ$�f���&j�ztT�mD��Ϻ��&XGEM9�䊿�l^���	a� �����2h��?3����-�@OYڮP�&�'6�0���Go'u)<G�����Jyu�ei+�*�b?;�Ow1S��_y���TH�SMjx�����F��)����s��V��~��<Xl�%k�Qm��.����W�M�m�&B��2�|\J�@���EqkB�X���+$9� KO���H����5(M�u�~�/*�M�������S݃!�ĉb8��K�2/
�֪̗Qb����S�?����F�\�
"��\���L��-�)���/�%9��L�b��j��##���U�O���?U,������0�C^V�v�5P_JM�;xqұ)Y����}n�VM&���uǣk@y�L�E1N����5҆����>o��Hu�_�	�04!�6Ğ���z�Y4�	���9
�������m�$�,�i�S>�(��?��4�_�zO�o<�`9���o�^s�������3�f ��Gv��z�o@Wk�~�k������F�k>��e3@����DP�ru��0�&0��޼@� _6|Q�Am�h�b�����=�sk>����h�P��СE��(�zg�h�!�Ook'*��Yϝ\~�I��|U��nA��A��C�2ߏ�c��H|݆�����,0���IK�iA���,:7X��\A�u8�R���!��bbR�T|d�*:��������sMn5?���^b!�������N����J��v�#�	�}l86۝��@jק<1S�N6�P��r��N&���9��_
�({{ƼM��7�r	��I�3��9����@�ց�[�㑣����\�r�l���y�-5�l9�ԣ%�Qv���a>��3��"AT�ɇx:�Q��w���[!�&���h����$_J3u�*?�Ҍւ�,�~e;�0i�j!gwC��:����`�Sc���;)H?>�ZA�gV�i~:�(%8�|B���(Y��M)=�K��R�'*������"�"&�|$�R�1���r�� ����>�����
�+E!n��i�S;�*d!A%�3xe�/�"����*E0 �Y��/�����O��!�BE�h�~j�oDM	/�<P�U�f�8e �!>-y��!I_�����+��+�+����������Ē�i#tϻ �`����&R���z�R>�i� "��/�*X�H�k1wǺ�H��bɦ���k}����wAR���c���2�ޥ���s��o�_�ܕ���0{{��@|}�7��K���S2�J4_m�ư�{�mtDq�hN�a��
��}?���/t��9�O��� 8�plٰ�;�8�BI���$nG#Z���<%=�Pڷ�axG0�7?�d��ZL%�2�sT�N�\�����~�P[�E����z V�x��)���0UU8��9@� ���1K�V($֟��0`C�sPf8bu1c�[�L�}�1�#Ca��Ý���/�t��Ax�3D��F*�V��(�*��x!��{f9�a}髰d�2(���J�,��)�i�m?��\�1�7c�3��O�u���H<3��&G6�����~\���[��0+:��l���}`�j�� �UQ2[o���m���}�w_���;7��]lK�f��ɝ��
,�|O
x{W���P(ۋ��$��	G�:!�@�#���r�rj�J|N�'����	eP�:�x-^��Eǝ[�>qJ�	���)
`�?�[��#����ܳ�^�w�0��{������~_h(�H�/��I��?yA�V-��Y+>BP�m>i�Lf2ܫX������dTT5��������n�z,�V³h�.mq���L�l �"�̑��L�)��׼��n9P'�9�^�����R�g�]=8��Kvbկ��k��pZ���A6@��{R\zE��� p�r�V`��}�_bGC�Z�f�4��d�Xy�?���#'ΐ�]��/��̧�⽶=�k�e}��o��G�5�$��W��*��8@t�F_�Z�8}ȡ����;��iM&ͣ�1��KS�uA����װ�N�+>
�x�n)}�H����^�=��F�nB����IL)*�� ��a�O)�蓺2��ْ�f^��Ϩ�N�������9��+��0�5�����c�R�g�HR��/���e�o�t��6)�}��Q)�EdX���-������묘B_�9
	�3�mLV�{�R�iW�:�V�F��*�p=ǑT��f�\<هz�=m�H�nZ��������m����I/\L��ض�A��Nau`t��QFE�d�����¬"Y-홺c�pJ��u�����7��qI&��􄝦K�v�iay�E&�lؚ��}�A۫=-�o���9���h���ղ�q[Æe�VP��7��e�7EB�t�6|p������R�phrk�n�w�a
zɕ�Z�։:r^_�lZfu�e���3G�����9� ��W��V{Q�@�|c�Y�!Q��E/x!���~f{�m%�t�_�w���B� �4�Ih�3���E6�H�f�z
��~��\"PO�Q(�LD��Y����t�/{�GX��H���`kȗcS����2g���Q��E���&�2�#�����- ,F��r��Ϯ ��_|�[��8G�y���˾!�Y?*�d�1?�+g�qf�?��F�P{��nľ�������,PW��V�����UV痑N�*���t�$wQ�H��S��m𳾵B�Hƛ.�3t���y)Vś������] G����~�ވlW��[na�����8j�/s3d��No1e��k���)��jl�.@�U��ņi�Ȳ�F�:��{,�u���Zw�Je�Ŗ*���De-R��E`�yu�ʄ7�b���& z��~ ���W�U�;����T1�D3��C�L�?/[�\��-Ҕl�w�{�Y4���3�WP}���U����1��� k|9,~O���@Kp�8z����M�� �P��p"��@�Ӣ6pRn�0���*��to�L����]�ZZ�Oo�����ݪ�G�ǩ��R�uMDv6�StA�2��z�ܿ!n(�Ն���k��:�����e ��9j�	��/�\����*p�F��$C�26�I+f-�]�<��(9IY�}1�K��ˤ{�І��nv�R�%�x�U��O��H6��x���=�,�9CG�n�8�]M&�\�Ί1&8,�I72� �����!*��Ϡ��<6Q:2�����<�yN�/6
�GwP� ֿd| �_;��]n�#�5�׵A�?�sl���*s�*1y���!I�B^�T(嚰a#�7GY��>��T�.�ӟ��\�w5����Y�����Q�K��
	��ٜ*�	�6� x	��e;�!�0\��'E����Lt����l8�$Z�1Gcv���Au�L����;$��y/���Z�,��-�X�UWo)J;?>����b�Ĥ��c��S�[�"5n��_���&T+�Z:�����iv��%^m�5jx�~d1Q�K�-	c���~��Iג��cVGr�e�
y�0��Y:uC�LeA��ɒip�<y�%����݋p<$O��L{x�gkàt4F��������m�rAqm̩��	Qs|�~��YA����i	6r��._�,.`�$.4OD,��'��kBg���Ū���~��Vǎm�J�[���U8�}JyA+䖗F'c���S���pR�����rԷ\!��Z<E�/)AaE%v�f��T]�g���0���ә5e�J%���kد�S̮�Y��||�� r#+�@��F�����#&Iܷ���`k}��Y��T*[�+� #7O�,4i1�{N�-����:n�}A	-Oc�������oW ��E�F��$4X�n�	��7DH�1���S��[����LZ��oe5�Ox.�t��M4�;�^���r�7ɡ6|�����L�O������
����T�L���#��	�1 �\T�?#���2��P�)��#���N���A�ʴ�� �&��лY˱���u�F��{�^Vx	U�SrJZ���>����fQ��3�rx*T�k�ȧ��������蟼���^�B���W[�����vZky�J���9^�/|�2_��L�7����ЉH�Cf5�t.�R�Z�ᜡ�=��)gM��tؓ'1W�|�/4՛E���-����<J[����.,�(�=H�_���p|�fP�1c�f)iB�N&rO�¿}���ݼ<�� �4@�<�[p��=?�QR*��ltg����OF�0󙥳X�j��@-�]x��S�}��0b�ڞ�+�����~#�;��u��1�Rn<���� ��m�pL�E�.������tlS��CD!�xZ'�n������b������@����M q[$���ڃ��
�W�V��6f��oم�z,I���r�vw
�pO�N�O�f��<�*O�\�"4�����F��ߒ(͒���&����+ܲDy�G�m"��61�6��V�ĵ���k�_��,W �~|Qol�W_j�
����P���`�(�r5��_����h������ԮV��ج���T�텂dI��ЈK����d�R�K*��+��Y�HK��{30�>�N����;x֮�U�����͓����*�8��n��G-�z84F�����w�TLm�p��D�M�@�+�o�3z:j��9��7���\0������i���@�
/�#Q�k��D^��3�DىUY29�lu�ܦEZ;��~��zpħ�;N��]��AqN�o � ��k�r*��ctR�.:�T�R6��%�Y�����f�X��D౫�q�_��L���c�e�ড়��@y����Qop]��k6>{�n�>KF]�V��u��z�&u����NDֲ��ͽ���?��z�+&�T���W��>�q
���>�� F�R������83+���fǯF7�,&��x��&ut^FY.�`��ʳ3e_�������֙��k�95�0b	'��,r(��~.�7�v�	����^���2�zsh��w�G{L,�-E��S�||��1��E�e������A���|~nB�V�^	�v�cx.�r�~�T�⽌i�C̹��A�(�9���n�(e�bj��1W�Ƕ-aH�:�+/�=�u��_�DU� tF"}8 >�ъ�L�Jl(�p��I۱��CO�V{���e����k 6F��n ��Yx��\]u�!W��I-�̤���y�B8d�B�B�	��_��p`�iK�Q� N�Ĵg��T���df�Ƣ���\�*_ڣ4�������J;�&��W�� b�=>]t�#<�@	aP/�
�S��%�:)�|:���
�4K���W���b�94�1��[	D�5���J#]��è�1|��e�Jwݒ�6�W�֜�ip�<BSգ^��?|;��8b�=���M��� �T
EeL`����ȟ����A��n�Y��x?�&,_��>�3���Ih���A I��ڡ�� |�]+(���Pt�rPj0���ݫjU�.
��Z�Ml%^X�Ā�s���#^a4�Ye&�����k�]��c��9���*�����1�{N����j�"̛OE�ߺH���� ������N$��B�G��t쯏�����ӆ�����P�Z��vpNC��]5Y��b�~��G��<�[a�CQ�n��7�@��8o둂��0��U��Т����Mue�ϟ�mC�yv�D���)�^��OssE0�n8�7����^Y��j��,�����צ���G�v#!^0��օ��(���&6�[�Ĕׯ�sy���Y%���ҲBU{�>ψ�I*�ѳ�������n�hȘ�
'G�9}7���/���aM0	��~�Z�]��/T3�l��S1�L�����d�O�X3S��� 4���}K�|�P谙�p~r<�36������5���r�%;8��o�2�+v����@��-3��ٝ��y���یԟ�:���u�2X���Gy\Y2��#�k�q��8�ϭRg��5���e��$��&,%�K&�H�vL~d����B��Up�c.�Kk.Xx	�Ki)�Z�YX۶�ۃ.�ӆ0チN��lO?QG*���̢>�S-��|��<�����!k�d��\vF�m��u���v�r��}�ɾ��X�Φ�B�Q1�|�:�L':��j����+��u�������ZQk�s���������]����Z��^'�/�Y�a��
;q�{�՛��W7u������N�:G��m;n�%D!k��5�l*��6��q�#����)��8��15���"o#���h�k#���y?�����\����`�����Tr�բ3�_���?\�+�T6n���/��Vh�_��I��*�˰�_��+�ղ�8p���W,��!4��D��]�p�r��OR)T�fW�P�|:C��|lQ�X4�Ǽ�`��>�Y�"���e����E$�3�S���<��/�<r���V�F��`��p[���Iq3�5^A�Mٵ���O�^$�`s(��b1oT�S$����hb!Bv��1S��f��$^�����?�/��`����5ѻ3�Z�;��)���k���b���+_;�����!��],N����s_tVP^�qIWi�g=;��)���yyk�I�H7���K6���\nF;btz�Yy�F�?�����iD�,����CޛMe���O}���	un0���n���SՁ�mܒ7����MJ���Q}y�s��\�Bv�°ZMx��aq�_īy%�l�L�Q�pǫ|��hd�ƶ��.�5_ިrD�����Z�������,&@��@�u�4���ۮ^�Ҹf�#ek�wb��Ε�=GI�r*&��򿺁vF��,�UɊ$bL)���A7{O�vBK��ٺ������p	l��;��e�C/�k7àE����ٙ59�U:
��w��g̞�,�h�"�4G9����̰;MO;�`���(B�X�G9;~YDw}��\R���_M��`Z��8#,6�����I�Y��%���40m�t��CeL�?�kJ�b�Ƴ��� 1��q�i[�m�	?�c,5��t�
ߑ���s~� %E��)�٥>%�\�YW��y-�Ց�����n��V ��M�ꂃ+�=�Z��M����%3��?�ͼ�gXga�+���VI��Z�W�04�Y8:!3o�q�V�ӛ}	�n��,"���O�#Ȓ~�yg���
,^�.m�.����MP5��#�*�y��^�3?D���=�X_:=�ժkt�.��(��6�*���n�$S��|��C�B���Q6@l���!��!ͷ�.�0��d��H���m,�2z!��z^�;������4��+N^�`��|��}i?Ż1bE���iq��|���|A}�#���=��G��y�)�'���� �3	��m��蠨�f��Lq�7��� �-뫆'�ܑ����k�