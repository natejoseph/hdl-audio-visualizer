��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��N(��)�A\k#B�L/�:V�J�P��}t��L ��
3����J0�+g�2{�1����1�&\�Յ�AB6�z����L�bR����C>fc�ͅˠ��QO�c��Y���<��c$�[gw�c�| ��J��)�6aߒ
:tw�z-Ԩ��x���Y舵e��\a#�ʶݫ�������IT# �aK��U��l`�����\�3�gN���!���7�Äb��A�%dU������x������;tm���|���	�ޤ�܍�aI�Y������Zߣނ�f/�c����z����C\�r]��&�H�Hљ^_�$������*�04/y�A�2b�����j�(͕(���v[�ɭ��y" 3�D��/#��77\������� �����h���e��wϱUg!���o�d�v��P��t[܂�ٮ�beK�QX֠���s��hq���?l%R�60�`ⱱ����27�M��U��a$��0�P�T�'iv�FpoM^�@�Q,5�g�&��M ��+ZY��Q����E9�r� -S0�w��.�ױ��,M&�9��3i|t������	o�@���h��e�%� �y��}xh)��T)��l���uً�ߥ>�6��
Ʃ�)�\�BY$U"�Z2��y6�[��c��3������s7��C*#R��9�����@g-�|��ނ�)EJHt���^���⌼�e��Bt�r�t�dӽB�0�����z	�d�=��:wR7,os9��9�8�*|��F����*���\bqB�������4���"Nk�,��uXn�y�|���-)*,KRz/-�\�Uǻ���)r�	CMX��`l*����jY�����yŕ���U�Pb�o�� �Ў �V\շT�7̈�&�o�;�A��K�^��]�,��V��J,� Ğ�.��.�-~:CY�+�c��"���J��� �l��wΡ�Vc�ES\:�ob5Bsz ?vc�,7`��;��m�����wc����b&���%Sq���Օ(��?�(r����c�"��ڭ����ƽ�Hm��b�6�Qưhȏ;Y�&z�����G��\F�r��
̆�����n:�kqg�{�H��7�'Ȓv`_�ƺ�V�]b�'Q�ө�%�׼_E0"}S#T���gG�)b-\�2?�g���k#�,�DӤCp��Uu �9M�t�%;^x0}[#ֺ�H�����F���}�SKG���z�h)�dح��:27\�k�4BQ���⎙����(������<�@���%q�8�x{��Ͼ��w�h��N��j4f���=�0�,n5к�
�d�M�Θ#���#��d�H75���9�Ru�%�`$��"�yX��e@4VE�w������c�2��I�(}�.�@�bZ��5	�M��S�>)e�L��J�6=�ʠ�ɛ{�Լ�-�m�e�!��u��FE��ٹ�p����Z%1�����h���ߐق#�B�[��$W��bB�E�Q�בI����[��j��}�]J3ג��{8i��SM@��+;q�#��	I�Rr�Ƣ��5=�d��k����D �5o5�%�ȗ-d�`)�<�C~E�<a��w�\$ՠ#�BR��O�"�I�Y[=��?Ca=��<�ya=샥r4~4E��V�ڏ�\G��Nk�7�R|��&�N"���|����M�)� @K�������ˎ�pm^r�P��Z�	�L6�r*�m��qɾ���F�@�E�c:A�PY(a8e��'��o&�Zĝu��>ӷ�QG�[h��?�gC�h�����əǄӓ��#8ޑ�IDZ��H6��ě/�$�ڈ�Rh	Y����YY�ͯ�L�˪y"���oJ��G��<�W��[e~K����|�3�r�y3�%���˰��MC����>L�����FA��-T��|+U�S�R?z��7BL�]}�CG�`��|))�ߧw�*��;o�JIo���d���Â^���p�*T\�׭�y+�V�Թ[�my,�ȹ����8�;�2����}p�ļ_�t|�A"�2bb?�t:��r�Z��&]�rMX�'1���N��|�6�UO(���ӧE�Y1fGXO���DZ�K���ly��q^����j��J�s^����'];�e$�%�Ýح�;[q���h�$F�>�(�a2�J�RWWg� <�>2��,�"_�����%��Z]CJ�ռ�3�7��A7}JGzr��b����>پj��n��(��J����[
���V%�h��?{�'~�H������&!r�+e{���'|7�ׇ�-A�0��xe���Ӿހ����k
�r33�H;��������f��F�]�����/�b+�c���+�/ l�Y��զ���}�֛�w[�g�h�3w��Ȩ�+�bu����\����e�{;�����n��3�F�4kl�D~�oS�r*u& ����=���U��â���ȏ����:�[�?TI�`���_���[]�t�^ ��-�3�d6��[������b����fA���e�#��=�'N[\�2j�:�j����Jd�$h/vԌ�c|?_R�+8Z-�6���utE
S|��K�5�$�˝���p�)��$��w���]]�sQ��l��FB�tj%�W�x���������Պ��]`����M�m�=d�E��qE+P���;K��<I-GHz�)Բ+p�j�wܓv�B�ȋ�c���$zu>����v��uA�J�b��5S�sC���&j�����b�~��ߨ���]�v,����S��Y���M��b�:�7���=�m �F��+7�b&��*�|)�b*�b+z.��7��a/��+�F����'�f�YRkA���ū�<�y�^��@���
2���IO�O��!d.BX��'���鰀I��> ����[�^��h8�����s�W���qJ�@Únmd�,ދ0�Iٶ�W�Wy�+���>v�xd���,L*�WWe|��~�d�ף��S��*��A�W��)������M�&�G��
K6]>E� /�S@8�nV��n����Eh�bZ9�E���]�6T?�U2VE/n"c$�@�j^�8mX�q-}�Ժ���+����Q�DN���g�"����Qu�@��F`�Hc��=�Q.������CK�p��L1���n-?)Ƕ&��\�ч�6�n�R0ʀK�2ޠÑ�!]���f��Y؏r��r{�s�sj�Q��EN�]h�=o���57<4�*��H�	�L�݁*ZU��HsDL� ��L9�G�9�W��-n`[�ao3,�ތ��h���ڿ���5�C	�����
��<���*C�x�|�i��x$�?jN/G���rr��܁�,_@OG:�.�O8�	x.J�'M3[U�s�쨇�9�YMML�l��SDaB\�fj����ݤ���ME���5T&'��W}1�ѳ�Cʒll�݈�ރ[�R$�d���V��To7�ACȧ�i�Ӥq�UJ%�`����f����M���4��!}����q�P�U��`�=u��J��]���Hx:�V��_���䉮0�V���Ck���ߗ�M��"�. ��Zr8-9��"���򊴼��&,Gc~���Ę���,���%��A�M_��[�HaQ����FǗ����tz�?K?b�5K�B��$�Ir�SqΓ����y�qx ����!&���O�q�?��,�������
�+����bA�RJ�����y��Ο\V��LF4�
����:	m����-�1'2�+�:�?֐]
��OD	c�G�`���=��/�G���'Q?�-j�3R[$9�~ޫ�{$��3a �42��i��c����Ȧ=�T�pF�R:�ty+��butBL�tՑq�]�ue|;T�y�kĈ�E�ָͶt�:g�1L)�AĞE	���c-�zF}ba
�"���?,��`w���?F��5��b��&K����x��l,|��|J�=]��wI��j&��K2�[* �����w��Z �������n���1���N��I~c�����B�ALl$��Ƈ�V�T sv��e��+X�Ϻ��ry��X��wx�t�v��q�}���u��J���'��ci�.֔5��$AQ�1���Ք��3�C���� ȼ&b�������;~P�)u��	ǣ~���;L%��� �s*k�sd Gi���;�~p�0�V��{`<�2�\��R���"V�����[X�'c��U{n���*_�ƾ��oM��`+S�쓟l5,��.I�qV�
�7a��P�y�)�&�(�7ؠ�|V\�8'�ҵ���ܜ���/��Ix$TB^>5Z�'m>���uW�Ɗt�,A�C�>+�|+i.��M��Ц��d�X����Ye�9�E����l�ӄwC��P��g���E��9�'�A�^��p�:&.��p�}���2��Z�Y��(M���\�qv�K5+ƕ92�O�K�TS�{�fM/��1ai�pyOi��U��+����F$)Kc�7a����YUC����΅�|`��%��Y ��+��7�����>�Ah�9\Y�陕����7�k���ˮ#�W�|VL��=�:�%b�Myķ�m�6-�3�ل�<g��:�hːO��J�Ȉ��b�x9�k��S���[6u����:rm�hd��N_�L��[�x�Yk���|�%�I9O�Z����1�M�K�F�XB��%t�T)�W�P7��
�R��I-��s��S#�Zf�V�gލZVe��x�Nf��㫡|a0���dy_kc�a�����_���I�8y���=�y��M�=��Z�$B�{��M�����͎���\'[��o�W�Uza
,50�����+�s�b� 	��d�2�*�?�
�zq��)��M芒�:���Y�\P���~캅!L�&Fo�3��{k���XՓc�VB�{w��pU��v6oΖ�OT~��i^o��?�aD��\
G���56��&o���s�k�Ǐc̘�l����;���po�������4W��h�\���(A�&
u0ft�-f���͓5,`��>�2�~>[��v��*��R%�����iqj??�������Br��k�#|����5��bl��`���8*0xE=� ɛ����P������J�����H�(��,������'�M�� �%ZY�%����ǧ�Ϳ�(���*�(�8D֪#	&2w��4_W�*¦���'�#�{
WqW>��Cog�f�+>W,��FV�kAV��:)��L�\�>ւ�u�1Wrz֜��բ!�'�������.]Ι�-��-�B�W#�*�i9f���[-��n�U"r[���՞*%2 �@�e��߬|�f�{�$=��^�N���ݻr	����b+����F����Cb���-/L�/���:х��U$P8T��'V����X�.�?�BI�q	�K�4%�L�1ŗ��}����9�Ѧy����C�;���un�k��m'H'Q狮
��*Ska?klEW�D0�hU��Nt���!#�2R/�����GO��*��L�-�Y|��0����W.�N�����p����W��~Ц��tq�`m��7_���}ORN�v��ռ,,�����~����2�둢�iNWP!�e��AwbM�05���<��?Q����^�ɝ�/6��L����w�`|�|�������!��ns����ˎ�"�z�ZH�8��$x�4¶�=��>[̟���m�޲�YB���Q�8cё���Bθ]�}����Ǖ�M�؅=�q���{�"�v6JE���6�|�Q����?VI����M���@��9aT�/$"i���8�}tܬ_1޳&�j�	��A�;��#*��8�V�멄��Wh�X^]DI�3ݨ����#�I�)B)��|������86�'Q���$Z�$W�6�S�=X��! �#g����4��`'(vЧ��}�uRϩWa�|�Ĥ�Y�mʎ{N�r�U�Ϻ��y]���O��ޞ?��a£x{�N�뽆Y�@�?�\w4[emO�5��|��y�r���#��!:���)y4���=jl��^�7#��@�w�m}_��}��+?��K�Y����\�#��XS��t
�n4jU��yا��]���\�&��5s�;�̅ ���\E/1��j�<\�5�+��>5����b�yI�aT�g�F-f�q0�s �Z��첶 �-�Pb����S!�ʳ�j�8%f���oٞ4��Y�"sH$�����n$�[rp1�6�����e�(\Ln��������z��l-��uT:Q�~!J2y�EK!��~����^iɡ��.�!?��txy�l�����;���{
�rQ��wc�.�%�OK��8p5�̍D����+@$D�zR�
fm;x23�'ϊD����:��;Q�"���9���u���7J�cs6����T�P�/aC{�ILA��0~��~v�ͱ�EoX�L�"�+Hp`�=�F6��{4s��t��41�M[-��N��@�\R�A��6��]P/y[�7����E!kǣ��Ӱk�h��<�|�E�t�Ƥҫ��>�S����Yb�p�s囇��>9ɥ�zw?����#�V�/�Rvw�����i��H����Zη��&�( ys`d�2faV)=&���\X�f%ѷ0$�%�� ������-�ia1+,� ���&$f�XW�c�^Ͽ�U�i@�"����ig^�i�i����\z��2��Df���y�u��L��C��T w��9d���n �����=U�ro��ݺ��-���:fuJ�pެܹUn]��&9�.jřL�I���]���(G���u!�n4�����M7�'����QEO���7��$��w�l�e]��w�X��bW�E;?�����瀒G���c��N�.�zq�C�3X/�S�� ���z�aX�����6$~�ɕ����/��ʷ�����)��P�TN	��ȣ�����5]��XN���!����@r�_�R�@��ˋ����
��۝�� �?��2�&�!;i�=��df��q��jOs!y������Z��S�%-�Si)|i��e���;� Ok5�^H/O�}z�P��[�q�%((������b�y�'���,��/���1�_� �r3�\�������;��o}�h_]	(�0��g�����ڻL�v)����ع����N<�ͱ�
��B��E3�M���o��QH��9KJ,��t���C� 8�{�ߦ���d;p�À�[˗�L����T7�T/IM���̤m1C��ܩ�a���*��p��:��%s���<����SBˠ종"!��^�Z�	>� ��?<�P�Hάj1À$
�J�]�1�N������@�8� ��?w��mU P�L^)�v��Л��B�����%F�߿	�$�5ꓬ�ث(��I� ���h��&���eӫ1��w�;dzr�{	mJ?�ӆِ�~��c� K(�-/�6���[c^�+ܮ�cm�s� :pC�s��I�m�	$jg�����eD�s�@��Jt1��kl�Ҁy��<�0�?}�(�§�	��:Ti:*�m�Z��uںy ��p��~�����z�L��`������=�zp��O���(F	@V��8��d?Ugy}u;9�ȟ�ɏ��i,&ƕp`ج��wkrt�XIR�]]p���J�g��'lxnԇ�hc�h^d<z���Wȶ[? �g/��
�>����# ���[~���Qs�wD1ִ�'�Y�L��c� .:gH�X���~ܓ:�	�L-{U���}~k�a�@����|ZCR(�ewf�^u� I~S�`���v�,�C\�E�,����Ɖ��o7:ɋ���$�a��Gc�y�:`n5�����a_�	0��3�Q%�ZԌ�n�2��-R�.��[_�k ڍ(��}Q�i=�B��<����[��գ�*��<P8�:kj6ѓ��'8���A�N����sxU�l�@��xyQ8Fw�2��皪lɛ���o����U~w<��b�߯�|�K,/iܐ����ױ�I���ebFv���Nn݅�h�� :��8��ajk���j<�!�%�� ��漀�tV��Sb��LЦ�e`>�?U�U��8�'��oR�''�uJ�ɻ���֦�ᆂ���8͒���1�Y_�n��Α��u B�!�ݐ]�k|=��z�S<;I�n�-x%��w���?/(�52%HB��6VB�/*YѾ��(Ũ�P!�$�$��
�s����)gY�x�W'�
�Th5Qf|/����Z�k&A���>��ּ�N�A�	�sZՄWܱk�?�
��S�$E���skx]6� 37��qK�U��א� f���4������+[5k\�=��+��e����dt�`AM�w;�<�����W&s�g�
�/3���Z~�� ���^]�#�tރ.�9��G���ǔ���[�료z^c�4�`� &���OU���(�r�b�H��>�Œ�	�1����6c�ƃ�Z����B����hą�֎�!�U