��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���֚/�뤕:/³��  ��NH�7�)\�ʭ�Y��4��@4��J\8qJӋ�Ц"m1�Q�S�1�3H K)����0���Y:�B�-�e�j!�FW��`�p�~�;��W�]�6���R�1�b������RR�Q8 y���%��8J��3��w> �]c�kg@p�i���ݔ��w�F@�+gk��Z$ޑ~���R�4���$��y˚�d�c�+rP��4pW�}q�V֝�٩���F�yF���=�� ��U9סGї�	����+\�g�o�{������l8$���í�9G| �3̡W1�:����KFW�@�� Kh|H��,u<sH���b	�"��`���_z��U�P'�f�(5D���6s�*���v�	������1��aj�o�CD�Q=��|K��Ju;�b�vߢ��-�_�-��M���`�X�TJ�c��ճ�\�+�`w��x

 ��)�Uf˞e��K#�1>���m��ty�;o�~ �)�c��C�3F�q�~u���m�O�`��v��@ǆ��=�srFmNv�����Qj��5�
�M�~�Ta�ޖ��7h���<[<�MG]���8��^6�B��A������s#N�v���?EP:��A��݊3ﾧ�bIW�i�i�}��*����I��;�ܣ
S��J` s����׶2�x��=\~�N� �2Q0���%�lB֍�t�ؙ3�j�㮮^��aHR�.C:3��B�)��_���vj����a��3����su���:�q�MlN_�N{�E�񗵽��Vh�;��x,b�tG����(�U��0�$.`�~�H=�l�w2R����
� 
���	仲R�1�u��Xf�z��g~�^��K1��ɖ��5	paR+ـ�
lx룱=�;��<W׮��-p��a3ų��gG2>ɕنQxOo-�8��r/�V�и����|����x6� ^9-��Q^|;�
?F6ۯ�=�=�f����\!���n^\�XA	���kRnؤ-�)�b����ǲ�R]����oo��0��G�~O<CU���E��eYH8'Qݓ�j��[�AX�M�N��PϾ#�ˇ��5�����%`�6ڔ��5܌Q|k��<���2��^|�[1SkÃP�����BM旉7×�0 �=ɹ�+CK�v��Bs��m���ߖ�3a*3�?�0���}���c��_���;N��p&���7��;����m�`�[X:�7���҇�d���4��; ոkڹ�����KI��	�c��|�G;\�a==K#�'��Z�y�u�h�K�����֪D3��߾Iy���:K6������Ö��)`��҇�C��G�W�-e\��Gh�
)��4���~��j�<H�+^�f�6�{�78Q#��&����f �&3k��b�9�U`3N��
p��OKr�"f#˿,J���aQ�ݑ`�!���iAPU��t:��it�Z���*T����s�Lvl�56���u.��?�s��� ��y?b8�s=�$�>�ﲓ��ט6�7�9Zl�ӥ��6>�#�bC#�"��Q��
ȉ&=����p�K����\���
R��DmY�&垧�1��wt{gv���O$�E������0��k����D��& ���"�C��t�a���h��!(��z��P���66��߻P0
{m�V��љ��Ug֯,�N�or�?�oD��Re��rp2�N�^�p��=Ǧz�͕l�yIU�.7��]v�3�58$�s��tEVe�.�Q���ѓN����.*s�$�]��V�,Kq��f+EȨ���f�;�m��5�O1��M��csV`h����`s��������92{����J�|ͧāgu(֗}��S���W�2^F6w5*>
q3�㨖�V/�0o�� 5��{�M���)�pѿ+�\��Ɣ�^^�`��d].D[N�$�-�2���	������0�!s�`'Q��96����J�CD������.����n�Ď�7�z˛�b�l�^��o���Z�W}�]O�U���K��η��t
�����~h	�P�5_�H�/�������ސJF��vz��(=h��;'�4�(���a9��A��5�����>��ª���׭d{\�_�z�N�AH�N�ۤԺ���ث��68K�Y����&;TT�p�3�*k�rM"$�8�1z��n��	/a{eyG8���J�����ݞc���V�=t�q���3;��((��
eER��M�W��󸊨3�ɲz���I8RU[{A���mm�
Pn��%"�\vm����u+�mz�`[��c
�ޘ��*��U��P.Rݞ���Ex��
�	�te9E_w (���V9�mi�l�����b?ރ��351�-��؎���k���l{���\+�����h�P���mx�nI� aI������K�#���n��yf�	�.QaK"]C≉A�p���"�W�ΠV\�U�:�a��Ԁ;쾑B�#_�J`�Ђ�m��Z3� ��E"GYI�ew70>�zp���[FP	k���~�c8�pRI�}�ű�$�$Y��#1��}�N��P�1����Q�:��27��¹�.���.�?�%��
�h��1����a�r�1�Ȯ:Iiqx�F文�E+q��Ak��\~Ý����v%�3��&~6�ʻUq�4�����#1��oW��c^��RAR9�tg�E���4�����kVM�٤:����A�����0k@���8��`!v�x�t�1":�Q�]�S��]��T���#M�ި�E��m��t�[�w��r���Ud;2�%��	@٭t~m�����&�D�Ó�N�9��#��:&0�-H߾y��G�aφ��Dg0RNN^@�0��v��A�ґ�Fꐸp>���?�4����?Bؽ����{biB�DD�S�� ��uCtV��N�@���maANS�唚ݣ�����Jf��qúe���0}���ڬt�럾*T]��0����P�l�׻�1�M.��z�#�k�(�Y/tW�Å����2
��q�BcßASo�ưz�0|*����- mf�6˘]�n�s��Z˽Fx��(K���k�B��n�@���)�육��5!�B�@�3�	|]lк��z�ڦbY�֟e��W8r���[RD���	��W��N��Bzβ��������SBS*1�x��U��YEk�fq@�W�1����11�s�&ygr;��\���W�vȣ}c��_�$�!=e�̧��,��/��"��$�֪˧�|�B���ِY��u��#�y��y��+���/{���^���z:�Hg�oG�c5X[0X�SKN��o�"���������H;��è��&�9R:��i����`�P�1����_|Y�DC<���+!H�:�e�S��9���� �Y�g�;3^�u�123��1����%<����=ȇ��ӄŖ�B�{��3������c̜Ow��*Q!���f���n�7���J�(+�aD�w�=��-D�AL���)���0h"��f�����U>�5ᦌ ��mF�Bѳ5����ϭ�e~:ھs�)�?\��Ps����N8�S�Nw8UA͞���1��R�':[j��^9"�#U&�w��n̈́��S c��^l@�"zj�'���t��^���>�TDOG����e>�2��(Zju��2��������	x:��C��[��嚮�z�S��+�:�tt䯼*>��DM�j>���|7L�4(Ў��~��	�����m����'Z��1H�~��}Ѓ�%e�`�b`�w��j�Vqf.��X��^&;�H�\_�њ*&�Y�hg8�J�,�B�6��j�	�w2_:
�"�8�p��p��Zj��qY�����0��-@10m��st�[������AV�1�������w�3h�:؈Z����h� `��ۅR��D����8�SC��c,�2�4%at���{pÃ��O�בf8���7�}��GZ�`�E�e���eÅ޺��i�+���q�1�^����=��ꄀ"<�W*Z�U�K�y�␞(8z���
��BKNgP���Jg$�n��.:�@��d�U�2I���)�p*-z�d�&Sl��CԺY׽v�\oEP�"beHY��تZ~�����Vl�Tc�V���A��W���l�v�zW!� �����1��yuܩK'���g�Ѹ�'���q3�r���*�|�bw�N��4Rx�(׭��u�B�U��rM}E��)Wo�p��.�s����E�N������7��cby#r?ض��ϣjs��E�0�}T��g%x���{øt>��FEK�-x��v�O�#���N"#��8��8����,���>���>+p��;N��*<��������R�<nE�Y�.�?����x���������E�JCQWBΉ��q����T
�A��j'�����������vN�-��MC�Q	��|�5�le�V��	P�	�"Xg*��
#/��:N�\���ۜ�X|����Z��e��W�����s%~}0޵|#�;'x׎0��j 7��UB$1Z������6澉BڣC�A����{���(��&�K�O��.z��"��**��ň,y�S3�ҫH�3X!�Ig���:?;p�mW�f%_�#���@�׃�n���,U��?!Q�G���uFEA�bx��'pӄ���u9��2�H5�	;3/�x)��O�UgM
�|�����Q����R��Ye�:J��/�x���{K�z��:K��ף�X�m��p��E�(���ve�A�VR��t����%VZ��7��� �/L�0\��Y��q��Y��$/�8T��H]!a���ӥo��5Ό1����t��{�1N�=��3\,�$�����-{�5��裛k�
F�9儓����_k��{˪�!���`\0�O$H(������N7����j4�4���{ue,���q/`ڮ�Od�	�b���� �_ݚu]쵂���l��8����ḽ6m^����n=���޽�y\��e�Rm�cX�Ԉ�rҞX&����ƛh$��#\��m�7�xQR��O��T�PW�G�l�*�G���F*S5�Hs���k]c)X�a�w8$�r�y�_������v�՝����TU�b+�]�<�K=uO����}9Q�p�,?�@��+�>7�Pr��Q�����,��M?���
��s�"f�x�#CxI�
~�J:�S��F��d���DL���'t���VUk��ҀQ�X�������ٲǤ��KV�g�?�wk�*��:�j$�Z�^Y�?T��F���6�J�Bj亊���ӊ�W�٧��߮��I$���Uħj�2-`���M���$���.=dS���y<�z����3s�n��PR%�(��KW�'J�K�P"q:�r3�(��-zce �2���[�>'���q� ��*��x����<n���2��_3p��ϐxeE� }"�p>a��Q\4�
���~W�xI�a1y���Ub����-�P����N��;l��Kkm�� �}E���3��{OY�Y�P2>�� %����e��z��M��PR��i܄pZ���{��w\��6/s�R:ӂ�!nwT�%�í�U����z���zAO�9��MFZ�;n����8�{�EI� �b)�#�t�s�9���a�߷unrΊc��U>��K���8h�19xp�c(Ɨٛ_��^�]>߮����'+�q��["]ӢЩ��h����m}�ͱ��
i�v�!(`I�����}R�����~a��y���)Q5Ӌ�c��u0��rP7ߤ�^2�43BYׅ���%_;JHO��.r>��Xӊ��6�O�o/kJUW A��7� L�'�a]d�	�g�fG.�G�r�`�;=Fm�
��%�}?R,��²��?2�n��@=�(��fxi��y%`m�[�:��F4��:�����>%�~��Y�� ��t��a��p�K+�>�C6��P .�*m�>�@;n�Y��䍜*���5e�!6�(|+���A��Tzq�᝱4�WX\Ɏɬf��/���}�d���;6�"�DY�s}���Ø����\"8�v�ԫbr]m$\&qC4糯��+�w<��s�j���e������C��i��V�ׅ-b�[]g�_�X�+Kw�-N��yWG9�md�wM��c3�D1]�I&0�6���@�	�5���� �%B%74̰G7,�+bnVe+b*5O�S�j���"�{^�MW��������[^�Xl8T��sq]@�E<͝�F��@E���:�H�CIb2�ߊ"9`2f'�O:%��/��A�(���0��Z�L(��	uP�%+�~�4v|��J v0�=l�� ���&!�.����ot39u��_�⾥��R.	�&��+.CR,�5�M5tc�yW���)um��i��uRq��#�k����Jd}�s[�]j���	9���DQa�&W���UH�G'����_�;������P�i��N�ˇ4=���-Z����9�r�]�.o�.�(�Y�f��� �,��3K�A�4��(���P�$:Y����"��U"��]�)Z���9Q	y�e��>��jl
�)�l��56]=����	r"�q���p�VKU���q��5��@K-.�[)���_�cW��1Ņ�x�߿�wV�5*��J"�F:���"s�Zӹxs'f1Q&nw�Q���� �6����)��v���?/�4 ��w��0�l���m��g��7��"����7:��8�XS ���A9@��ؔ-ݬ&M����	��i+l�?:A�ƙy
Z��n�63�C���Ł�sZ�w� wCX�����w���Ls/rMp�.�`؏k9�dVSZ��뎣�j�	��O���{IQ2���]i����2�٘�ǡ�zN'|���@V�c�KL�<S�����ՙ�'��
E& �p�}q�݂�Ɋm 	��/2+��)#�6Wo�7H���|��Ў��/���O.����@��К�.�3����w�-�1T$Ww���o��X���H\�f,�9����ⲇI���ǡ��Y]@�,�[m�ͮ���p��Q�xKl�^��]�a������f��|V�b�Tr���'A{��<����בZ��SC�}��K��`7���G�I����H7��j�1�՘⩌�H�~04�J��#v�U�]�f��\%{=]��V)U��Yt�j��cG���^��6A���_l���pp��
8�t���8n�DBHM��o){��=vZ�N�I��T������ !S%hȈ����߲sL�a����4f���)o���}��w��"��L`�b*��Q��6G��:&[|w���I�����E�>sIPo̿�J(���cnlOʂ���"�J�a �J/��Ԕ8��`�HX ��LN������5ՙ;P��r�J�xx;V�ۻ�j�D�-ߍ�����2>����-�%���f B��=�'!�����HB�L�q�í��ѽ��c ���n�{�Sј��Y}�^YW�U�
K�i�-���6%�^e�Q���	(�'+��p_��u�ցP6Y{�qx}/�hȨu�����������C/Y5֦C��+xޠ�<ʦ��BjM�^�3��X�E6R�VV+e�EM��b͋'�����7qf�op
cA.PF�e��M`X��Q#�X �@��ƈ���!�rd������d	O[.�J�;-G&E04�
\���r�u*3��ۃ|�͜��]
��)�׹�1�%Л �o0P.����hy5���c`��d��!G�d9)�"�LbXP�N��ȗv-'��u����X�����\O�����CҀ@Y*�p����ܑ�}�ޏ!�- ��ώ�B��U,�PC���嶮W4�V����HC\ȵk��0�)�1��t�ٟj���2L���A'��ڶk��j�b[bG��V�9�nU�ͪ�d{�aU�h$Oڨm�uҩ���T�.�	�3F���$%ÛNw�Fi�^2�R`�2L�*\;�V�H˧g�h<@)����YP��uT�3���w���6&����h-���Z��M�"F`���UAvp�OpD���0J��\�H�C�\��F�4m��ۂ,�R3��AgVn�h!�|�f����\�(.�����VO�ʡٲ7>�>}5�	�*g\�>�@��dx�XTOJ�����.n��4ط�n�8J��f�QbBG�c�к��G����od�ܤ4�у���%�y�pDR 2/���N����g����܀A�h�rN,��<����k��H'����B��?�'U�}��6*�"�S
rї>����A
�������a/��-Nl�9����U�<M�l%�ep+�UL���������x5W�� KF����������N�ׄ-ez8W2���Ś?���ۉf{�iݩ��� 	櫘PeIZ�| �EMB��NA���Q���Z�[t�����Y��L/�<o��`yD���\����Z�e