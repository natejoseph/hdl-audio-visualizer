��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��"涏K}��L^�L=����RZ��i���)�6@dS7�έ_{[�2Ъ�҃���j�׭+j�Ӫ]P@��HQY	đ�kp/�F�z�5��с�08�r��w"t���E��|1�>:�hj�]	3)m�+n�[��(��
�!�u<� ��@�|`�A#K{����X,�#:!r��o�2��V��5��0�L��4�u��2�?���E��a/u��;ܴ����(L,�=)��X[&8`X�$���B�Qi~����y��ow����()�qmXHZ�B�K�w���L�+�:�ըw}�� M ��lDw��	�3�?�T'�c)���m�Z�{#`,�M�ii��/�u5�Q=!�A3��eG�w�K�s�ؐ��󮒍J7���K_��O����}f%��c�i��l��B����9%z37p��Ǯ�˂�<�	b�h���zVMk����E���>gT�5�?���(�EՑ�(*e�����J�a�u�+�����;텂L��?u/6\�d��}��WL&W��1D�E�ÑZeЄ�b�]Z�2��	�Ƅ�,Z��:���N�Վ�7C���ц����m�*'��ܷ�Sen'�F��0G���ҩ�e$w�`�չ�O�;�Ra�ж5b�6�HW���S����I���>/;,i�����&�~��g	H@H�b��餤 pw|'����82A�o����6����D3����
�׽S���"U��I��kz�?^H'x~�����u�;�����|��N��؏�~��\MN�N�e��^�`�j[�=S����y���֪����u�\�Ɵ��(�:�4Dl�z(9P��3/|?TD>�����u�|�j�aBj�;�#x	��'`)����z8�����0��n;ߢ��s�����O��n�MThW����[��jѣo��`�\�qqzӦ�\R Xp�5��3�dß4��h�-����ga'*fg��ˢ
��ߚ�Ys�Q�A�l ��;�ps�wS��I�I�hs��d!dR�߹��w&��B�R�Ӄo 	L�S�����L������C�7!�U���+�� �R}����*&�t�*.��3��PP�<�z���P�a�hyCɼ�}��ˀ�/��)�&�q��im�/���1��`;�<�V��焭��M��30��a��>� e3�i�z�j5S���O�F�=�qT)*gi��=�e���mS�e5HsY��`3�g�aR-���]0�4�X-�>�λ�R#�ʻ���-8�.o*_uYCy���r6MB�
v��a�����|g�_~S+wg���yAKx5ckz��ފ���Ҷ=)��9�Y;j!�efT�0���s�)�h:�s�4�
�����>c���Vk��wd0���S��䔃�π�ъ�@��/15s�,ֻs�e�V�f�gU���L�q�^�q��'pܔ;2&�7��@�OiD1�T���$V�m�6�5�ü&g�� �v;�6�o���PGњ��LG��2h6�I,��fbl��y�%�?��'��P,�K}-A0�����c+ɛ&,�q �t��F|@j�զt����}�Y�'�>�<FFO��d�s���gJ�g� �EW&�Z��z-�9��.�,���D:`�9����Z,�,���+9��A9֪�֬"�6���E)�:)�T�'f���P��U���E��l�>�g{��fZ�Iu���N�A����VV-r�`\)��F����ɗKm6�����^dp3�x����w�'��tX>�
;c�E{��Q$�m��y�pg�m��"��F�Q�|���}�m�&�,���F�Hp�V��p\��c(ڝ~��l쫮��a�z1K��ϿWO1�ܰe��]��/��r�R�����:HcP������q�%6�� ����l�GlNE��./�.7v:(�u?*�3_3w��vv&#x	/�(V5���Pi~o�b&w�/�ӆ?ѯ������_��C���j88�bTOа6W��u�u�eޒ���j�h��l��G}�$Ҏ�C�%W���!��\%/�������dx��p���GA� _�5��P�u|T&g>'��?���^:՝6�e8���i+ c����m�P��rDw�Eo(c�ܗUk�>O��c-��D���w����\���2�4�1�����g��#����{N���� \�h��I���e��)7o�q�=J�����B�,OX�J�# ����T\�����l�Lr`oy3�.�ȃ��+���О�z�>`�7i,�o�N�	��|�����Fz^�	�^�/*�\��#�">��ֳ@[��� y���(f��T(}�8"�n�'�ވ6ׅӛ��A�Wh����N6'���Ylؾj��wdW%�1A��;)l���M�N��WVY�JJ��6��t^LdX��[i!�A#׆R��5��Ѱɲ������7瘢Ue2�Y��@�!$U��A>�Î�/�<���*4Z����?����p�<WDA%o�3pLBKf� ����9u�DkP==��^�a�;%��"�E�sCO�+�LP�9T��м���'�k�]���,h���y\�s�9Z�mb���D�,k����c0�d��BT������d�t�)$-�ݿb��?	�����N'�b4a̓����+�G�8��O4b6��Z��^1"�=���Y���l&��Hg�N'7���ZWm4�Z+/�?�9�Ϛ�&!���kqw��X�������Y�#Vf�3fAě3�B��e�ħ3j(~�A�)Q���\�4�������6v�����E���}(����]�9��H$G��m��0�	�.\uF�gӚ� ��|Iۀ��O��פ�UF\9s�J�ن��N	A�$�C�W�Qk�����l
��^���.@kZ�ģ�ph�U�O�˪�O�t]���!���別�oY�ǻO�_���lU��	Ԣ=�o7����	
�¹U%�
�`�a�֥�A����΋�5�U�ںU�IvI���04�P89�׫E�����C��O�*\th�^�Qa�[�p17�h�p5��\g_ra2a7�B�Ej��w�5�1�P�O+�fQ5�S/6S�+@`;�<#�,:�,w�=�-z*@�:W��jv�����TKѧ)���[wOx��R=|���Z1�LXj��1o�4-5��paӱ�����t@�R�_�=�el���	Е�~;Ɵt��ky'~�
����w+�9���Q7��G�2�_� $c?�*k�oЫ��Z�a�*�z��)�S�v�FBzw��ϓ��~B�����@�M;�q�"����"e��;�ZI��dtj���%��d�JdƧ�r5�>��dw|h�=2�"!n�e(��0���*;J���İ���I�9MG����"�}����k�x	1�7q����I�>;�ߑsv�#w��T���zƲ+���?�Jk����K��r{m|�uғ�BG[�촼P`�41�ls?�GZj�5�ߧC���bk*�t�d�]OD����_Q ?�ī��
E�{t}K	ne5��&d�{�z+�Ro��Ro���F�Gz�,Iʡ����C�T:�[�j�s�tt�ċDM-����C�/@zWV��+2<�1�[���9uQi~;��n��KZ�K�ىV�I���(���j�I"T�pO�ەG�׀miQD�y?9Dj��1/ќ���|x,l��@RX����53��Y�pi�̻�����`�	����o �U�������J���s���_�_m�R��wt����D���pl⌎���S�	��Rpau�r<���y�,��gM{K�q�h��fC�����z~l ���[tb��b��ګ#����)@�D`���V���Q/�Ar(�o1�_�.!ԫ���;��l 4�q�C��m���A�� �A��Bk��#Ҩ�)���j����w��B���|��]ю���~�����dG���SC �c�״�QA[�|�P'yN��+�$���ҳ"�R�m5K)Y��^��l�>#]կM{�f?�p���I��T�<u�|H�W�w���o�f�;�y-�Dr���P�Q�O&ΰbDc��/Fc¾2�%*Iwd�$ŭ]�u�����X����n���p�jn��@w�Ԉ�?~��������j��v�^����<
�@�Q,�M��^�:�qy|E�&l)�P���
��Ѕ	�9�����*���F0���f�zK����S�%�朝��&�R���B?{�/~a�I������X���� ����87#�y��F_?o)�˺
������6�k~/���v����k]:A�����SΘ U��� ���$��f��bNK
��Ku��=���d��:��3���Do3�^�
����c^�/T]/�bK#�!�[����fI6*6=��mf����ҭ����������L`c�5�OPl�<XA�s�3@}�/���!t���qH������R������4���g�d1Y}c_l�9�j�? }����B�(i'0���0��ͳ�8�Hdf��Ҝ0y����^��H�>1���7��1M��ڶa���GR����i!������66�AL��2͝, ٕM*����z��
�5(ШĮV��S]��F80z�A�_��,�����1rɭA>�9B�=�}rl{��f�uٙ7�9���{k\8�9��-p��5����͕1\ �+�f��C�;c�N���ĺ�z�[['a��xb���jL�Ζ�h́����j:  S��R&��GCZ���|#N#�`��O:�� 8��mI�Wx��`����L]8c�����$���}m��%�g�e�8�
��D	q��������-+(v�. ���Ȣ�,c�w��'Z������qw��9��0�[�6)&(p���a�J��0��7�|L�I&o���psR�˕�)Ձ�ݜ���3lڃ�Q#oUx�+��\jC�O+��8�nV|o��"�$��Q�ޒy���p�'���.r|�����"��k)����*rg�w�EV�4�&���H~�@�ǉ+�}�B^���������)���%{��(:�8�,\c�V�9����e�/�3�P�J]%,$�mOj���r`��?��M