��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��=HAW��*��d��JG�Q q �$3�?b�~��S�APH9�C�q
��gft%*.�M�����Φ��eT^�ېiM���|��
|���i�%(s߿;����g^�e��KW�W��5�>���}����Ι��!�E̒���Q�Q���GX��C��l U�(��fT�o,C���/��܂l��(p�m'R�)8]ѩ�^�Z���Q9�6�ZT�\��J���u8�pS���~-�=���r�=�x�x�� o.��jR�\x�,^���g�����l��d�F+6�6$"���1g�hp;��PS�G�Ђru�x,`�0�)	�n�6,6E���@�>:����w�&���{ E�]��4WB�F�m_Oz�I̯d��Z� �K]��c�	�ӂ��Hാԕ���==�q�/�aP.�)øy��
�;A]2<�;�
@�	Cx�A��?�)�i,6�uL��¯t���eݏ����J�\ΚM��߆gЮ��H�Q�4H߯�.�wҡ �mX
�׋�pNXcx��w����Д�M���^/�1cf3���ǁ�?���4�`�GC��47����K���z�	�e�6m�r8�����x6')�@U���ˏ�R�x��n������X��47�����_su��A[P����t27���7������x�a�)��ފ�ٱS�
�W�H���Y�eE�j�T��6*R.^���Q�!b���r*newz���
E�~��sC9�����2����U#��ϋ�Of�p\W�.�Q�w�H���3�䧠�����`���x����襯�� �b�T�`�����=�U�+�#fTg�R:ዄ�0��+\Cu5i�ݍ�^B��,�{��:�!�v�|��G��J�д�<�I�rRQ��c7��Ԃ�s��Z
��IW��)ׂ�u�8�7_�Ec� G��c��Wx����C�.�ݐd9_�H�i�L�+3"��!�/�� �4�f5�8���%�τk����vt!C�gז�9����P
��(�1���q��.I(��BHaB6�A�o6'��ò\Ɛ�\(�wʟhMy~�l���D�c���!/�+󉷲��ă���sR`ۅ��]:�P�D�e K
S�v���7��iL:?M���cj���X�y`=��9��0^�ʆH��r�\�2p� Ts4�|�C1`�Ep��ȶ�&o��u� Lz��#[�����1hWs�t̤�}�����a�n����7�)G��v(S�����:[�����	�=s)[V(F �� ���j�SO�A��p�[a� ih$�����b	��Ы)�:ȏ	���k���E�$��K�}��Uv/�iu�U�j��;�\���^��rU�o%�D27�3-�`��wj�W#�h���R���0����Qs^���= �x�n@C�m,h�7+��B��}某�)E�u���S����wz���[�9��e�{�I�I��,(���ؗOZ�Y/
3��E�`�h�e/YV�W���c�QT�T���Er�����#<ّya1����]J&3�C�e#V#i����:$8�I��Q���F�l��y�BC(��Ay�j"��cM����������]Hh�1��#�Y��x��i/��)��R�撱�j�
�`��l{?���Uv?j�3���4��@}{�N�UQ��b?��ۓ��a�9Aj2�HR��>��U�*r,	���\P��*�!�����F<�琶յ&N�(H�B)�,����S۪����q�%�kX?k����"��ܹ��e�r�f����?�P>�B�iF!"��v�D��	��1����a�^o�(=ɉ�3n��<:j�6yt钊�E���͑�b���!��2�Ӕ��pn������I���|O��� pfn<)��
���ѫ���0��N���j@�y��_A;��Yp:�0��#XL*n��ȟ��nXj{�u!Z39Y;NEk�X�����.z� �&o(/(���ϭ]0���G�O��1�𵬈�E��{��K��a-�*6Vk\u���5kEոH2F��K��n����H|/��_._wKؕ��R�
���5�J{��9�I��2 Bz��������iYJ��M�,/��J)z��Qd�%!W뫤�q��}��l��s$Du�f Sן �\�bol���ub��R�M`0�4٘1iS�Đ��E�5��T}�Bw�ͩFz���oN|��Xb�QEۊ"���wjC:��?u0�E���(��a��)��ϼ˶���K
4EIX��<J�c������n������{�~4L���S//�ڮۋ韂�=e�MP�CR1�A�|2f!V�}����߶l�x0�Vi� �À'�lg�q��6��ݬ�-���>D��������>^"����$7e�a%x�pO�4}���f�� �E�6mx�^-��.3�o��B׏-V�3���A,H�B�K��^~4�oҟ��(*�_����wuJ�Z�G"�9��5�v��M�-׳n�K.$ \�k�k�D=y� ��1��ͱ�f6Z�]�ѣ���"#�?���HI�Ϙ���|�\:��"��{0ڭt����Z����ꨅZ��:	�T����*k���f�b�V�]rO���k+���p�5�3l'�4v�i���*�hIz��l�j��X/3�=���LIL�b�3:�uE�4}t�x������Ͽ�2�u��$���E��V��*�Xw%T�F[l�cz&ъOO�*`�]�Ҽ�}�R�b�j�J�,�"'���b�x
�v���L��a���_R�t���:Zz��<���-.�����4��폪6��W�K#yC+JN�Cpa��:������l�g�@(9^�c�ωB5^�ɑ!�S�N�ۏ�Pd�= U�m
��r,��^�⌽lD�d�:ü���$!ST�C��:��:r��x�B(`�ޅ����<�೎!M�徿�	�� _�l+�����a��]_e��47jHS�������	��I����B�w�����2��~֖ٶŶ8��WlZ���9h����He�ъ7��p$ȋQ ^�Ѯ'S#�۾��\��''����0��7�����MʵÒ���{ӫ��]yp\O���o��	^�a��܈#̌u�, 4.��
c;%�Sg��^����{�!W���,����ւ<�DQ�0���T�k|_@vV'�l�1i�@�!v:��[�;��иBǬ���e��pCy�{�\?���c*3��sq��
C]��9�:i�G$*t���|Q�](�kn`���[�8�����!6��lz:?k��$|#�S��:pZ�����%���w�KEg�?�Z��9����L��X롣Fc$j�!�..�;�vz �TK�[�<�U���3(�ta��q��xl�C�[;�����"B�ۜ����K����Z+�B���ak�a�0>G'���"@F����<AD�ːx�%z����*�@#F����1������7);��$v�Ma�j&~e"HP7�>}Y����R�'/���9�40�������+l�PX$�b���3�0��zo��c�Z�J2���ySt�|8��)�X���#'ai����zI>e����K_�����6�dV�D��a��P��V��I�O%�Cd=7���V��~�|>¶���$+�fM!�����ag��gc-�N��\�!�8m{�cdt�n��r"������g��v�q��y��X��<,�\�abt��uz��ۺ�
sGj�nu�1��1���Pο O� �
�HEV�Sղ -�����%�������ϒ�rgfTS���xݪ�e�Υ��W7�O��Q�i�?W�_��:��.x�V�D�KR���&ChN�:~���&6�2�^�S���[M�J�4��E�ӳp�=�(|�º5�(���x�"�D6A]��'����;��Y&����CA� �����4%������Cum�׾w��L�k� oik�������</���]v�T�'���� �6�ᮽ+�s�I�o@�.�B��}a�>;YY�o��җ;��ї6��(�ҕ�kT�~��K�:�J�C��}@��)�v��{�6�Kβ�s����ϖ�������*w��f�H!�E�E�&�Q�r�[��A<_^��� ���FJ#u|+f{�az�� �@0�b[�"��K<�k|����f&]b�" ��!�JV���� �ۅ"����N{7rO�A}�Z�2Nk�E���5Fp�>�܈jD�� ��5��[i�J�p���"�~)�Gp�z��!������ ��$��7a�>I�����u�+��C��4����Pp�֤�-��33ӳRj�M����g�����m!i����������	
��Y(���xs���C⑾���y�.T8`=ѳ���l-�2Îf ��=mT�̋�L�@H�����ցj��viG�Z��i���V���\�&�u3�Q�dH{l���q�{��"W��0=G0��[T֗��c-���[���IIG8�P`1������E�5���n���ߍ:��Cm�@�׺@�(6����5��"Z7��Slt}{�p5�?9g�F�������p��k�����z����e���y<��>�C�ll�ų^A	��}+p�X�n��l���?�h0)���ػ�[
z�t��⢇�u��K�W}���%�(�Md�EJ��"��ˉ��s���#��4q�Q�?�=	)��-��/n��lc�x�S َ�+ت���M�b��$�����p@_��$����Ny�d���!���m�j�#E��_-Rj-��\I`�F�f��Z�v��=�p�P_����`��]��1��^���Q��\�5ˍ?e+�<�g"P3��j����o�g?�w߅��L�ڒ��?������9�#�ts}���	(���0�Sv�(�m�O�0�B�;������&IFޙ��.]�$0�k7˿�׳�'(\6��7���^G��}/�bՙ�k��b�wm��זqNr���_�t��;�4�i���iUE��?�D����M;�_{0b<y�G�<�w�px"-,U�YWKFex��	ʑ ?�Z��/�.Zg�s�ݍʬ�Tu�?���*b���Q��u!�	��n�eӠ�xo���eOm���hI��T�<�K�2�Iݝ.��>]}>y+�'�V.Q;Վ�i�K
�ۛu�SIu�-7���C.em ��{���P��4`Iږ����V��#b�e91�Y5�ji���ؓE������s�e�2�p�����������үs9�K�3����3�$@?�%&�S+�Ȳ���Z�U��Lꯍ�����uw�G�5�m��8�Y�֮b�#P�����b�В{׆C#/:_k^���֔�B,-���dbT~eD>��ۗ�K�kfԼz �l�Q7�?q�o�!p�Q�c���2=��j*࿈j��Ek�@Ԕn���7X3��.[ԣo�1���͂�
��&��̛QQ���?3^�7�`��3uN���V�Z���U��z?��wmviO��J�q���=��wZ��3��9/M�Q4u��K�[�
}�� TW�zՒ�B't��O�{�gi�s�r�R/�0�k�l�x�ly�˴�y{-u��e-9�N�.����k�z�����FV#]�$�X�m�S�ˋ~�Ap�2~4���>\�wWm��{�ڕ�p��B����`�!�m1���F���7��#��j3��_b���6�&蓓�x�b�@�j' !tp���W�#�!s��^%���-�n<LYC"Zɹ)rȜC���g!���,�#�Y��.��H"��r��3���Jx��]DLLx��!�����,�� �S���E��/�;gg�$�݂,�/䖄����P�bz�UJ��W�N���h�'��J糐�ɣd�T��q
67�ON�"e�H��V}2��_/R�J�|���M�	���	�%�������W;��+������i׋��wܰ�1.��.����eP��:VS�����$@-�vѕ��ޫ�'s|H+?r}���?�%lhїQ�j�����Ʈ�ώDCo��_��?=_ȋ�z����[ݐL[��7�^�q�N��+�d��_�+cb������x��v8WO��ZU�t��EM�"�tS������b2Mf�޴_�B�.eT�0���I�t���^�b
�/e+�dK��%?�5]X$�e��LD�&��oS�X
�Fɺ�T+���&��\@���NΗ�A����p�PR������:��$e�8��:D��x]�ᒨ��*��,-Y��$+��E�ٷ*N��>��D�q��#��@G�%i�D�oFNh"���(��q�N-��)���SڱU}TL#2���H�C��ɲ�g,�vAs��z��}�4�$-���X�	�K�r7����hΐ��R%-���ّo�uh��X�����$|3�|��9��l����܊�G 0��38���/�	V8�Jj��[�o�	�x��C�i��#f�%K˙��z�"�]�������f	����-R�I�fcG�f��QْP��1�6�����3������E����6�N[� u��Y�a�ؑ�["�߬���e�ɷ�x҈W�z����wB�S�<%y��V$�$�'z�~Գp9/�W)d�ݫ��e{�p�_����֥�����s"	��僪ċ��]��s��Nބ
�^��¦��FkR��戋�q����ty\�&�7c�^�!���.߭e����t�6��1� G T���f��aP�2�WS��ZP��םR.�Z���[a5ǐ0�
�qӘ�z����t~{vbz�Q)� %!�­L'7]O6Α�8�m�T�'��