��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�l�(���qrM �Y���L	:�꜂���kL�t ���%�M�}^�ц�X3�
''��".��[���SA�f?�Bk%��*!>���o�K��HyJ�~�7��rl��P��n��B�� E���5NR���l��?���b ��v�{+.&��Ү��ȥh�@{[姟S�1 f�$ �,�_�R��Ψ��'7�c��M?��Y��N�Q�~��B�ِ7�%���?	q����5дy�N#.+�u�����w ��3���c�M���Z�����w%��<��ze"��<��Í�uMSq��Ee��;h�a�!7���'N��BK���վ2���������P�c�;B�j�W'3UI��	ݝ��Gr��[�J��F�9�n����4���
.YF�Q�6�N�� ��%��!�'	��Kg����|��?aucs�^1�Ϸ�H�Sžǋ1���,��!I�Xɛȡ3RҴ���@�1�n�`O��`$25��e�}�6�ZC��f�l�m�bՏ�z2���y��;\����T��n>�4+�WS��vr扪�tg��H|�e�4J�򁿖�Z��L#f"6���·.�v!��0���*%�U��D�E`/������'i	��R$#_��ώ����?;���Y�������$����e���g�"So��'@&lL�����D��ֿ��sF�"5%��`�w��c�����"�%��c4�u݊+�Aɛ`���E�9�AD0)����G���nl'M�	Rz5���_�F�_FF�����ܹ��~2M.������Z�3��t��q����%w{vޅ}��>�0?z��<��8���@��{��6�s��SG���(�P\��A=C�C2i9�k���{L�F4t:K�G��ja��k����T����4�ϒ�2VD=�Z"�0��c��Ī���t=(��rk���~|��Ш��cc�bB�Pmmg�����,�Q!]p�����ּ&]�4֪��%�Й"�<�?�e��S�q�W���؞����P��"@�Y��`�%l�R�0�S>���E�e9��B��蚭���~�3%��7�4U��o���1��;��D���5�� u,�i�eT�cV�|��E�����M:�uk��XPz�X�W4~��{=�7z`�_54��ܔ�.�!lD�5��!�i��e����<D96nc�����w~�B3��#<K��.~��f�s�e�x󷁿&J`�4y�|{�t���r|�XBƿ��@w��F;� ]�`�G�E�k(�g3ܜ����-�N�^��zX�L����h7_�)�9�>,4��h��+�F�&uR�,Ch�ȷ�o��e*�㒄������J�`�1��?��oм�H~О�k#�P�� U��Y�U&�KQ�����J��0X�p���.�e#�ƺB�\L��]��X��&����y�5�K~��S�'1S��":��W7����7㢞�p77`fpeF`|`l��D}`��JK��͙"vj��	PlE�e<:a̳��yx��^3��E@r՛�@�e-�P��W�����1��dS�y�4����{�PG[g�RLL��61�9��4T��Kr�m��8iQ�/8N?�����!�rW$��E��x��֣��ژ�[go�[���A@��ǡ�Ȩ }1J@�=+��:B$�n�$/8Ub�j�M �>#���7\�FIu�ըҖج��lJY�6zV�@1]��|]sD��cg)�u�QI�=��.(sk�-���c���:N`�Z%�y-*�l�A��#����J C6_���<D���52��"�n�i,o��o�(�5�gU`�*X Y��*����o!{#�I��۠�t؎�
#�b�i/J)N��g)O�p��o��f�	u��	f`�{�##�����4�b�9�CbPt"B��xZ��4gόZrV�A��.�܌)հ(y�vj0��������hx���{���/4��ܓ��-��2$�����M7&I����k���$�� �Z��������w��4Jo��a�s�����s_� �OoC/>ù�
����܋�����X WyM9�e��Kq�M\���<��*�ڒ�K�B"q(���4U�Aw��nFWQԠ�o��V��"A��u��pH':/m-8n�sr�/k��EUo��1��A�s�B�[�$�y�Kp��MƉ����.Ђg�ˀ��<��N9������ͯ�C�D��Z�=�D���-J"8RD�!��8ǑQ5�+��(�O[Z��=Ŵ�]�f�xk��C$�y�������D�9:;�z����57f�i?�#nOK?֚#Y��jWt$IY_��G��xo�/4��7��[�%Ոe"�>�����b_�/�h5���
!�?Mq[���u�"��>�g@�+�����=z����psw�u�{wy�VZa��CM@[�o�ի@��k�N	�3��P�5���i��Kr�acx��}����;�L'Xՠ"@h_
��T4
88ϥUKo�<�-;�P#�0�(�8�u���� ߗ~�-�u7b̊Ĉ�H���,�vk�o���_�����E��Ұ*�`m^l؎Ěח����0Y��B�>)[cc �ʭ()-V�D]iӺnlܪ(ڍ�`q6*A�T;�7 ��<{�,�����
���BP~�B�֒�*��̘:-���	��1�ۃB���(_��&�P{3E��#V���L����H������z�$�j�r�K�q�zEE%�f���/��o�d�(���QK� ,�2����w�#�6�"#.I�V�|�Cˉ�;�  � �0Q��a-�+�KJY���Nzl�
m2+�kJ�/�^Ȑ�����'�k����$J4_�(���^$896 ��_Y*�1T��_�� oI����[-�~���L{��t��0+�j�P��>sI~�`�G��C�
.'Gh���⥫�N	kF,�Hd%�P<��m�J$�����}�?���j�EQ~�o��|V�ۛj �-���4\�j4��Õ>et?NLϰ2 bp�L�	��͘mgsi�Ŏ G%tv\���������ە�몥�*{��&��w�lr��T?�_���Y�I���l5��E��2��U�ړe������p2L����2hl�k�TX::�Z��	��{bx>w$��˩��\�aYd��؛�_��[�Vx]:��)�o������2Q���.y����qQu�jT��<@�͵\�R��5g�D��}"#Ԁ�g$Z^B��gѰ*؀�	�_�A���ɂ@|f���@[�Á,�/KY}1�n�Z6��A��5x���l�瘅w�t�J 2�S���
E�QK~B�C�a�#�Zi��R�[j�����#56(�G�@�,�{
�f�'�By���K`m��ER�^/��ߐhQd��<�!�J�� i3��+i�������V����0B�p�
����{�q�� ~��@��e���y9=+^f[֮��!�����}x 4BtbM����_iF��_�u��p����t��1\���U{��j����$��Ӷ(1�`%g��6u�?�i]I�arHZL��W�Ļ������]E��5K�����}�g���7������w��Ͼ��x ���9eTC���$�Տ��s�{��|��$��V*����D������7jXm.���w��/�������7����8$Qڝ�b��e�� �Ͽ/b%��H.)�R�Z���^�nN��{�X���g�����!ų~��i�+y��D=*�x9_R�� xeeq����%��њ��`Acף=�o� S<���~��Q,}�t[���7<��̭��L���4]
Z�N����N>�>�	1W ����I�IY7u�7�o��r���_u|?Dak-LX��W��ܶa�j�n����f�$.����j��C���!㝦�:�(�/��<I�ewA�初Yn��9�Ngqzu	��}b���]�q[�Ώ��,'��Jp��'~��/!����	Յ��VGH&E]����Y�Tޜ���"��.و�!��N^�վ��/�����U�pjF��ڙ �^������+D�]�ɬ�l������\�Iu	����Xd���Z�� �g�T��"*тn_�f�E�oKofZ����_N�F����$�o'	C�OkN��0�����g�!X$��G��K%vc�4:��k��u$s��n�l�'C��i���`�=oPHl�zC<�	$6(���@�^WR��M��%&	d�T�i<�#�Js���vDA=�х���?'*F�q��F�Z�[��z�Gl�}�*x��+�"�dh�0p����0�y���fR�:�GWm�{�&=c񪐤�0�@�� ^?_K)�~���q�5L^,}�R��rWu�	���7Mg|
ԜA���AN#�7;�Sw~R-����sбL�	r�3��rIz�w��Od��M���S�2T��.0[�5��/$���8FX硛-�X���)+y�<~����������/��pP(bƋ;Ў��k�1H�|��q^�B~���ӷϋ4��AK�H�8)־Z����*�l�n�+��_rۻ��.6�����9FjD�h�> Lci6>�)��N�H6��	�A݀N�X�A�]EI�x19�6{��j������Q{�(]S��
��Y:�(^0:�?@��~�|OcY���9"��\��!�y�y� ��.0x��dq;�-���������0T�d��n?ˉ�#��;�z�S��Q[�R�(7()��G�q�%kO�_�@��?��C�=�n��������я�Y�����j��M��� FyH��+�x�=�rKQ��^?>k5Ov�b�!H����G�"4�C� y�
���6������|凂���S��z��N|�$���tk��eQ�3�D+RM'q'�]��\b����O�����TCߪ�7�C��M"��2BVd��E��L �|[[�J�{|l�C`�{U�����o��̅�H��"[Iɳ�EF��[�'H6SF��&� 7�������+��
Lm`�����'K �j�����4;Pށ?�΍�58B��U ���k+q������`Я���y�e�����ߞ���#3W^OE��t�H�.228v�8n��3� LXH�={��mg�.q��%&j�d���Q�!�{h��_��P���$�?�!<��*@���s�tLD�j$��sqC��Ľ~_��[Z�u>���W���qx�bǷe)c>���[w·�x^�* H�%rt�e.�?	S�0^�����#m�@Â��8����.xv�XMc���P1����v(	{t&�@��]�^:����ogXL���%h��v��MU�2I� �v�p���&��X^�j��L/wmV`��?��$-�[_
O���g��Qu��/:5�-�����e���A���
=s���cS��5�\s�Z�O7�lJ�Р�3�T��F/��g+x�mCI�4�ys�S�R(M�cJ�U�wb�U�+����j��x��nc��k�M�o002%m�n	���2ȓ��~F2u�iXH��7�(k9�����Bi��]��z���	��2҈�jRc�� �O��#!��P^��e�1���7���=ݎw"8NK�z�3�e�1�8��'�G<Ns��x���R�<��+�� ����nn�I�-�I����9�;����"�Q˓��h��W�j���
D�(P��x����Gb�2�b��L�a�"�#�]�Ф��u�$�.˙���rʧ���+��,��у�3�c�"�
No~��w�X͊n,���w�J_�(�7�����*�UC�H�����$f`X�lV��G�_�-@��![=x<�u���� �6C������?ݰ����ι��Sd)Ʒ1ݾ>
l2�.(���Q���Q��Y�����\[�� �~�ȃ�Um�3�0�h�����+���E(�� 0��"ߚ
CR����~k!܁��ĥ��$�:ޤo����LF7V^�ܙ���'���La��c
�)<���G����6&�/8��v�o�æ<��
���8�+rg����dD9����h���i�K]��
�$K���M��`7�;�i�M�:{�g�w����~O/ �R/��:��
)�4?9�ѱߺ�B�4}t��jr�6\�T�.�B#2�7�)��$T����g4]���-�B;zn-�A�rأ�+Ffd��>D8~d���W��[�>7G�>�流���C=��c�v�h���"�0��?��p9F�;l$����BeojUˠ���ӇfaB=�+�a<;�lT�>����:�^�w���
��ĳJ��g@�?8��|��p�&3?�Hw�aw_^0y��Q�xR6�yB�5��Qi.�N�y;~��&;#��@=Ly��@ܻ�
3� ��u��p��=h���I�05��v���ެ��z���
�(�5Oi�(�.L��K�5��N��]2��P�*��B�!�'��� +�C���-à�m���;���`80X��#��Z�FW��ܶ�^j���'�b����ւ7��o'�ET��,�o5�i�3̸���9�_b�5�n���}I�gO�d���p	3��$�"�A9;B�t���.�����r�s�R�����Y��{�z�����o�п�l� G �X�}�颮8�O0V��,jt�uB�,q��"Ďӿ=�*�n*���JE[,���~�n��8�ʖ9ŉ�Uܑ�s6\��uh�����&�Y�~mx����cR��݂�8�*f�i��-�� 2!G]�����G�6!�^Ϧׁ=�q����K"�:����~�����1��Ɏ?EV�F�!7�Dn?��8�_�"�tA���YuYxeZ7j/�7�ZAҘ���}O{���EY�#4��y2���F�勱�5z��	�6��A<�_C�L[V�WOl��ѐ�tY�#��ë�g~�D��.����U��>����\(:�lRߐf�#��L��z�N�� -�Agظ[(0b:b�U��R&���\��r*����n��!�~~҆lp`.n_��]ڠS�!R��1�xv��Q