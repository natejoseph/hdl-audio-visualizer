��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CG�ʜ�S��m����uf�+��K7��'�3�JՎ6� �*� ��{Y�c���H��^�\vov�*��F��N[:G"*�ٻC�p��0\(���ix�]�
�"=��UQ��v���TL�A����U;��!?B)�+���3��L{�m����G������.�$9��0���z�$ ؗ�ɗ1��,����&��Pj�^-�-5�LXA��?�*|AMA�g���=�CWH(�A"��&?)�\��	�Or&�L�	�oT�6��Y�*��(�5���h�z�:,�^a��Hn{��3�@�.j����ʏ�����y�t2<5�0��&���bo]�E��V��Q1Q�q�z)51��8Q�x�����a�r ���KۿfH�[cM���m��[�A���!�m"�E��P���؃ ��̦��Ϥ��y=l0���.�|�ЇI�0.)1!�8�V�y�	9v#�h@3G+.� .���W�d5M;]p�\_L�$�l��h��)�Ϯ#��;sOtJ�ם�wt�=~�����z��rv�c�l!��lħj���eΛ��Җy�a;6��F��
��Z9�@�Dz��
4�
��:>�#��<Ri=�:;�d��-�sbI�p4�;�J8W���R*DXa�ؐ�J' �5F��ILr��0���.gg���g�C�X��4}i��J�����悮�O��� ��#p�f��ξ�ʏ���|��l�n'�My�q�=<
����V�t����d�cR}<&�����ap�ʤ;@׏S/�J�����u���¸�	��BԜ���1b�u֯��-qѸ����V��EQZӮyh'8��3�A�A$"����`�@<�&�����c޺çl]���w��
�-�YO�K�06,��)����Z���E�M�>�&�����$B\'��Fg���P{�����`4��l u���հ	�������I�9����WJ��0Z�4뜐��g��^�DM<����e�ЗŁ��xA݇�Fa��4���
O�Y�Y�D#��D$�X�����\��)tu;�mz1Og6m�������Z�
�^��.�Zzǋ'�˛�-�i{q�brk�r/�-�ȢN鮀C�9���l�"�5v<}�+X}lBȤ^�y9 �~2<��Av�Ü�mP�h�� 1����m�	g!-���RsKm�&&�,��ϩ,�h�[^��d�e�P,56�%ꪖ m4�%�5�y��@��~Hr����Ó�?��G�	�]Ј:j���4&*�M!!��#q�D{W�~'���1��#��../�����$���u\�"=������  iK���������g��;]ډ��H(�I�Y&M%>�� 8����ltV�/���%&|�	�
�Gu��)۾��*���\��ܖݑ+Nj��ќnSw��'<���i��c�-��΢`]���>��,�+�.]����wQ���'��nM��F�AVX4������#�O�j��'f=2G��Y�)H���jf���g�N��|9�T��:t�4��!��w�ڣ	§�P�dy��)"�X~�dM{��\B+�焓{NC}ƏDt_ӷ��ih��(x<��z�H-�xx@(��ff	�x�
�u�KCI\J��"~do^ p��L�T�����P���i5Zt��[�I�6��hH9�e���OM��Aݢ��oy���J'#�-ު�l3��|t�1C��K��;�F��4����J�)]t�}r��|͕�봜�`\��нd�Ӊ�F�����q<�n=%��s�)���&��l1H5݀Sc��D��`���Z���W�/	M���ꂰ��!]\D�=�)���'qFbMS��l2��O@p/�;㽬��g�1��o��4�­�@��z��2YuU/g0%��yq�є�\��{*6�[+1�60���'H��8����v��������~R���Fc2���������2 ���%�%���V�!&6�.�?��ώn�����'{��ă����@���i!��F�gyҹ~������TZ��?[�!��{�>H(`��[��xO P��pc�e7��+��Uc���1��蛇,�^f=v3�<x��Z�N��5x5��`9��/��b)l����V_��7S������,W��$�<�������B���-/[�9:G�I��~�qBc��&P��c��++�B=X)�0;�y�"l�0͉�w@��a�)��)~M���zjje�
|���K�+_J5�3�9C��~E�;Љ�s4��8;�����ܚ������z����/%V(:�}���k�fZ�6�x�$Euunrc��JE�U-��$��\���-����b���D&*�-9o-'J<R]��~�Q,�������{����פ~o���H4���ź�eT� ��Xk=��r�U�^3���죂;�ݸ�#]d�}p�����F�r��֘3ߟY�󸾲傗M�H�NwWy�O�>}��I�?�?~� u%���2�^��/&�����I9��cT��D����^A�i��eK���Oop�^�*�4}g�~^D�%q0]��&F���+���|�tX��L�Sr�Zo�ż�;��!���{�{���s�(�2s���yŧ�ic�p���=�#��5T'��Ն���0x���YW:����酊�E@�J�N�y�.��S��ӌga�d��桢�c����'�/Ȩhh�@[���G|Y����c�	/��>\����+4z��]��:I�n��'��Wr^Up������(��1Ye���s3�G���n��	�no֗^ۊ���)�h|M݇Qd��cл�)O�BP*%�T�a�r�x�=o�&�K�M�Mkй�� �[=5�d��F�^�q���W��@i��J�p�L�4I�-6D�a�.���e�ڎ����6�}�Y�TE���~�� Z!�m9��z��fQa�l����q6��Yw ���qJ�<��t�/�q8E����x��@jÙ��8==%ɂ|1��6-[�w뺔���i����Ol�K����9#6TXH@m7���dEW�S�P�������d)��B��PU��\h����v�0�=�Ӟ��W�V��h����m���ǩ��w�F�[T�0YY*�D���'G����P=a�|'�~!�-s�Q���Niw�o�
L붋�~�ƽ�؞Й5Z��������,�[��������}	�:i),B@�*�KM	0����y�0�F²mi��AB����0�O�}$ox.���М��5N	��. ���>�����l`3)�2I*#i2�*`+�el8�|��5�ǂ�w𚮑!�=�������*����7��F�ط$��(6���P֖ؖ�;�����(�2�?zz�n!��#��vF�h��?;B�N�u8�c|���3����T>�]�YQ�j:o�"�bY�3���=ѐ�4�x~]����*l�7����&E˫q��:зO(�nB+��\fx�׹�8����u�q�q��l��� �.���Wg�<�ɓ)��Mi�ݓ�k[n�q�G67kWT/sN�<��mCK�浟 ٵmRlp �|\|�Ҿ��$Zp5�$`�P'0α�����4T�:�:�'uI�Ŭ�B�2ŷ"�Q"4<\Z���]�@�g/M�a�'܆����+��8��ASIT�����9�,
�7j�偫Z�]cxk���"����жS��*�;g^�����=�;���7<�A����",�0=�sy.s&	Ӻ������,�L0qN��:��"�	�B���r$�㽲����D�<�%Z��f5z���"R�� �]Y�T�u�ǬIz*��S}���I�[�5	��*�>�2<@AI�2'��(K���<�R��=�ӺDǭ�tT,\�\0���v�L���h,tm��ܵ�Y�:��+�ș���n�t���;FCPˠ���coF])f=����!�:"0b����(2p��d�\����荵\wf��5�z�Jn�7�������d���6�z��e5A,�O+Y���]�܈[�b1�v�Z�zK"�N�u��a�=���f�"�ĘY�w�?��8j��73��4H�u��'�$�=�5�v�op���Jb��}B����~�)�&5^�c�TГ(v��t�����O�9Y,'Z�b��+l�d���3H��"���Bp��dR��X/ӌ0���N�aעv}m.�JV�ic`��x6�~��,B�XxB�~��t`ɜm���&�H��{���K��l�$��4����"ս�]����R7t�]]��y��]��ߜ�H9��;}Њ��#���X��>�ҿ�W��2`}ucܚΑ���l�8�-���|��N�4F�X鐆y&��qYE�{�S�'Q�X��=Ġc�@�����C9&���ءU������Ŷ�?�u�̢`�B\��Iԓ����s!�^2�_>� ��,I�I��
R\�Ș�3�&(.Z.�}��k$^%(U���]�?&z0�
	v5���p���tX�������N���&���BJ�R��5h������"~%% �KX�����w[۫�If�J|�Am:�I��x�!IV��x�Z�fQ� ��3�w�m\|���[�*[������p�u>+�<l;9������T0Ƹ��NVm�Lѩ��H�o����܁�=3�D6�N閿�C(��4�A�`*Pj��a���=̶p4_c����Le?�q4%8R��~�����j{�o�ڡ�fq���DfZ��kp�r���<�1��C̿[}O�� �S�P��ɐۇ9\���l���o����R\��d��;a�z�h`�QF�� G��=�ܧ��z��B�	E��[<�~�/hE�(+���5e�7-���<��;T�/ܲ�%uD��m��[���
�4z��?'3u�/�{�
�bC;��w�I�=�lz�2��B񳁳�P`ώSΌ�L$Q���Bg�TR�TV��j�S�*��bx�nb�	�����!��<(�ƹ�r9n	��3���mZ�|��c7㪦
�O���d���o��5�͊�3H ;Ր��d�#�i�½�1��@���<x�yI������Q9�`�
�"�� $��θz��5�3���T��>�'�|�z��+~�Z���>�;�H�W�3�Wx&D	�o�&�S�x)�~�@��00:Y�t��P���90�n������T���ɝ-u9�Ƌ�
7�:�z�J�-���b�.�TI��搢/+����e�͋|��Vs��9�>��a&�j��Ys")�����]if�Mڡ���:/c�<���l�Z���/YBi�d�Pve@��|�u����f��R��W���c)�m���g�Iy�9��/p��$���m�ď)oa['�=N!]���/Ϣ�5Z��:��e[��>��;X+�C���&G������UbW2a��9���O�X���P�[CR���!EQ�E�ʨ�O�,+�Y��x�\���mh+̢*�΂�wk�F�ǩ𥥑��"��Q��*W9���d�no1
����=��u/�g��&u��Е[tۡa��+C��̦��O,��(�st��s�����= �F�hY�V� �_����'6��l�V��]����G��dH^Kk'�=f��nP���1���o{�\SH՗I�_���p�þ�uҹ֙��^��Oͨ��N�zYZ_�]I��M�*�Xz�^f߁b��ƴ9;>���F�P����
"MbVc��1/�� .�}~*C��d��b�Ba\ÔR.�I��ͣ�����p狘�wWA�Uo����?T՟�ч�n���U(@N�PU;��&&ǘw�2�Z���:Q�r�)��@<��ϽϘZJh�7��:7o�n<��n��Kk^e�iU¹����}|�g��3�ºk�O3$Ap&6���f����qM��^6cն��!G��̭��ձ���y���y�>
�����U���� �Y�`]��l`���[pq+�s�a�r5�2["Px̞-#��Q@���3��R�������}�w��y@ͭ�18��.����v�h���m��K/8yd������=�tcz�3<��BT��	^��&\�	\%(	�������g����ҙ��3�.��E[R��
�z�\]���C��Vk��?�B�<^`�����oE��G:L����]���t���Y���d�O3����m�k$�H	ф�{�'���k��������o��ol��6_���;�=x����mt�՗�����9U������kWB}���'��H��qk�$���@�]�]CQ�D��M�h̦���T�j�O˂ζ�:Y��|�9���0�F������[�	�譞D�C�F��c��ғ��0`�o'��n�uM���-Xմ��f����~���iO����p�������v	?J3��l&*1��.���rX�>I��қ��^̐TP���V|kN%[������;�O�����VM�B�-6��.%�;9����(US�7��&J��K�>C��0 ^��SɅ4�-)d51윷�sn�
�K�6MF����p�j0G[����f��8���*ӥEg56c������y>]�Yn�W��Lo� �(��`�'��B�4����Kyr��]����:��c'�g��pM̛��