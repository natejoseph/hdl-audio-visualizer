��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O������.�C�zWݽK�#���V\���?`Lr�M��*��'����,N`�Դ���w��<۹��B@�1�'5\\�^�w��L��9�x��ڨ�g`UN}�E�e��sb��J�x� �%X��p���G�CT=��#�0EŁ�������y�,6�����|Λ��AJ^Z��]���~�=��-�۠�K=��sj��Q��EtWDA���8Yh0*	�J��@`#&D�WD��R�-������vJ��]���SL��UF�VY��9����i�B��A��tx�p�o6M�����;�j�32BK�(j )��c�w�j�.c>�;�Ż�W��;��f��m�p� ����%�5��� ���L����.(�Y·���&������+4M���k-!���m,6q#���o�;�dB�)0��)�K�>�����+���i���'2B���G�ھ?�R�ho��.
��7(0��.���.e�cj�'�c
�'i��z,��bT�
]�Ӫ�ޏE�ｦE@%��^�Ƣ�
b��fl��4�9ȥK�f7�/�QPe�ϴjE��),�D��	�)�KՒ��C�L��Hmٍ6O9�Xw�f�G����1�:��[2�H���6%*`ek���r��~�'�;�S��UhQ���]*>���4��Ĵ�L�����fR> VT���(���������+J��I+�'MD"ģ�dC?�e�IC�''h�:p���
:���v��;��G�A5?
ſ.PfV��E{.3�E�ސ�ΐ�C_��*�O��Ch5X���Ì-����4̗o��Fs�MgAz�����.��h��G�M6��L�G�es�g�o)k���\�=�o���?^4�-),�x4�E�.�@�����'���:Г�5�qerKN�_U)/3����6��Y��3�x*g!i����6����G"|��ޞ%�x��kn�â�Zl'?�����#��/����}����,/Q�s�z~(�e�Qq�E�heh|[u��_�[�޼w;g�2Z�=B95��*)c�ԭGE"���Q�j��"�˼���	N#�c�vf�n!4>�d��;W�aЁ�k?4(�o:��- ݮ7��k�ϯH�?1�;S�5+����ܫa��m�~��Ā����*M ȷ��DuY��A�_�#2ߤE��;am0R�@<���.Wu>�]AG��D�s:��g��G���ZbT`� r���O����H�;7W�(2�Ӆ,#|���KGc�˗H4��x����4zO���ҖKb�^��W��-���t�4�A�K��E���n4��ξ��黎m��?��r��%O
�x���$$�����h�cևC�s�xھC
�Ȉ��O�~J3�7�@�!h��܏��V�m�<
p9�7�G��DD���}�/Tb��\T�t�/��E��R��F�+�� ��hS�2y3�츢������e�d��@\N�����F��}`��I��]��l�Jq6����D(�|rH}m�St�����O���w�Q�=��i�ŞX�n�0�^}D�eB����V>�ujh�"�<үn��jϢ��gj�-�Q�cSw��� 6��#���j���>��ǳJ���MTOfJ�)B/Eۑ�4�k�����\��x+� ��)���d��Q�<��R��9���`�p�!wr0"�1�_����)�xFB��+�{F0i�	�)�z�[d�=��� �l9^e�]�&n��%�^�����q��y/��#��X�~.�_�G��s6��{W2X$E*�cI�����P�Q&)B�t���5`~GF]��K9:O� q+& Ln�W'���	�1�quvz�^�y/��[s���"
�˵��p�d�8��b.I����i�ـ�I8f���i(�>=ۇ�����5@�Ό^%�� )��R�	��g�Eاdy�>������߽��@�=�2�H�X�ݛ���	�
�t�ef�ڔ)5A@��J�<�.��s�uߝQ�]Q6.�Z A.F����_Bt�g�)\Z���)�m�'+��Xu[��&]����N y���f����@�Ų��,���m��o|(4}�z�z5�gc����'��;H&��E�w?�����ۂ\@`���lz!
Ka�I�R
������9b8E�-���>6J�����a��9�2
q��.7x[�ky��$^d-�j����4���K�
j�uY�%�5⟞�-�L(���B���f����(v�\�o?�)7�$]��'U$"���I���#���[A����2��.Rgz�Q�	}
UI��]L����L����.�<��5l'-#fD�4ǩa-c3ϰ\�����c�C�jB�
Y��k6 � ж�8UC�5Cf�N�K��%�+�{�߳�4P�1��fn�2�ZQ���0�=Ւ5`��S��rE[��oM�h-K"��4���REb3l�
s��t��<��H�8�`�� �;�jʩ�������8��/#���]6NCU4��n�Ez*�5�~'>��sWn����o6ޢF��E]�ⷁV$�A�����ِ�IUr���ٔ���e�Í�8�2��Is1�(^��Hy~�H跲Z�L�ղ1�лW�,�W\j�ݦ�Q
|�*~$J��-KQ}�Rw�#Is�LJNف��G#F$�'����b�OAн�O�k�{����9Tƶ����0yŽc/88��w/SQ5��J&��Li��^Yޠ���
ػ�U&O}��3eͤi�H��
7Ьs��A̥�b���ݓ�ļ�B��~V��w�\]_�V7�ٶ�!����p��+�^��Õz�s.��?!�i��k���G�=���ybY_Q�)#�]I�_��;��_�q�F���u���a���Z���y������;����#3M�$k
�y������kѳ$�(��E1��8h���A��YY#�[<�^�h�jXG-��9u�L�<��2����� ��#x��3],�|}��)�/wDF@���g��h_�4q�����A�`Ӌ��ol���_���K�\���#���I\m���?�x�(ʦ�qfEÛ���^����h:k��>}\g�vS̔ `�E�$�����h�= �^�e#��{#�+_�E���!!�ƬIRcu9u�=�fXY	Zf�������-sB���ǂ��T�ۤv��ɻ��-�cQ���]ģn�C���
���_i:P���N:�r�^��Z�R�o0�}�b0x7��m_R��ꖣ��@�'>D(�|5�}���Ƃ��J�Uh����]$t;�%�Rg�E=6'�N��e���`5y�0�f��!�g����aXp�P�*>:e�&\�=����{GA�es(l'��0�G���9Q>�2�y���d�Mfa3d	�*�_�L� �D�Y�Ӳ'��	�Jl{4\zPT�[���5~'�z�s�q������Ii:��fc�@�R��	��7��ۗ�C���)����fl�ps�����[�۫-Q�[ST|�R3�؂DO�綒6Z�rk�B����M6mf�}��}�݁�J"afݟ}�S�/
Y4 ͨ��o�$�͕`i�hy6ҡ���?<U�hP݋�>w��)b�Y1C��CS�3��zC���w�����:��ɍ׃�W;yK�&��(���I��C\�y;�)�����������fO�K��Ɏ�K���ųόw�?�0����=db� \�q>Qħ�P�kҘ���wg�]ſ�s<����:��Y�1J�&o�>k�]�}�L�՞�$� G/Ɍ���B���mt�T*Øs�a�J� ��^�cnO�V�$���-��#�!~͝�5�`p:7��[�棔�ڈ�� �tH'��mW�����8&C���� ��U@HI���46�T%�}��mH�4�fk�l㦿��x�ޘ7�4��:d(Ȼ5 b�}�����Ux)5��CXm��o�5JD���M!�c����7���o�+jfA\��X5G��0���C���<�:[D��;���_v�[�>��n��񓰣�c��FU�z��}�֌]�����\�:���
�i12��m����y�?\t��5�`�"t�����I�eP�,/F�q{ڪ$� �b�G�f� �-[4����՗͏��?���0���X���w>4�K����
e��Ԟ��\{�0^>}r�[=���K
V/|{W�V�o���1C�f�� C XLm�	���z�������4�lC�͞Cj�z7K�Vb}�L8Y��?؆$���k�g	��'}�.rFá�C3|k�)����g�ױ�8W�K>?|$iUlM���qh����]T��,2ɐ�a[�Y5&�E�&��Z�E�6��6�2��O&����6�A����=�6�|�|��[�a�qXO![ؾ�uHj�*<����򾥴�#ǚԭ 8�ޡm5&��c<��<�G�2�M7��C2v��Еo�Xd:�����?���u���A�v��/�͍��P�ֻg�u��g+S�)��0htB�I��{0���B��p��k���m�K(#���	H����B�� APGUS�;m�~�zo��\)c�bj�H�y���SN���1|r��Y������p��*=�)�%ܶ,=�m^���ў�(���:�)6�dKͿ�M.n�^�;ta �6�-��޵%h~BX���A��}��U��@V�$7��J���&���v=J*��D��"-;�\�Z�Z�u��'8���k԰�g�����8��6sM��)'�2�$�!�OP����?�g�om\�����=Fe�M�O�0G�����]ج��?J����R~�(�s^(@(�<�`a}N��fN�J&�<UOo�!%��s�C;q	-���%�hT��X%m��Ay��)�|�o� �yx�L�����af������_�#��T$%_����l�F#���Kl��*;���4�c��^,�^u��O��K�k����@�b���φi�Һ�2���D*svS����$'ǟ�{ %��[3�����MB��b߻?��
�T��/J��ZϦ���<�-,�x/�j�[ʸ4��]ui�T*zS��7�b��[�v����U.���=�$�wV%�T�h>�۳AR�R2j����Գ�S�"����줓��7��<RU����Z��ІƹD�	�K!A����� T�*��E׆	���o#�vտ����$�؋�E����2ۍ����`Gn��".�������vg�I�[yj�����'�^����IF6��}h#�����ti̲��N���Oy����JQ�>k�:�h���@U��=�#��z�����b�|����]j��5 Z��AMw�\��l���s�@�P0z��X�4m�Q�;v]��"Y��G���dN��I�'��M��GD�h`��a��H�o���L�R�L/�s�u�O��Նئ��'k(mO'wHO�e�؄�Ec7����Y�.�{)��[�Ӡ�����4��x��v�v&��[���|2�x���X�K��ț�8�^\R���S@4z'������f��W\X9�&��w]�9�#������M?�3w�Xq��%��ڽ�~99>�;�S#���>ܨ���/&Ӹ������L��HG�ck��7�^��4~JI��Z\t�ң?��U���(B��i�/��?�r�s����Mi���ό�7��ϳ�-kx�꒸=P�-�jf��|��gv��"n�"���ۆ�-ܗ��Gr��FT�[t�-pn�-]l
�Z��?"q/�Ԥ�g�{<ڈz��8c�m�W�ì�<l)�ز ���k;�y�}��S�)T�A� Lk��[��P���o5�آh�Jk)#@BҲ�Xu�+��;��
������F�`��M�Do�Og^I���A;G~��@���vuTh[��,�[���l���r�����w� @�)uyƊ��ѫ�Et%tÒ�5�7$�$|��K�+5KV�T {��}���%������� 7���%��ſ�ݝ+0��0lE�ݲ��B��fWi9����z���,ר��Zκ���oAk�r魬�׊+�����d�^k�v�Yv�txe�^[�.�7Hq���:���7V0ܴߴ]���?�`��[$(�'M9y-6�j.~��^R4��zi�c�i�-1/`�����t�'����aQ�I�_�CG�e�jw�����;���|N���g9͏KO��?Dx�����0=Ю�S!�%F���OĎ� f�K8�CT�m�Bx=/����v���ü���9��vC��h���&�"C 7;��У9[��{�4-&mP��TL���*}�A�
u�[�[�@�~'��̹�Uio�8�Ĉ!��u�O�>�C�gf��+^-ZBı�Ѯi�s�p�1\WB�����*�F*I��ϲ����Q��^���Ƀ�~\`��
��C�h�%�G�C��jGF9EoBQ�J���;�U���@����j�9�m�jW#''/~����YED�b�y���Էz����m;�?R���!�h�V�%i�>�NO����{��
��TOd�f��K28���'�f�T�#ɱ�@S��	�8��H���Y�smg借5ȩ�d�K�����h-jɪt=T�EM��M�`�5:���G-;�;���U�+�M(��ܪ!�]>�u�5"�7���l�89����(�#O�iiL�8��8y�����R�����\��Y��G �~����Z�]�}N��k�)#KV��*Y�9�u�q�oh�*���NI�e�6,}�	��P)�*i�cT�LX��$����I1B���J�F�p�QV�i��*���쭅��p��|�-��}�5�b-$�yY
@Sr�
�Ný}g&���
'�>CR�7��I�l�cȞiH��@�t�u%�r]t%Qt���"i��/M���:�TO2#�*�V��	���u�kw�дGO(��q ʢΜ�襯\�>rՋU�9T�����R� �_���o(�x�Kjne4��f����3a]�گ ��J�qW��Bu3b`N���iAx��>�D-v�-;����4��^$5��M>ׯݒi�qs�NN�@`�Geg��!�9�k���`�q��~��7MXk��=��i����fa���`
m^>���!�4'ѿt���>S�B�����x�I}9�黐:Gj�ͣ��XK��n�|R	�WK�/۾��p��)�MȾ�XY��0n6��x����p/4T	��˞X�$b��/�*�1��<�9����Q��I��ɏ$t�LE���+5ڽn���c��%'�0j٢6!F��%4<�'�!�)���˟����5���0L��e��u�������Bz��t_}������a1�ߛ���k����)�tK����Sɏ0WM;l#�
�uMt�ɑ�Ĳ*��"�ҿkT?�,���,��FV����K	�=�B�I�m�JشR��W��M��ఐaϾ�
*���-NOQ������{rż����&�� OY�g��Hb�gYy̕��n�7D����SҚz��=!�#��f�灅�gNW(��L!�Bw̼��|D���Cѿ3�j ����wg�b:�g��U^�T���r�X����`e$��k|z�e�!͐�2�p�[�\�vD%쾑řj�_j@�A;�̯�����`'+c������-��Mi��+�w�WS.� h:�IA]��=����0�ߵ�Āa���Y�9��>V�`;���Y�<\�R�Y���uE�<^�UΦ��+��qr�?ip<] դ���,<���`ţ���J�Y�\M��M5M�2㰃�d�UW���<�[����ѯo�5�(�M|3FP2������Rߺ!���R�0��mwy�󥑛l��rq�]��6
�Y��M���B�/nygh��*��t<�˖�^���hC(��~��������q��; ,&�MAd	�B��p���X��&��0���6��=��.̗V�_��!�#UT7���<��"��7�-dwA��|a����J؃�,�>�A���Ӝ��EA�t�
��;�K�o����ژ-y�F��_���������m��Q�����cc���/�H�X$櫣��;�t�O���ԗ���罩)�<IKr{!D��g���Xo$���JxE20D����p�"{���h7\,��H���gU	�F��<띀�M]�&��h+6VDe��r�'>�V%�D��T��܈�C����X0��ѯGhU�L�#�����_�t�ܗk�Za����|�~ò!���|���89�|�B�M+�s���Qk'�\x��2f�ו��x	؞�Q>����Iڀ�ͩ�ƨw�tI?����'�v�q�U�F���9�Y�z������w��g�?Ļ}����^�fDG�Me���v�xN
����n�xI��V������@������>_=�׽�#�����K#p��!-7S��p�M
up�O�Q�y�}1d���[��;ܡCjMv!q���O�[����2�z�de���~,$=�����rJ������~�������-1,�X}��7��f�e,�y�<Fމ:|PݖH L	|���h�s��e��최�dX��~�ˈLMQ<+K��o�u��B1k�=[SN�GZ��ZX],�X�VS�$�D��O�V�c�g,V����S���	6r揖�5��`�4�7���2��}�Jb芬��#9�0�]�K���������c5����k��_LDI�;��Q���ff(K���RA�.��z2��iF=������B�)G�߯ɍ҄ 4u��G���d��P$%�M����������(�S�j��3�v|�t�H�w�yP��Ց�a�irD��t͘�?�*P�1誵��1sX�H��MYqvM�@�dX��X�@@�D��:���
���e�
:��E���rP�+�Z��QXs�R��m��Xt����<���m96'�B�,(��RǘZ-��t��ӻK�����f{�0J1��̻�~��/��,�G7E�*�p�0{��K�3@�����Pn9m�i�'���b�x`��c�3j��g�0�踓$"4� x�ǎ
�#|P���B��E�Fa�i#Z�4I��MQ�Q��n/2�&,f��GKB�M�Q� �Dp8Ga1/[E�ӝ�c�d�ǅ�� |��?8X��៟�@ެ��>�P�}s��gL��+�Q�����g��6'�_9�̼�OE�����^�����k.M�kP�����N'���d����v�ʵ�9]P��	%�68u�����c�	�|���t���F5���+z���26��L!|��ܐ(ҭ��Bhv�L^|>Oٖΰq���)ٛ���]�B�Z ��G}QU�K�S�� ?��*!-��
	��C=)|��k?s (T�t����\��](��Q [f��ݛ��0��.\u5�i��G�C�y�>PZ��Sf�U:���H���!>:hf��a�1TR�w���`�T�|��i�6� r?}�\+��:#&btJ����`�$4��y�V?�x���T�z�U57�d��}$�q���HZ"�I��0Sٰ흠(º�;�8c��}���VZ�� ���As����ʦ�y��Zа�0ސ�SY��i:w�35�RW�`�e:H�"C�ՔKp��$�L�N��� �W��������n�(�� �"9�!�	��Y����?Ń����ѱ��.�F����Ԯ��怶����~n��:�����	D�Jz�����7�lw(�-�%���R����s�Ѥ������E^�J�y�7��S9
g#�>���������{� �B���������r)ZKƝ|T��N#gKJ��������u�D<��|�&��\n�)u 3H 檚���r�R4?�6���Ī7®ۻ�oBz�1*��E�X:������qx��s���qz���=FE���pY�f�X
/���c3@�����{�)�-U���W����V�}�4��>��kM�P�s�,~��U�{l�Fo��F�S$ݤ�7	x������B��6�岯N��~1*߁�$~��:{������̯�}V�kZ�j��<���tZW��3���'&�j'�;�ɉ�iR�������YV$G)�Ot�W�:]�8���;�X��@U .2sY  ��o�%n
�>-`���ʮѯt�V7�F�x����v�����<U)���Âd_�Ը&�hug��#BpJ�A�$��p�tû�1!��V#���_�.�[�-��}UHTe1V���`��0_7d��y�N��"J��o������s�؀��7�TT������	W�א5N�6����}�BP�"�$�(���% �Mw@��R-.��h :קVC���j���P�ReD�5'4����˻��o_M����&*�|�H����st�M	�̨�%J,\iq��!�����V<�؁��.�,��}w0B��g�}�bDu�X���ݟ����^����]k�ޅ��lFg/��ȵ���4�m�﷒j3��] P�j\e�����Pzr��O��"d*���M����ػv\��[��Rf�z�nK��q��b�����3�C�̗EXe@�ѠS���(���G�=pHg��}� ���G��ɒ��vO[Q��U�J��+7ֹ�f}Q�ȿ���"	c�2J���/&��e��^^-8���@�V| 7���c$��Ei[����M�Ee�R������\�tJ��A�l:|H�E�0
z/���)9,ޞ����/�֣�~��`�G�������:�"������ҿ�P� '㕃!%�y67k��Qԭ	�M��~}X!�i+[�m����ٍ#�#���lK�GE��Wx�g7�W���F�ħ P��6c��J�6ɚ�&����R",L�Xd�;�)��ΰ���,���r�y]�HG�N�.ȇ_�x�-�j(w���GS��Jχ@H�o�Y����EŌ��A���=��uN7��zc�>X��yR��W�,��G+!���	��`�y0*�K����-fi�J��l�/sN�.�'{�ْk��Xu <{��m7D<ݹ��vِ�\,��ܥ��e��"������Ln
�!��%:WR` �]MD{�_���ѩ�ʲ:R�c7��!�W5b��#�:�U�5>$��ؗܮ���?�V��,��IO�N���p�$�X�R�u'7o���K�UT���Pt�����B{B'~}��7�7%���"�O�~����%�tq<�zb�*e�+F^j��G��Rw�\-��P՘����#�X�I�rʣ�յ����1<ߣ`j�wvf��^�r�U��B����R/��\ȇ�<e�|�2[��n(�Ě�<Ý]@�>7�zN��kH13���Y�~o�"\cn�|�qgCd�#�U��.a��|ׄ��x��־\j_+?�9�ej�����Ø�TӝT�=Oi�l���zV����H=l!��A�0�h���\�խ�$oQDk��iU���EF���3TV�|cX����:��>͖�D�=�����$)���(�g�Б�AG�b<�`;!���
H���)�����Fs�>� ���X�"%�{����jQ3�D��a���%�<�,�x��6����]k�i��p,���xE����и�*��G�Z%�����i|��t)e5�+�m����L����$B������ħ�q��f�f�}�ˊ�ې���,x_G�lu�/�X\��"�j>QX�;{�����C���q��H����4���0:-�G���$4T�U�w<������	�!s��]���F�jC��njg���&�qKi#�Ezc��-�5i�X	:����Rt����;�wc?��\<��!$mT7{���y�ڄ����5P��6C5���O?Մ�hp�U��>�JÇIL7!�a���Ȳ�8�W'��m3?\��nwCi�X�k����6�pF��{m���x�ߛ��7�;/&$ts��CK���\���C���s�5�N�1&�h.�f�pe�t�2��%ߘ^�^9-s�4�5�ز{�"L'$��>����� ~ؽ�4�8ݸu$$��9���$Q�� ���sR;�3?�c�
��.K���h����T�9�`�xQ��-���Z���K�f��=}�5I���Ž�m��CB�*	��}!W��\G@�<���$����}��U�sJ��CzvH:ه?b���/a.��J�[��w�7�zW;�40�(�q�����:@#�s71�(�m��o�?���2��ڒ����-��I��{E���K��p�)��UP��������2+�x��cPY��� S}z�|.������w�����3,G��)�Q:���	��'jm$�m�Y�9�F�u��5��u�FGu�cY�Y\�>DKt({Lkv�Iլ
=�umh�&���4qug�2�Z8U.�ې,�g(���G]<��܇��b�t�\:�|�rP8K�ͪ��5�7���m!0s�*^�ŜA�%XB;�l;�u����KT=�����;H"};�v��,�{���tsq.z+�9�����`��\Â�ىp�<���urG�@_�l��G���qo�w�-P[���Q�N�o��U�<Ǽ�8dG�6e�|�GJ�o�3o�it�mX�:��L/)��of��Y�b��
��t�ކ�a�F��W�Jx����]{�����miinzn�����)9���BJ�����Н�x?�_.�����1�%�3���$F@�s�x�	d|HF��57���x3R9�g�/�%��"=l�8T���1F���Ka�%� ar����8O���Sal���kE�LT��Jt��c��{KI�U�&����,=�%������}wm���M�H�3~F�C�9d1���_&�x��u�+�QD?�ʀC��Q�T��[o%�ߪ�G�b"�hyơ�N�R;���/�dp��~��%���pY_Y��P��Z��C�ݳt����/V5�x
o���&h��`a*4���{b����#sǵ���AV<@�t�R��	bq���)�N�4:�s�_j�iR^]f�k;���(e��vԚf��&��MX.7/v�{r�H��{ GC~:^*�b��e�*��7w�8����=|�.�+Z~�Е�s��ȳ2x���P^�K$l'ѭNO��Qp�0���`��?4t��dA$8\�f��!#93����%)��iIzd�L�"N��4E�%BP�	�1��%=z�ʧ�'��'�o�<*�YO���H��O�sC�2v���~���4��K}����������5�_��BDV�.�`+�c89�]�^���6�Xkې�8����k-�n�4��3��55*���"�:�H=5]�J�ԁ�m���iwwkyM,X����܎�)�X�S~Z.�,�箸�?�0fW*UsY���;%q�a��e��+���]����#����xi�e4�W���?�gP&�l�F3�X��O��q����Ͻ�mqZ��I ^}���«Y��z@H8e�(�ܬI�=���˶���5��;#��m�d�恚�ai��K��
��Z5 �>���OU�X7��,����f�>o��Y�Cj��3����<��=v����x�m�Y�=�3��͹Ho{�.����1����icm��[d1
!�E���ػͥ�2��
_2^�zΤh=<�o��V��Z��UB��7vut"7͈�H(hթ��$r=�B��&K�j1�qX1�.�T�0J��	����ĺ��>�r*�wMY�l޻&�mRm�&����;�����L�i��9��G�-�⨮϶k}�՞f�"X۽۸-��	
�04������;Y��-�F�q!WO�N��o*1��ϡc�b {����ޏ����s��.�=�jh�Ptr��w>���	���,�����3�3Zt[�u��{��Xs�`�^Eҽ�a��a�4�ɰE� �d��6�7-��6VY�> ����5��%�\�\�^��O���PY��$�H^9ȅ��Gxڈ�`�ɠޏҏf�Rn��S �M���E[���+j<aMA�� ��x��7 |Lh����	�e5Q]`��� H��~��n��פ�g����ن��.aA蠘�w	�p�(��nu>���|�A��61��6�I��*���M���܃T�B�����]Cd�`��֫���-����6U�ᖚ�#����쎈F\�f�G�_#�Qk|2��:��P�mʐl�8*����]Ղe��Kg 6ͫS�T���/462-��Fq�|>�Rl�\W��\�KQ���*X�1=r�^My��'K�8�+�|��k֏Xu���Dڲ��B��iM�ox��&��n���F�y��C%�~��k�w���<��o?En�[�s���f�^���b�w��q�'φ���Y�˒�q�Iqs<��y�د��*����H��+NS������=ȲK����XV�D�F�� O��=k$�B�%���P2��!�<�\֙Fڒ�%�u,_��srl�K#� (��E:vT���`݀L���I��q�i��|�ˤU�w�u�ĵ�qf�W���Zkx�f���"�CcHu2ʁa��܁�F(��b$D��X���{\�H?鳉�%�����ҵe�D]������ƆPQ�׌��]p��lE�N��rW��qP��x��rW�́{�;����R�$��;Ex��n�g������M��\����*�gR;/胻5��
2u�����Mt�o�_��	��7�˸!{uB.MY���d3��~�'����S=��c��d6�"�7�{�3Z�t�2���{��+Y(��3=����=*���~}���oi[�V4�pM\{ń6 �C��r��IFro[�ȓ�S�
+�f~%J.��6�yܹJخ�[�z
��-/F^E=�m�x����~��s�F�;.ۇ�e��x�+�����ߪmА����r,s��xd?I[0M$9AP�c�C���X>� riCůd!c��h2�~6�/�%�����ڰ����]�E'� ���W���t�H�]��������v��u!g-9A��^��J���Q7�v�������ث�b�'�v�����'�b	&r�����$���S�����#�]m+��膏�x��D&���{�ң1bV�Z�ڀ���Z�!mr�������Z�M��l<�v�މ7n7�+��:��"v��Aڇ�� ��E�}��7�+���MߢP��0}�t�1��9^3KB�W�6�R������_ɲ���jC஭�~�\�Z�T���ȋT���v~y0J{7Q<��i
�7.!���D���ݽzFDL�D��a�`<�z�XCx����D/����܍��\ASc��CG��BZa%nYv_&�ǆ����1�*T<�����=�r1��@�
j-��8��&uA}�D����$z�^Ff�?Na� ��:Ÿ��\S&��Y� �Π��p����<�V�c;L��$��Ԓ^�N�e����;$tu�&�R���L֤�[���ib'Vx|{�0�/��f��g��?�]6��C,0��&M����|S����}x�ݎ�Hۤ��}�]"�n��7?r�4�q?�U�\i�	�ݔ�|�Q����?�{c�d7�=�#iM����-�}<{�A�[�����/�e�F ����%��j5� �o�����]t����oGl�`s�&��6�n���V}��kS×���������ļ���nl0��I�VO���4 �:�7ݛb��M�L�Ep�$;I0��&�7�*� ����%	P|仄Ԁ�l	w|q�>6���}�}.�q4�Dd��p��袶�-�j!�Vkav��V����:��̂���� Gޤ ���+#/�(���פS��ِ��'�"�Iw/1UTaHq,�P��k�!?Y���N���j�