��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��"涏K}���&��$��f�gp3˅�E!J��(�gB�p[���me���\tgg���}5^���p�[��J��0�lϨJQ:KH֛v�~P�e���*���}s�$h�ƺ7������G�`=÷�`�"��o5Y����yTs��6J��XGir5�>狯�mJIq���29��P����m$ɴ:��<P�k{~�Oa�^Yr8��Lv
�C��3�2S,Y֐�� ��BJ�~o�)A�j �<�>�����6O}�sT�C��-�\:)^��37Zʪ<�}��^������5��o���R�.y�B�	�
��~|����v5g9�N��h����
�I(�x!�A����δ!� ��,�-w"EVyr�q-��HO6��?T��~�z{^�\�oD	how����q��^2n�{��#�0�#.�?�
��T�,o���J�v��I��U9�ϫ\p�ffC�)'oo1ϡN��,@F�{��es������).�XaàԪU�\��3��R�67�{\���`WzDz�G����t)�������� :����#�FJ��_"T��2E8����Xk������Ht�4U�`��o>�,�Z<�wި��3ه��Rb"�BE�y�i�/����Ξ�h���)��P;������#�^j�o�)A�c|ҥ���(hM<
/p����NV3�
Bk��M)�d����[�ȀN)�\���eϖ�����e�"�N;�/6�O�%k'���C��6��N�73��βځ@����|�,���W�������d_aH�/��V�&T�asz�����j��s�Py��ᰛ�{7�yan���'��/q
�2�_����u�IR����q��~i)]��WctM�%ݘW��p�J���p�E��s�V�Kь|Q2'�0������᥶�sP�j,��g��K�f�D�Q�J��X���3˹k4�nY�2�
�a݋�jW��;���#
����QR��($�ں�p�8OҊ�`d�?�{3q��
!<Ѹ�~���U�@�����_�P�QUoå>Mdfgq!>�t����G���Z91�^z��B=�L�3�%3���y�~.b�k��CX���a��ξy�	���t�9�n��;b�g����`K�>2������S�s��2��cw�{��=h����0o�͌���Q�g>��"���6PY�K�ߏ;��шoQ��	h��R�;�u��#�9�񢊂�d�ikF���j�[�m���&{8ő�2�E��uG$�,��!���Jy"�ݾ��u=A�8���):�i�խA�@�u��(2О��?�@�Y�����C�ű����9�lzE��MD�O:��� >��ok7N�gm����ٌ^��nrP���nz0�1M͑W�cq0��������!��<���v�B��n	�Ǣt��@ı�:�n��Ǉl}����o��w-<��-�/�����;�@i���>�s�?����y ׻�ۚ# +�����|�������6|<����ܶ8��z�+٩��a�@L�;����!�#�r�pT`�*���(�n�%�yZ�1��q\�ޯ�r���K�*ljS:ww��^.&��]ï�A@ς�`h���Ϳw��z��k���pH�;��}��p(�?q6��� 7���5������?�2��>`a8���Td�|������Ir�+��(^B�������0�l.͹zN�I���8�Ѿ>�e�@�ĸ���%�����^� �S��et�q~���JX�~x�����@���6��X�'�H�[7�C>��s��ybL���p)"N%�jJ�\9�Є��w����K�5[-�����r�4g����6���E#θ/+��7D�k�Gw�!d\ <囧=Ol�艕l�+����a�7��dBD�#Թ��ժS'�o�=���0|O�"Y�r��V-�p�uڊ�� ��5�J���iV+��w�K*�N�lJ�A]�'XY9�� ��X�B�ã�� k`�
��6>�{H�s?4��#�G�O.�}��-�\�?��q����-A���N�70RE�@��$���G��x��ɥ�-ԨH�ORM(��3(1�za�Q�j%�`�<)��!��j�S5
��a{�M���"x$h/92�
�Ҿ��DE�x��_W�%�d:Ǎh+o�N�w�n��0������tǝ�; .�V���.�,y�w	?��_�P�q3���?�4o�Y<S��:�j�Ϧ£YƵ[�I`s���ߧ�wfh�"q�����}��mWF4������\��7v6;��B��nUMe0!o�͑�Ƨv��M�D�M,�I�=��r��js�M�e+�TC���M������&'���4,�O+�x�&=�/t��3߼>9�o&�ڴb�~�z�E�b��KGc�[;ҙ�I�rкQ�om	y����$mߚa���4`�4����������t���d]���~.귵0:c'����H��V�{b�m%V�:cӚ��
��:�/��T��s�k~��E��2}
��ũ�����X�'�X�K�iO��cR��U�-��8,l6;�_�WM��)��.G`s/{!^��Td��XV^?2w:�4jL�g�E�\���MUm�̂z�og=�������$�֎�-!I���|jܰ��p�f��>&_U�}��$��ԁ��JTWx���I�þ��3)b����:B���[l�z��=�/w"'av�b[������U�n���(LZ�0}Xg2�8��
�-W��2�Ɓp�"<�'v|��0�
N�@�fu�2�� �|i� �o�1󔲢��+`�rq�H��>���̀u;��1.�8��%'ՔKl��	݋)d��Z럵- 4v�Bl����</�f���}+Q�_��g�����&����T�1h]��e��/�c}ˤ�z�<M<�iB>*Ҟ��6ot����t�|���Q\?��F�CZ�����~����tny'�Q�J�j��­n�O\��4�إ�� �tܖ�^���׀�[y�|�G�l꽌��WM$���wƷ2���	͋K��-�#o�iA/����j�M$��8��+�})w��\��|DۡE����$�`�jՖ�`�9^�t�T��G�T�\�?,4D�b:����w_m�?+��Q���
�4B6S4��l�e׆�a6����/�R�O�/S��-I��C�T��CNO.?)�X!�u0�%�vc�wQAR��nys.��M��U�Q�l8R4r����=s��X��P����^O�{�CHp��ؽ�mun���}�$/�9������I*���e\r�9rԌ���h��	`�����i����a@����z����݆�������ua��/f:�(���/�n��P�]U��ذ�u9��Q�������5�kZ���냾�k�(��S��x���8�5���J)p,$�goz%SF�ѐ��:�,ݭĈ���h�?ћ�(�%sO�\�ab���K:� ��BV�a�o�>ChĬˏX�U�����:�K+�����%dW�T��-�3\��w�2_E\zj���?$�,D�1)�\���R���R�8/P�������%�C��8������Y�\���%��������!��4B�L�KmL����gL�|xk;s6��S
�s�X���6c���O7#�+��/V��?�:ϓ��@�@�T��Y�L6��`��sڶ�����w��V�M��م��T�6���e���
�h ]�8r�{"�@�mV��?FP�Y��;F��`\�	J_�=n)��*�)/�W}[���n󿰮&N�"\�(��.���_��$�(��\tE-�O�b�XX�
�,%�u����Z�Й��!U!�՟�h� ܀o���r&�Q�ǽ���\���C\"�!���VsP1�E}��ݶ�!O�VH��9�H��	]� �	1�9PU�����k1s�o�I����.�G�ٛ�5��ު܄��B
��b�0D8�G�^��h��_V�b�w�ga�2�O�daF��o�����dcpb�;��Y�l]�23��7����q6��x�B;H�s������OO���D���|��	7��!�w2<�h�����t+U����3�iԯiV8�4'?�(8K�l�Ȣ�w�Q���.�'��0��9Y�|����hP�B�>I�h�5�"� ͷ�����	���t5�5�P%�I�P�[0@�j ��D.�����>�Z9RG��h�TO�uǀ�
�������'By��ih{�������O-�|_�;�S8��� ��P���G0��N?=�)�g_#Y�5��X��6e�.5��[ѥFe��j���o���ٷ>a��Ld��%:V�(���!�8�U~',��FS��dz���p�~�sSt��g6kt��FT��%T��?4�W�8���̮^�/I���,����D��ڒd5ڱ̆����h�\o&8�Q��Z����LL���Y�\T}��B�^%.�+�u��I�䌴�!�k�!�[� m�f=��v�}�Y�?�ڸ������7�H?���[V<��)�d>3��Q+�qv������t{�uc	me��@C��JW���no	ax{z���9p/t[hh*�}�A��L�S�{����ǫ�>6(.����Z�ʥ�I�_CT��{��ror��n�p��)l�E-��eR��朡����d9�r��2M��� �%�벐��6`-�8�����S�����,�����]^��yOU��Ы��2��뤽�~�mhD�(C������Yk����!M���<Vv�~�`��f�8�Zs9;C&"E����ȡ��z(~���~�ϩ��o��S9H걟��a4dֹ�5~�R����bs ���r�Oh��%�?�#v ~�V,���᝭�q/�~�w��U#)ۉ�%	�% U��ǟ�\Y��Uت +�q�+��=e�]uV�dUQ>.���]�^�A@u������3�y��Y�:w鱸����	��Z����~�h�	���dզ��Y�� (�d��F(��m��QHf@����鄿D�4ʯ��X��ʐ��`H�ojei'��JA�%���qھ��8}��\\Qл�O�����E��	���a��o�YO҉2�jp)u3ৎ��!f���r�J�HM{]�a����� ��j�sB#���	������u�Ce���I�D�~RUsyad>���\�h����ִ��'�c�6r�\����a�'��[�wo��	r�8��M>���f>U5�IҺ�=�����-�KJ@j�P��������}��B'�����^}wh�nTd��EF�j�j�90��gm<���4��w~�N�[H��"��	�1n�3��\���X���]F]����a�,�*`yw1��0�(�=���Tz�^�8�-	5�:���ڭ���6,���3�<4:����D\����[J�(�<���.x�~��P����Ͽ����8 �d�2�Y1�Hq��ǡ�[��Xﮂ�,��H��r>;Ch�晻�~�dﺽ�x=����E��`��)̧�\� 8�@�9}���/�����s~���] L~�,�$�>���೙�����l��(x��_�!F��FN�M��<��TA�yi������l����%eF�V�ۻ��q�*�-C:�x�����4
.V�~R��Y�Y&U��8�ԊF��p���BJe3V��/�Rg��`�HN�9c�B�����jK�����ܵz��0�p�WJ!�P����399P����P��ߦS��!�:6�R?P������i�x#Ф$s%�E)����A��CE��83gYDj�����S\J��s����e}҈����C�lSP��&},�v`{�[g�1�9Q�|҉�������D���Fz��ۋ��%��g ��W�_+)g��kI�t¢5��,����=�7Z�!�
�칋��:ȶ�f��F����aԬ/
; Q��W�����}�8�z݈`K���c4�8�[�p���a�Z��&����e1�:��د�ފ����X
3�n%m�ڠ�Z�b�Bs� ��f��b���;"ϴF�|�]l{�L%���Ǿ���=RW�yy��b;z�sn�����~�t�2lњM�9>�X/R��������-�oj��.�& �颪iE���򛖶2P9����*L��7������o)�Ѹ �W&�L~�=I��&��q��}��c:I�%A� ��&�gjݝyO]���奲�h)�eB��\뷦4[��� L2�~�܍`�s�7XaI�ސ����b�� ѵI�:���N�����SN׸�4�#9��2�\k/h����
�������\ar�Sڋ��d�$4�{��2�&����dP}լ���zfj��>7��^����^����.O�&H�����js"I��N�dٌV"�J�R��iN5�-�SPk���%ER��.�:�`# s�_X�������i���Ӻ��?A��zl����b�䵷�(�J�wH�%�Z"�����J��Z�B)#v+7B��G�h79�^Y;��_��^�04l����0j���`uV�1�2H����Z.}?�i��ފ�M��ɗ��1���%���Y���~b���vz(uT$1�Nʎ]A��t�	����A3��(�c���c�Fӎ+��|��̩랫)���
���P&���y���{���;Gm�&qG�Zt�U� �	�,�ch��?�w	�[�:��g!g�ہ����Ç��~\h��;%���ѓ�Q���;�Px*W)R3
�K�S�E*��2���&��,�����E	x�-�O(��pL��p��`G�c��=�A^��b��R�L�Y�6i�a���dr���ە��V�64�}� NҺ��lT�h|O�3!��]��I�Ŕh�k��!|ܴ�sO�b(�\�~,.�d���;0�^@5�gOn��������뢸�,n��\���seDeEH{Bx������Qs2�J�`��&���MpP6��
8 ��t�u���%�p5�8^\^`X']�{�
���D��}i� v�`��_Zf<��%��2s���M�e>�٥�� ̼��^��2��`����y����q��\� ��W��5��ӛ{N�K(�ϤH��Ys��WZ�#I��x��z�hT��S��S��(}]�Rl�͟��Jr�K�Ρ;J�4�{"�4r.�����@z�=h���y�u���z,R�۔�m�h".*�"&WCr�y�1N�|]s��[�co ï��n1��a5��P�Q�_��e[V��&~��k\�%Aw��@#'[x��Ъ��֛S��\���Z�w�j��<�@5o(�H�#	`��4?�_��I͛�F�c��GSؾS���j�N\���Ƴ28��#�pź�6Zꭎ���@� ��O'�賙f�fO�rW<�E�Wl���h��J�L ����L���Ai�˶��0_�B��7�ٟE!�C	��x7Y�VY�Ԉ����34�T�/ZT'!W'��ڑA~�|0����Nޱ��������P�!����f���uʁ(��>�wA��;M1�Q
��"�;�%`!��9�򝥎�A�RdU�*��+e\	�0��y���V�r��|C��P���4dۮK�T��2 �r�HS��� 	�ݵ�&�T6_5'�c�`Q�����;�S��>׬��B5I&Ɖ<1�"D�Gf/�ȇ6׻e�/���6�3�z���v"�e�\S��c���ch.Z�ŭa�r���E�[�OK�����4��JkpO�6іEl�[����E'a�E����U6�Uz?*���~��㼻���Vh�g$�]���J[yo�{��T�j�؄������V��H.���5�.1��ǂRo���UP������9>�7
�Ԅ-����x[��ba_.��y�����@�PY�����P~���3f��@��O�~w_��#s6kl�S�XĆ����a�G���=��A�O.D�}��������0f�@oD�bn��;_��a%z�s�(Z#�ַ�r��8���mG���I�t��s7XeOyK^�!n�5?n�2���oKiTqb�P/IF�I=�Z [��(,[}5�M�-˞��_�2��F&��&�<�J<�)� >�w�ԧ�[0%���G��%��'�]�K���D酛i��ѡ_�,��p<ś; w#�0����u�U+\�D����7G���]V95ze��3�WM�Z(�Վ94#�Dԛζ�GXi�L�.�g����i��m�>n#��m�*�(,�vh\�r��'��@�nFx}�R��rƭJ\��[v��/Â"�P���`��7���/���哂�
r>̴�\4���x/ݯ��2���������*\����N�} U֛7F�W2 �V1(Kvr��^��+m}��D�1DK�yx�|�l%����78�7�Q'�Ќ��6��dg��0p���/ޭ�!��H!X����ST�a�v5m:҉����<,R��C>e�{.L.C��K�#�p��ط�؁$;�g#��_�����8�%�8A�l�E�����;�G�R�$��X���,�YL��C��7�m����?��Ux	JU�Pl�v��{�\��B\͈��{i>nf}��ۉ� ��vO��4���D8K�v���^�E�V�
�(�-l�Ī�w��3
+ �9��	�sK��^��Ȥah�9 ��A;9v�yb�B���M��o�v�຿H��V���/	���Ҿ��G����s�E���5:'�d��9i��Wq&2�d+��(�ǎ�1S�@P��g�����Y~��>�B����;��� �T�c"�������;%