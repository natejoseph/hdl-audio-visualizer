��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����uc�1��x�ak����L�z�~nz���*3و%�H����p(��y��A\�G�b�����@t�/ϣ�*�!����g�3�Y{�ccO7G�M�����Yعm�*<v��.$������,m.U?q�v'M���_�섔���-�z��آ�� �`
�-S�*�b��^��uPD�UW_dH� �yՉ���	�n]����5��i�2��-I}-��Czz����Q�ЕM�@c���J�^?bc�ׄz8z�xWp�&�k^�����O��m�?��G�����ɰ2�q6m�X� �W�x=��9'v���}�����į�ߚ:犡��0���tm#���V�5��Dw:>0
Q�܃�}��X,���D�����WM�����;���rz1N5^��st-ʚL(e�ʐ����6��#]Ё�H�@�<���{�c�%	�ུ�>&R�Mep o�f�G�Ϸ� ��A|�=6���2ѶP_��0G�<�H��� �T��l�:� :=5��w��o��h\HzGd�l�"�
�T��Ɔ�t3ҙ�c���H���(N	�j6�e����Ɏq��z��E�g"�Ζ:T����-��	�B!�5�i����`8��y�`�w��`J��O0DR�L+�WL�wQ�ǃ!�_����/xɟ��,&����	?��y���<w����/��h	��Y�Z
'��e�W'�1���dST�M��s��My�k��=�+�P�,�l�Cᯕ«�_�����������w�%:��~Ȭ���;94l��((���/GW���'��.��OA�pS�ϡDJ�,l֥�	3k��	da�δE�#�IFh�.�ap8�W�>�kڋ���A���C1TJ�#�R�m�����X<���ҡ��+�S�o�����:��u�f�d�����Ux�ؗ{F��-��d
��{r��>�g%aۆ9ԜЗQ����+9�CG�J
q��2l����������B��@#��y�:R�=�Y��pl���3��꾀��߿�����k
� ��D �� �����|���;�є5��<ř�0nR���̥=9�1�^�j�C���x��(J�B��߽�(˾ާ�̩�G���@AV��dNaI�ID'N�0�73
���ؕ��~��NR�f�*78��U*�RŢ��F�׮�fC�����;�[}���؄3�w;D�J��L�J������؄Q����� �K)�llſ2�W���X}	׷~�1I[6���������^����%y���<l���M���S ���pі�:�c�Ak��n\xI��;��{���sU���+���#���<� ��,7�EC͑���?�����4�(����$�VJ�iOG��� R^d_��B�Е��rY���G���4o�����
Mm5^ںl���jϺ�_�)�ڏ���2(ʒ{V�
{|z�Q�j!
��d�dv��x�@�������+纓��sdd#�7��Aػ�O��(4ڀ~��G��DRG���{H��#2�9m�S��y7W�{w�=S-��!v���Y����3j��3��a,'��y�<,�N�O^�U�N6�	�1nM�
���=<��
 � �dl�L�~�PI�;Y�����_��*=��&G�;L��� t�<���:|	��֣"� %2Vvsı���-SL�
TL�:���J���*R��O��w(l���]���3+��HKgP� �@�e{�Q�X����j9t�]���F�Q��;n�a�#CeT��՝�����hHN3+U�m�S�nS�^oTq�uP1�����!��[Jl6�x{İ��6�Yܻts?��i�GC�v�c���E�+��C�����K�H]\���m�_]�!�43���bE�z�Pf���Ě�R��]����dFT�7S B���8^x�{N��߽�|�y��LlFDD��g-zɩ��V���⩬0=q�+ʷ;�"����|B\3��Pn�����B"��� ԩ�4p�J`��ln򍴎���oyDm��{Q(8�N��%)������Eޭd0��^���(�W�"Ej��m����ӟ���Q,7�Uۊ7/a4'�r�sl�Z�H�1|����^q U����[0�T�O����e+qT�FB��
��ӈ��>A%�:��&(�9���>�����O�[�v$��IR�G$�({��M�2�.�����:��1���)��$`r��bʌ�B��j'�c.؉?�rWqfk��#:��A������k�󩄾�3����9/ s�`k�:)ζP�`�z�dw����_�m0t�3ޯ�5;�3Е��?���)�oI^�� �#�Qѐ��NS���{٬<�����06�?�N�R����l{L�5���a���շ��"R��� qr����5�Fl�":�K���³y�+��s=2ݟl��4�?�����&�"�S:��"@�������&&`]զ������:k2p�uA��`�u#ӵt?!���H��Ka�P���q�%y�W�fI�(WJ��?j�E�(���ƃa�.��V����Dn�.4���?�ҋP��1�PNB��)!\�W�V[2l�/3	�!��A�ph��S�e��<�#�᪨��=�e5���Uw}EF����@P�G�C��ω���S+4?��x�r�y^$�>̎P.p��\�|-�G�#��2+kᘇ|e
_3L�oAg�V�<��O���ы�mv�<ěL#Ԭ�[$;����m�Ӿ���ej� �,����=!algS����$���xLm��P�[�"�́�B��W��. �i�42V8���+|?�=����XS�̓	xvRp�pX���
\��kC�K�3���Ʀ����ʠ��R�A��(�'h(,�Cֈ?�A��*$�8<�����C����l��'7��)��j%&�d)��7�e~6E}���|D�30ҡ���D����P}"Pr%�0����!�}ȼ�pGշ���ǎ(�Ə`-��f�b6�Y-��)��7�M��WU����Nꆌ%�I��8}A)I��iS�ʻ���>O� a
e�o�#5u!Kg=��h��%��WX�fV<�v6�'*�ܝh:BK�}���MZ��}u�3d�5��:�1X�w�p���y���������Txլl�mdD����-9}�2e��U�<��R��/��d�a��h,;﭂X"/b�j �4 �X�S�E�]���e���OcX�ͩnG�k�:�����t��fWd PDǇsNB�o�\7>���['0�n}L/�!- R_�Q;U�]�\pR����<h{�|"��r��Z���R<!��(u{J��E���<�C��Yc��䪙~�!ٍ��bj��Y����yO��B�9h'���CS?���x$�6�/@�#���\�h�T��E����ky2�v��Y�>*=Dpy�mcS�B[�QC���<�B�����mJ��.:��Y�R�)�
&��cv����c�e/*��̇Xуqޟy@�*@��u�Z�����-��I0�QrtJ�V>8��X]�W`i�3l�,� //��}Y�1R|G�ٮ�O�v�cG��\f*�nm]{��1fܓx9��A���*�!������۲7��1����K����f�`�ӎ_� ��ӗ��p�ׁ��z�2�+�V���ր���X�ks�`�.^��)p��|�j��t���aꈳ��F��dܩ����[WL�������8!ش�mL���=4��m�/� M���/G���\��`��K�t���&5��{��ߤ
��pf�o ��3���[�䐅�Qq'M#z�Tg|Ֆ���� �2(gg� �L�]���,�B�c<�$�l�ߢ��R7���1���O���$���
J_�N��e�&ş ���<\㾟�����/=��H5��ٟ-6x�x�:��Q\L591�������xP>
Ѷ���2���*����u6l��M�����lk���E�d��Ê�}����J�@���p:�g�r��qm�=Jb�&��E��H��V�[p���si~Ā�K6�h�[���t@F�,w���㶖kWW�t]b{3�O��70���yWW���j�J�9��w�e����*/�W'X�&25�}�������zP#<˰�.���%Ht�ǲ�y�9�ᣥ$�����F�`�/ ��wf���I4�Ք��x���/�'�q���y��Lh��4� ��̀����g=����!�Pk��]x�9�y�
zY� 2�]S����v�H;�6�`ә�8�6��p�$2�
�e��E=�;x�i���꥖���ؤ��	�V�'u�_Y��>����j�o~�ww?P�K��P,�b�sFaB5V�:~!z�[��zC� 0Z��X�ϯI��6�<i��C��X/���7j�����W�
�K(������g�����d�~���9!�f�ܖ����/k�No���M-q>��nͫ���O�-��^����U�dH? �*�Σտ�޺IyV, p&���=r��{y�Y�*���k&z�L2���;��w:��Q�7�Ԣ�d�[�G� ��'�M�%'�����z%~�8;��2�Bg��Ɣ���Xyo���_�3;���k�N{�+�P���V��9��'-5�i���%��cl�/
�O4�%d ?�XW2�9�)k,�h�#����>�Ŵ�_+Y�0��%چĳ%�o?)5�B�sN'�[B?[�ǐ�=Q�5�{�L�=t���t�@���V���8�ٓ]o)]�\E(NI?��NH�>�~w�}lpc�\V�k\Y>B`A�O.;��޲�Bs#�
�Tq�0Oz~��#�~r7����!���n�v��'PG2 qa^5��}n��}�j�7���y�����q;�Y�w���@M��n�*!���i���ޔ=u�	*5��
]. �v	�iƂk%�$�qY'�k���GXE���&��llX���ë�������tl��#�l��W��,��|�
�~	�k�s�AZ��h!�z�H�[9��+a
��%��wn���b��Ȫ	�a%�w�~J�)��&Rѫ�>>l�	?�C��9�Ъ�<�{CޗDtgΏj�K-)��rm�����B�/*S���'�N袸��J��
��������34��t�7��vI,�^���ӗ�S�Ic��7�O��q�UԜ��(ӂv!��x��@i�0j�ǋ���*u��FfT�>E-���K����Y��ЁYŃ�@KJ7Ns��O�;��C˼L>�=|�?�}EK%��&��L�ｑ��s�kt|��j4��	\4�6������<�
Mj��y�/R��!@��;a�jm62Wp��+���F��w��czF^j[�������e�S�>��~g�뱎�`[�cF M�{,���-ۃǣ�(�7�V�t���B�,x����f�a塨�5 ��Z�~h�b�y�s�k<���"�!�.ks�x���&�A��/�\������]N�*�[�o���'"�7q�脖7Z�3u�|��A�!mLJ ��
��?�܄�_P!O_?]�e�6��or�U�.�Iq����e*}���o]�^3U���e�@�&�As>�\�|��7 �P(���bׁRQ��R�W��=�Y���D�?��cb���}�S�fb��������M�
���CO�%�b���Q\����}���2���S��T9�p�N�m�x�G�'.���D�r�`@ݓ�_yY�3�l�)���=�9:��7�DB�:^�U4$��]�����iƌ�X�ĳ@iBb�<���*�\���*�=��65E
���f5:~s�%u\�	�7��Z=@�|��2q`kVT��e��vw3T޳�E�+Z� 7K��2�F.	���/��������P1��G��ᥩ��%��I&��8�;��'V�j���aԋ"���,�c�y�F�^`p���Y?�f�=��*%�8U|J~LV���G��V�":)Y��y���� �l���͇ftL��"��I�r�`BW��?i�r���m��G��q�ɛ��B������V��%�0#�AsG���u�g���P �ic�#�~��ٯɤ$�Q�5G���U=C�AR�S�*�Ї!������Ȑu��u����>�������D����L��g/�Z�q���*<��r��	��g/r洚�R��*� ���_�s���G�!d��fIP�[b��}1��e*9kW�mC�tpȘh%���aŨ�����b��|��*�6�S�j���r�=�s�\k���:!�Ɓ�ء��5����V�� ��g-�|����ۊ�A#-�6�6�� �Zz�c@:�rN�4��W�9����Z�s$Cṱ�i��,�8^�0��GY@t�d���t%���aC��>��U?�%d��Z��T%(Ɵp�P4\�T�i�M.�A��h�A�藫\9���\��^	�P�# VX�^"�#�F�i) vn\ܓ��r��m�b�{��K�P]O*/Qk�=��G̞��6A4b:�nC����^�FE���@�����#�M�^�4��A|���}ꯡ��Q�5�j�Rg��*�p���;2�}���oM�;���E�U8H�7��ö	b��Aį��E���V'і�y`�����$X���R>R(�nC��9h�/��-
�=4�j�R�A���E"�ߨ/�u�(QR�xQ��;��YPV�{���v&��C��2�����YA�r�Z+��ڬ�^�迂�����|f��Q��-!��K�a~}o��`���rߦ���J���F�q���铪q7E�u������ �"�ҺD84����f�fn_����yL;TKltMΉ(Ƽ@���AlUu���Y�	k~�n��q��D�r���:t�p�[@)F��+2����S2��?8�2����I���s�M����-sר�V�,`���^���ɜq���"B�$��+��#V�]��Ʈ�P�ޫ�@��7p�����ދ�Ms]���s�w�@�׈H�N��h�ǇZJ���E�Yc���~>�P�3,�I��ꠘ�6��'�x�@8���,.��H� K��ɬ�'���4��tz�!�,#Eyڹ��ԛ��-���4c������3��!��$����X��LW�<�;)�������nme|L���>!�؂���u�"9����h��v͋�9�R�359��v��"�]����gO�b삇���u�j�J��N��z�k����߂扌�����Y���y2,*�����yG�����W��#��I��K���1�3�{g��i��=xo;P<DE�{�W�m:�^�EҒ���h��UX�����*W�4:��a�"'����������x�:�K;ƙ~9LT�S.��?�K-D�=w�k���R����5����2@�B�lpXL0���~Yp��h�T��<��ejNH(Փo�2X#�J�2k��dw��yj]Q���7�x��a�ۤ���w�ܛ�,_PP�����,XX��M�h~�����kh�T��@��1%�Q?5��]Wĵ-C�<l���p6OK�`
3��4���(X���9�/I%Z�S�Rz�]��R�qg��w��D�M!q �a��&Yuf���w&Ҩ/l����t3/;^����(qv �Z��[��f_�h� ]�f1k���4>��B�c~n��R���%�/��Y4�F~�!�=����u�|4�#����d̀��x_����"ƝC!i�ר��8�;RCu��i-� �o�"��[�g���gѣ!H�m�!���Ʌ��N0(\�Ͷ���;���=7�G
�*�w��g_���>5����GN⇛,MÍ��py�,D(~�SM���c�Js���eD�dJ� �[!�w�7�G���~�Q�iW��$g��x"�	Jf�E�u�DB+6�wq��]D3ߞ����M���0>�� Cx�o��1Xn qD���`$��`-�=G4xfy�Q�g�,�b�+�n�7M����.尖�M�D�������O���~�\��~��`��?D.?�~ȏ�����=���q�#�j�/Pp�ooh���-��W���duN�����j��=)�	F#2Z\�͍�D���� �ș�~��Y�ܿ����:�َ]"IE�D�U��_�	S��Q^^Q2�MQM/�����%���{ov����	�'��|,����%a�2�����Ҏ���6�-�li|�Ge����B5z�Ր<$�Ɲ�u�$�(q\��s L5	�7�S��9�'�y�E�����yg%|Ӊ=\��y/��޹�1�X�@�z��P1b.�����P�����@�����RÉ��AU`KA+Lz�	˯~Q�<��eՓrS���K+������c�e��5dwn�(3
6���W��eR�`��~T���.$l���?<L@�\c�.���M���r���(��u(�X�sM����,����_��=/��+R�A��EP`~W�8�x�s�����m9����z�,�)�mVq���z��WO���)���\Z�1<��.����W��'_.�k���X�B�L��B �|G�^�Tk�k<�r׆ng$M�"���O�3=�>G	����6�<usqkL�����t�գ���e��_l4�;�+�z���<ð)��Q�D�Gސ5	����l����΁h�A1˒��:x*RO����k��n|��4�b��b&�ν��#~��5��!g u��x��m�A�����
�Gq-ҥ��o��L̏W���m+��䖖����+T#��������n�p�K7o83�]5"Nq���j��Y�77�����I=��i�7���`�fr��V
A�?�O\s=P} �oص"mQR��
��(�)g9	�m-��?�&�9C�&pP�uN��:�<B3��czJ���	��5�)DvR!�@��Fa�{��9��kZSe��1Su���=��5����i��6z��t_Rς!r�� Q�K�z~�j)c�}�}�װW�a1 Q�C���;ݧ¾׀k��D�;N� ���8N�B���C N���v4�e�1�؁�@��y��#r{;�i}�/�5ǯ�|}:xU��� P�A7���j �#�8�Z�.�XI1BS䫓��w���[j	�
�ִ�r�����3��Qj�T&�����0��x�3 ��λ��-�Oi�#R��5c�>x�� UZ/ v��S��� ���,t����&w�ZO�Q��3X<Ƨ+��o�j���u��jI	4u�Q��r|�:S�t� )�kj���!q�%C�-fH`���]{U�5I� (�u���5�:�Yk�pD�UB�kz����2�D�)��j��@���`2������ ���H�P�nF�9���f�E����Y_���x8���C���ڈ�P��'��F��yC�Zm��T��i��,�H3��;�v�M�Lv$��a��b���<����Z��V���,�sի��<�����#�`�u���"�`:�$���Q%� �x���1�N�}��9���|%ֶG8��~Z���$<�d�ǧS�����8��N%�ap��u�`kj��W�����EM�ȹe�NF^�}��I7޷�an��c��z�;�Ku>@�8k���Sf+�g=����<�d�|$ưK�h�1B�W�F�p��F�7����lQ�� �$�����ޡ_��_�P@��PZ��)D�H���A��JS��1�2�S��9����ɀ;��G�<fy�D�{��e؞*�/bN�D{�5�)�yP�= 3�yM�3#�6 �[�A�}QG�IšGS���4o��A�穰�0�e�t�?	�-u�@n
;�HܖmE@��k��P`�$P ���,��]���k��7�;V�9r��C�_�m�(����p��8��u�FZ[��j���!9�*8~P%,���l��dP��mˊ]/-�ӝ����F��W@w�~C�*WC��w��/C�>&��02����#�������ԅ���� F�+G��)���d�w�f$�c^��Z�V�$Dr7=3�[cJ/<�r2�h`r
<T�~6��"zI݀n8��YG����4P�s�}K})������Yww��;�����Ӗ������, �հBEmO �������Ѐ�)����c� �n<*������V�-h�+�"N��颱��J67x$��W2����$NjUX||-�y��N	��Ѷo�w�ex���M����6��m���<䂔��۟��շ^ �JPU�7j�.�=_#E�������4������gYCv$��9vU�n/�D��Ï���B�M�5�'� �痒�������
�������9jkw���Ա���՗��ww��/�X!k\d�O���7�`'��V�o��g���k�o�gϝ9��-o���ѳD�j*Ϟ��h܂��Ɯ����
0��<�"YC�zAH w��G�+��3d�ݩ?̪\�7*>��ͱ0�5�=��J*��2�☑	\��������3�)7i=+�,�dq���v���=�9�V�S�6BI�R�D�bJ� ��2���@lNHis2�|����'&��������	�����	����V3J	����(�% n��EH_�/,M���\vت���������՘�����*��J�U*xuJ+*�q�#��' �V=t�y���߱�X�1�V�)Ϭid�z3����q�}OӞ��Ew2ꍞ��-��m�ci�IY���%�A8�D:��䤉#�Oa釋�����z�3�s�B�_�����M��$�ձ�I[�{ckC����~�R����7�%7��x��U�@�C�v������,�'�"���<�����(��F�~��E"�eG]��拈��|tߧ~�Z�U�%]�׵=pߓ$�]{r�~�������$��ReM�Ӎ���A>x;έ�iA�<�O�VҊ0&,��8�$���+��E7m�����"�n���eu��?8�!�fY
��������C��]x�(�+����o۫��6+I���x���&�����]ۂ.�n����M�a�Q:h��^.���S5��d�L��?f@�5�C�j5�E��G<���Sߏ�}����W[j�f�x� ��v߳	�k�-��T��;��'��X�g��&פ��d
`^��-i�.��V�z�p,�o��Xh�_�������T����M%ّ�F[ �aq�)K5Ԋ�X�����yj����� ����W���
����m',�$`�Y�]
���5��#ZZ#cp1��"�Q"t���u�#u�k�{O����0��5;Un� �"���u�r��gK@$���S�l�}��QW�W��M�	�C6^he�'�N���If�|��i HP���Ǐ`���j Mt�(�o���&����Ic8��8l9�W�jf�a��I/j$Rb�oA��!\sp?s�& �����W�VP�T0�|ȾGµ��B���3�]R�]L���{����w�#7ϵ�E�6�ŊF��]}�W�S�����R�6���l����:$Η��B��i _?�j��w{�-,c��(����i����Û�m�\3S�))]&@u�MNA��x��R��O�it�"�kkm�d�$�w�.@w�,b㠹tk[�]��\�|e��˳��^��7�	�t��hPW�ʊ㒬�7��,��!��f�������p�3S�A%5#�����C��Z�pH�W�j3���F����*D��GNep^��.���|P��k��O�(�'"$����k��U�؅��)M�����}����O8oM{������}��ӟ�o�������?Q�3H�&��Ͷ��h��Uk�;
�p�2ʘ@����#�v>�^A�Y��l+wsC��І�I��^jY�I>�x��6���j���ZZ]�	>���E6F7�K��S�\�JyY�1�~��g=E�q9@��I;��O,mx �V�H�Y�\t��\��z����5���t�$�!�`o��O�������Xi�����a	m�3�(�չ�Ё9V�3_Ee�%+H�.�Y�4�$���Y�E�9����y�7���F���]�u�2;;��f�{�J�����|?q/JB�ؼ�;!�K{X6��o��<�GJ�ʜ��.���9����y�G���G�h�cjL���ۈYm!Ղ�GQH�����qK��� $�w�1�n���y,ށ=8�|f�	�Q	�i*U��0�P��T
�C����RU��M=�)�Ö�Ƹ����c��uh܀������Qo�����b�s�S	�P��SI�,� E�KR�a�u$�]\g/v��Wf��y�uWXy�mc�wW�����b�s�5&��&ޟQU��ӘUhYs����6�e%�0��Rz/� �@�Dc���-�
� v�{s��1���'u��F�C�Kj�Þp�O���́�C�%s�׉��q=���-�řA�?cUWC��S�#F�ւ���JPH
�@�j1��h��tќ�#)�N�(�ƮASܔ�J��v���>�[�����n|�1JE�6���ڜ5

�����G��ώ@0ȇ~"��r�{ʓ~^�r���2&ܡ��K��.�,ҽ@�\5�R?��)q��i���;y�S�����d��69
e���(������"��wN"��.g}��@Sٲ�#R]�쟕]l�Kd�繅حI���I�p���(�vg��9�M,w��\k!ay����vr�����U^����-eŎ��[WOd⸵?�=w��.���D��\E�`��ռBRr��tv�.��TTji*�3�N���B�}����� 7e7$FZ?@w����-S��9p�)T���K��xQ�K��+Y�]m���y抄�?	�N�c�Ƞ�WGrC��}+� [D���%�1Z����=}o!�50v(��)c�迅��S�/���i��f����^=#�D7��}>����B�IZT�2���/-M[��!�	t�X̃\ Ň#'2��u��@�ϰ��ܘ|�W�+
DQd��UԔk��e*�����9�����osR@~s�	0|�B)��#.�3���<ݱ�Ҭds�)�����s)E�1�f�u�% ���ݏ���*�V�3�8�L���v���d9�Fػ�)���5�څx@X�Ц���v�ZPpnܤ�	-m��$� k�D�"������)��+m�S�Tt�ݮ|	'��"�S�O���h���Ae!��))�i�S c+wXy�[$�jl�Q����.�\4���AL4�O��e�y���
0!=�yGG4wQCx�a)�i���֘,�L�ZF_mwc�~?"p�fC�F�K燴I��ì4q�k�vW�Ȭ�A�u�M��9{�t�UJ /àr��V�9��`|�eb��h@�ݾI�y3x�9-t?(�A�c#
����nUs]t��Շv���IۚB�	����q�w�'!Y+�$�J;�TL��|�T��cKD��Z�����ba�v�18<P�*�1~���x�Oʒ���W,�L8+!�t�y����+�@�(<�K���k�N0�a$�/DI�b6�����G+�)4��	5.������7\�l��8���II<�.�!�j�1�,z�@W�CgC w��qZ�I֘�� c�6$eK����*]���qs��t�Sq҆��/�������K�N1M�����"u�KXg�^�I��l0/���k�Ⱦ��&1��/�0��E�f)S{
R�p��cN�2L�x�{ZTx���?�0�_�m6�o ��:���@=�f����܊Y�z�/�$�k*�)���
5�]넧Y.��J�)h��6���<��m�!���(-�CZ��n\�{�׏����.Y����Fq剕�kg^H���"yy�[�Ǒ��eiqN�;|#���>/�/ma��8	����T���m�A�4���!*�bz�
�LN�w���/��z�J��\�pB��oD���t�~	F=-!���ڼ�k>���#�?-M�Zr�	�����$����,"�l�qՑ'_��zO��YZe��3����vT���������GD��f�K5����������.Z�\N�G��{Q��v�چ�6����%����'*�"�"`SB�k9�1,p�De���jk��٣Iu%A�XcR ��S��7dEa|��2�H,$�ĲͻFu�����HfVb+��s]
*ܤG2ݢ;C<XĢ���Ə�<��t�V��ZW�Պ5�C~��L ��I$����U�P����wvn��7�������>B��Y35\0�m���4�������~eQV�hV�-�s`�a;#�|�� 0�,��ѩ����_YI�8��@�o8�ڇ��.X�l@k�eHhwB���t�;���^n\���*��T����=��u�q��@l�z��/XXn6y��v���~M�-Œ��!�p�X��Ae�X�y
��̗����Ȅ�5T��:GZ�ʣ��Ȅ�N �A���&�zE�Tr	�����]0��ڸ�Oq_��}�m��Qb�2��=� �>�ZlDL����w�IgZ�'�ؒA�9V��Na�,o]����IF	����:��#��o�>����L�a8���}s�Z�-,�~�/a�./j��S�hۿ�(���l2��W�9q��by!q�XT� O$�X��)q���ܩ��,*���/�Ɔ��b�!�CP�䳮�ծ�P�+�v�j�+�B�]د^���'޽��O��
o�M�/�n�1�!�����Z�H�u-$�����=̜�j�Lh\7jE�h~���s�/��K���T=U�=�d7��=;�$C�R�n�J�ΐ&���T��.8G����fP�t@�3��Qt����$v��D�F�Ӿ�HR ��"mk	�N�U�5��̓֨ha.F��J��d�c�DT(�숪�"G��D:v3� ��@�2��IgVB��/��^����+`�?/���Q<�9l��iXg�7�_*m��2�"��ׄ�?L�.���	oQ6��7!a����͂��ME�Y��4�X<�>e�K�4n��y�S��jlTI�����8��Gm� ޭG�/�g�k�Z0o�N�ĂQ�G�x��r`|<s�di�#|fR�{�Ġ���W�kW���d�7�'��ϴ4�s�	Bo?#x�W����ͩ��0����1���L>'���b�C���PP�6���f�1_,�DqҾ����OF2�P?^.e��ul�r��\M�� u�����9�]��`�u*�� lW��X�� 6�ŵ��m�-7�F��S��k-
p��0w�\o�� �~:�s��2�4��1���c�t�9qߟV~�cdiH��h�Xu��7����w{�<C�m��~HC�_g���\�Kّ�'�L�n��o7��[jK���n٪[��6��`z�qH�C����)[s��0R=���xGq���j��"�ˋ�䬒t��RS�r��l�jD��.$����	� ��_�*t���P&@�ř��i��Jc�#��摋jH��1�:WF�R~��Q���'��kP��;?Q��-OdJm,?��O�
�x�g��zD��ߣ��MV(�ݙ��lp*x��+'��t����]�dg����,�M'զp<��UM�k&9��ܬ���C��D?=UFj����fsi�P���^�&�N՛y�����x0d�T���;&eʦ
��凙뺤��'��`.����tӭ�LYp �f�c'3�s�A�H���pT����A,G�x�����!��i8���������z��7���Ȫ��^a�ִ��{3��X[Ba�"�\�F���os��g�����#��~t�OZ������d�n��5�(��섚�Y��ҕO���;�$%\o!`2���ٍ�6���u�~z^�X����h��S��J˹L B�O��x���Q=NI��q����]e�1]�n~���D0r]����ګ�j���zg��Ͼ�o����qi��tK��&��!��"�ɍ�씋m���Fɉ0[ԔF*�?[G����[(�x��Sվ���a���>
ឩG�//)
KQ�_��!{(`ܯ�/h��vG���w ����������*nM)吉A��5��V��w���������veA��:[oN��M-��z9aIJsNx�c?��/�_k�\�X5"2܀���7�1C���~W�58��|ʊ��){6xI�\��S�(�3v�qQj���7~�L�<�PD�׳������ս���C 9=WZw�`u|M��� �����#�%��n�Ǘ��`+P�h�v}#�P�V|�d�:�L�I��C7��y��ʗ8��MK����:�?J���t��B&��e
:#tY��]+����z��"���$��JK���pN�(ɫ3ڎyq�9t:*iI�Lj�~px����M��v.��^s�y�aH6_�oog�P�L�w����M��Ja`�?Un�YKo��Vn�$�<�8$����2��2m�MA�Y��`
��k�P�B@a��5�q-�)��-s*��:��͜���
�G�`W�#DZR�Ó��	Ø��e�ܳ�����:Ϟ,��Z��<<7�����I�Y<{�a�_�,y@}n�K86c>D��[�>r1#�V��ga�e���'���Ho��.(_����p��vr۲1��%~�`G-��:��eK�(r_=�7�ͺs�p>KQX�|�]i�h�f�����K��v�-����~e�`��`�ފ�P<'EFx�2��`TS-}��%�^ʹv�.�\u�H��F3��x��m��ه�N��3���r�����RCEo�Iq6��w�C['� =\��G�~��`�s�G�<�j^
��
����!�z��eɥf�'��M�ˉ u�S�I�bm�E���І�p�B����fГ����%�Q)Ǌ�ە��.���L\��T�BX��JZ�l�/6ZlH����=�t-�6�ׂeq��N� 8��g�Z����!��ɾ��g��A"��m5xlk�
�O`��W����)��
*��"|ǝ�� D��3UѰ�ft�87M>X���.�i�IǠ�R�d��VBNB��j��*�L,2)�t@��L5`��Wx\̒�#�FǕ]� l�&IO;Q�r�!�{8fЙ�!������8�K㓿��5Ī�j`e%���W�X�!֞�T�5�*�&
`�n�������S�-��x'�d7�n-㧣Q/'��k��PbEzO��-f�.�����t�[����t��K�?-Бh����0L߈P�xD5��6ƍ�OB�)y}��NOQ�z����i����=G�y-�,��fZ�=�cj_�Q̖ x`Z��-kN@�����%�u+���6�O}�#(�<�S���4��|��T�����>��a�"�X���Y
TDE<'�~Ȃ<�ء����A��6s<zn���9%H�v� �(�����B�`��C� 	�b��2�Փ�+Ghj(G���?�PT:�����0�P�_/*O~�����Q�')����J��ŦM���_c<��n��f;��nJ��~b�� \֌���x_��A�Y����$���K	K8ʿ��Ӎ7^"ĉQ��Q�E+��:z����e�#�'Sp^�M�=u�vRȁU@?$�x�/�m�Qɓ���|9�~�~���H6a�/���B&��5r�Hة��\C�~�g�)�L	�(���ˬ���-y�w	��!BÃ-��n�9�
 ���k�$�w"l�X��4���.yqc� ��=4G
��x�L��S����A7���S+oaI�3Ew�����37��6�F7�!+t���F��5����j�ɲ0�b�&�����2����Ѷ����C�:��勣�ɐ�!��W"���'l����qd��D$N���w�0�T��:�}D��1-�%��Ģ�lI�-4���fҖΗ� �os)���� �p̬E�2�<d!�k��s��	���S&���#��!����v����k�� �f��W��9=����l�����c@��Hf6��Kz>干n�O������49&���I1���M>"�"��3��x�+ҜD���V���ǐ�^���j U9�e?$�kg��%2�����������zG�]y��cf�q�劯H�)��b�{X�v����k+�Q�֗�_w��\������H�!]J���ܪ8�u��<��`���fP�7~�;_�,������@���A�rlZ��:�q�.|�6��Zs��[�1��k:��2�wq^���"E� s�IE���z�]����ԑ�5#��~@h�ӽ>��=���d 4	���BZ�4~�_.0$�����J�R�Qŷ���z��m�`�W=R`+x��J��v�j�d<���XAѿ���ij�XJ�� z�9�猋y�_��b�~���vNJ�F�8�]�C9�3HU��h��� ��_'o,u�9�l�طq��d��\��}&J{p���_�X�U��5���̆:K�������Y�m�7+{&�V)D"%T��eT`��<`6gC<�s���W����x���=���I���Yd&7LB�힤���05K2A��1|W��돪3�S.��M�͜����V��*`V��?H���ݎ�c?'\VvN`�h�n³&��wj�g��h4�d��kŰa��ύ�r�ndS�3#B=8Im�K|�h0�i�Ⴣ�1�~?�6����j<�����ŚM�B>=�����P*U�d����ؙX`�Ӛx���56�r�J4����yflԽ�/�ԕ���p4�D3�lN/[>
Jg>�ki� ��<Li�( ��ѕ%<M �J��#cB�vh�Q8�ѵ]����[�p�����^"1{���u������|a���.�RH��y>}e��������ēw23�h'�鄠�!�����0�#"BN���X�c��@V�Y�=B.��z
f��d�J�������:�7�7�CvͶ���J-ʌ�e֞�}k�)�lICt���gUmi���}ݥx����1��/J�7�)�߱��׀ "�i9��a��J���N��3RcL�Cۜ5��G�O��  �J�>V��ǅ�1o�^-��8wR	�D�k�]y|e�n�T��4�!�.��&g��2�CSEP��{`>i������x0�S��(���ʱ����[�3��������
�WK�^�j�D�(�'b*U��Gq`���R��#$�2�	8�����/�8����2r����Vek;ө8�z�M�^��.�����vz��l�/�������ݶ��c�ƪP��I��a�&�Dk)��$��F?68���%��)��׿������>��O�U��F�����;8��9Fs|���g�$v��'�"��=]�zDȺ_={\%�Jh�U�!�W0�+�F�7��f�t��ہ,���g-;D|�k�{n��л����5��G� ����U�f���1)T5���_�Wk�´���GYȹϾ΢���������������X����_$צ-Åw?
G��W�!�t9�Ž��Z){�q��앑]�^+�p���n����,��������EZY�3)ZV��c���yG̞��hX�]�b���*�Bsk�{J�B���F�'�	1FD,��0�!'��a�nY��dn�/�B��:�K3cU�k#C(C ˎ.��6E[�L'��*�?8�'�dfc�ԓ\KI���� ՞��}@ɔ�Ղ3�䂨��Q"�8���xP"բKû�	{�B�}�h�i��3*� ���$�l��ؽv8�xVM����ۢd�Lg�NO4MA[�4���J'8������H�dvqfP�-��m�C�;=�����zq5�;������j�3.��K�7_�����O>eM0�,Vm��|i��r�2��Ci�K�ڑ����{,_�O�{%i�7��>�D#1:�����MU+��RR���6G��nvPq�{��·-��W1�y|�@ȉ���<�Ŭl���h�dƺ �&�ٿ�8���I�t�lIc�^��$�ih1���:��O��|�?���[��ک�q��G�� ��V]b�j0RP���:�KkSێ.�E��D
�����ȷ	����g�V��وRp�+��u*�hU���x�՘�I��W&�۴��`7	bC��f�42��H�U./FY��_��mz02�s�ɿ���c��D���f��7�?]�(G]mx,m5�y���'��=��t[���/!�K��@Ej�m4��{�-��ޡ��Tm��U3���w,�OCc�xΣpdG�}
b���t�3�g��}���6�s���~��=״x���.A�JZ�⦀88H��;��;�s������_2`V;���e�_�F~ \ǑqT̆��w�����
G��E9!Z�.p���O|�9kI�a[ۀ':�q�A��z���$JXd�SH�1�6qC�It&mZ)S�����R/���)f�>|ч1���ޥ��'+��dB�xW�oo)�B&`T�11���)�������k���ۧh���1q�/��Ӹ��������7�5�+�X��+Kn��&���U�;����S��FvJ/v	��:����eوX���:�m��[�imםY���E� ���h�P%S1v���ZFK«�t����QH�,���<~�nX��Tǿ�ցC�׋�P�s`�������sJD��ȘIç!�V=��{P@N��D�ŵ��\����������7N[5�
���OU���U'hM���w�2��ռ���a���4	�io�3)���]B|��s�[Iq �y��aΓό��G%�.C����!6��%��K�>����`�A��^KҢ��
�	s#|��6��̘Gt��]C�+h�h��+���"�I���Ε�]
��]��!������Lx��%&r�A�}��+��㎊�tӴ{b!=,V�x-���e	#؉�X�أ�_r��Q0�1�q�s��bD{��麢z�s"R
!���uz|���Br�nK�?���M�>��-�0��H����a3K�{�a{ॳ}D��Z��NWֈ�DTyi�n�R
�6��AP���d.�-�Ъ�h�\*-Qg*|#P�w�f�(���ſOy4ƸÃ��C���p�ڙh�"���H��>�=Ip�*3w�%��*��H!*�݆���yeWx�PR`"�],U�ϥ����ף�UEXlF˝�5�Èٽ��c1�!C"bQp�R4�(������E_��\�f��/'<��0>�-�B�|V�[�4��W�
\ �->���X\�)k'��
]���.\��/���}a�20�+sg����8�rI�M��b���{N�x�ϟ�z�L%��w����7��ZG�x@иVxG{E?��fu�<��楴�m��D	���@*D^��;�
�sL���1��H��5�����K�8,�<_˼��N��`n�Z��,\6��P���ؖ�?����h�� ��<���o�C��K:��¸��ðXp�c�E���sW���K��|�y�,��ą��Z�7NF�TA����qXP�{ Y�}�$�^�ԸB|&U�D�&&�HAx��X�\R���e?&q�/�oe���l��<�l��s�������k��YF��p3WU]XS�މ�>@�o/:�/O������	k���-�4\s*�4�<�5c!���%'�[�!-�������+D�a�,���m�M�f����eo�����&Ǳ��měp��e��fY��!~�Z�O�ql�.�G�4hG��3'h��$�OuP4]��9�����j����ǥ����zY�f����wU�|y�����bz���^��	�-��qJ��g������em�1�YQhcUp%��J�O�
��������4��m��ZUh䈡���~�s��/g�i9B��>��J���H�7@��%"�����B@F�e|Y��������sy����_��\�d����q�M�6m�+��B9�-�f��3�Av}����dN"���|qW{β@�����=��9 :���<K��[��oP���!]V��H���Ԯ�2"m�}�zgT]=�w�J�vφu:Gř�$<iU��q����X��=I(�y�q�>3w��A[���A��zWa5���|����Qz�G��j� ��p!m���LwFo�����aӧ�VӅ�HI}Ð�^��W��ި� ����(��y|�L$��>߯�^�5�T�(�򧸁���-�q8����W�4����˭�t`��v�?p�5gv�h���b�sݾ�j78�K9W��Pݛ.
�9K����~T�б�/�p��TB �ܽ��� h�&�:���v��>��xo˕~����7�Y�c�m)(�TIT������?�*����}�����p�^��
�=�:E��Aw��D���}Y�#b11P]�ܦ���`ϛ��J�l��m}׊�#����8|��N+EE��s0������?��*�bP/-���h�BC'W�:��&�^(=m�sfO���d�8c8�V��Z�ڊ��v�_�jc�(�L �FZȃG����[�L7����Dx�������V<\,#�HU�,�q�ߢ	�sꨊ�#1f�xB�`�Nd���frm��5u&�Ȁgdz(F??)����-ln ��M�8��ؿ0�׳rD���&��g���m��'
���]I3Z��sD�Cn��b40Ev���&��\d90����D4�y*��I"^������i���.�˕�����l� ip�[�R����ܑY���$�A�J���	��p�O�/����L�y�3o~���<��9-)�0 �q����s�;��MoO�乓�ٛb�L%\�����,?3[X���ʎ߷��*��`�1���?f�_��/;�䘅]���e�w��g܆
Hp_�~��Z��%���!��~��"X۴4�hp�Z��񽟭TQ�f>��yJz2��i�Ǡ��K����G�_��S���4]�������J[�-��6�Y4&�G)����̤lj~H����U ��<�O�����_$�(��F�/�b�ރֱA���1�%Ae/�~B�"Ѯ���;��IUH�v�P���z�fE9z�#�~}�T\FʵA�^Cj�d7?o�h�0��h��0��KV�6��ä�:�/�
���g���|��i
Z��P:EF��-v��Z��|�����<%�n�T���s,ӹ�@LG��~��߻���������΢.�\�V0u�Zu��}%jU��|ɗxx7�G�[aoL̈���z�P���]���*�v�����l���@F��==>�p�x�Ų��u�u ���N-� X'��/%:�N� �Xkq�o����|�w����u��	�& �z��Ћ��w��|:틭_R4W��#������*��ϩJ!���5���V�{�h<8��vK5Ճ�u�S�Fji��#�������-����� �t�v�U�7���s�3�����	�_����RDZ&�~��ƛ�Y�)�OOøk�Am�LZ��0b��@� )H{�N�N����
l��;E��Q]��~Sl��$J�M�:K=��юpX�ؒ��H�Y�+�塃���نDd~$!�"\.�7�`��*�'�E>�?*쨓OP��oO�\0���3���ػ�FzQGf��K���h�Q�2t�Yv��T�f�vi�6����FسT�w��Mr�(t�����ג��� #V��(�ƅ$6()0�����X�H�S����0��W��S��d��PA0���7L_�:�j��8i���GL�H���̢;;�>�O�����y����w]�_���֢M&�W�>���ǳ��EM�����t�4�S�[�0^�_�թ�'G:����{!�<YeJ�,�_�����:��_C��\�
.{_�SH!(:B�.E&�`6���y��3ӳzM�>����èL_��N7�2_R\���s�Ƙ+C�h:�Ħ	� �2o��2����S��NJ����-p%@�\����;�3�e͸(�v��EGť��"J�2۬�k����9��t!� �^�[tg5@��~�����z�N�u>kuIq��Y�"M��2X�m���K�f0���/S�^�J?�{����<}�����"U�$
$���2cޖ7}�l&A>�).dn;��%kw����	ޙ�y�~�p���v��i��12��L���~���g�FP?g���T���~�{�$c#��LיĽ��2���
DS���s�s
O�7?׽�:
e�]	|݄N�#��h!`;MQ��_N%�CКhE�,YP��Fr#h���yϒ�����**油ڠR؜�bK��Q�'}���O����7�L��D��]��S�zv�M7;���~��۝oSړ�)e�R���V�|�����ta�؝y]�h������ٟ�)��UQ�wK�׿��8�A"�G��vmv�i̲�+[��~#�/.(k�B*F��C|��:�6:�|AKO�c���SkۚA���o0#��9TN�j��pkM?�R8�Z��-��;��$B^I�p���@$�ʞ�cpo�ٓ���G��<E�Q�Ȫ@6�*�n���	��i�9�i��y'�^�̓�'"�Lv>��1mX:M_�o�Iŧ�K_٨�q�<�����3i.����瓳B_0���tt\!���)��>�|�8��*�X�L�B8�_ե�<���{��(��Lp�9��
W��N���C����s�\�Fk��Z�ߡ�V�\R Z��&:T���F_�*�z�����9���XQ��Ɛ�����
��}_M�J<~^RGW��N��&�M͔�С8��Ġ�-?>��>4��Z��� �!D}C������R�یpko�O� ���`�Hb�8%�}�VjI��O�N�����<Ϧ��&=�	}�!�N0�SCa�Qt�nH=���IP�-t�q�w&����?߆�Ү�8[�P'��x��C�, 2#�2��0�wA�M��!<Q��b4�(u�������-x[l��Ga|�'���EaT�V'Q����I�.�N^aGQ�v-&����fH�<2��F>�1VEځ��19V~�"�
�ON1�@���"|�VV�`���B�df��Ǒ�$w���ہ�j��v���q&�զ�yakތ��\z2V�q:��"�!|��j��ڈkE�8/M��rtG�,�'���_b8�yE�|������?t����X��E�ƵB���?w�-����?���Mt����m�������pT�)��K���d�x���X�C)�4�r�*���ہiB��d!����ϷA���>�f>��s����,2�`���D����=UH\�!���j'=4�.��sN�2?d�BK򇢗�]tUX���M���eZ�׮�~��AJmr�����"�6ZZ��SsC�@�p�6��+I8�k��C�w��� �e`�Œ�0`��:��%��b�X��P�q����+z���V��#��GN��>W�d�-�͘�D@�D��O�Ҧ$�k`5��$1���^��-3t5!���9�(��11g��ê_
[�������!���=�/�͑+� �>� C|92w*��}�:^h4�W�ok=�lL�W �y�=m8��ؗ1�OIG լ���h�Z�4�)�X�xx�r��c;ٱ����q����8�_h=��OS��b,(�A	$�Ek�&ݷt�M�sΘb6����b��S�Q\n؏ ��\x�ff��������^�{x_`���R��qy�T��<:'Uo��>%��Bs��]Q�e�=�4�:~����	���'f���R�/e���2d_f<�|RC7�uS��;?7�V���w��W�9<��IGf?�pˈ#�T���{4=U����=m�!� _E�0%�,��-DM�z���lb��׾_�ѡ�a��G{���-�",�r^�X"�-$�W��!���*�pz�HfP�׃��w���c�oW���m�/���r ��`�L(W�-B���M璅ќ�Dp��a���1������)�"���|��(�~K$.��B]�,ج%n�Y>4��4�=�<��l��� ��9�� i7����"���[���;��"�a?�W"�1��"�A��2Ueu�U��r?���1Ƣ�KZ�
�:'"�p@��F�@�R�B~��k���_~s[�3��F�~�r�a�!�[���	w��yi��Ry\ŇI��GP��Ǫ��97諳�����e�ϲ���c²W$�ke:�T�t�r�����	f�wh)����^�`1P&�d�&��9�m��͸s�N��}C��+Y,a	�B�@h�2d�"��/˝4�7��(�D�&Ҙ(�{k(����
�Q1~!Ǖg���j��)1=�,tO���8�(ڡ���'��\�vE7�`@^��ut"�ShJ��{0�ڧQ�lN�F���+��� �Ǡ�� }��H�����#���Z�u9�&�P�E��8��K(��a�1��7�a8~{fGF���/
�f�~3؀�L�wy{/E�:�)��5�ו��)�I�GCA%{:���dc��c�x�Q ��x����ǽ�XҤ]�B}�"]��M2������F��A�^~reNn�3��W�'�R	��͜��H�!0y�ڠy��0Ɓ��E�wvIA��F}�׼�PZ��;�.^As[F��Nx`��['��4�x�u~r�o�n�����&L��b�2"���k�N��O�`a`���{+�c/C#P?�D�J�{rη���u)���[U�B{�|4D�k{'_�}�*�Y vTuf 0�["�+�����3vΨBQ�iE��p|��d�]�o�dy2��0.��|V>���}�	{H��#�8qz6*c~��H�EB6�HVyO����[�(�� ~���y�F-�5��:̈/<�9_�E�rq��`#bC��D\:
��t"g�����{G��Ba��-�W�sU���1f	���h�� ���}tA��i(uE��Ī.Up����Vn���M�J����n���g(���WF
����Ul�gX5Y	ʷ�)Bd�Aq��_ĝprѪ�����kJ"(��Y$m �)�A���m���/I�q�(>1�����qȍ�Q�4(⩱y��?�>��"�E�8��ߝ{=�H1̊!]?��Z��$)L�Xv�� x÷�g�ܰ;�+�3'��S��,���M`��ô��5']���(�E�������b���B%����;�'��V5��3Z���j�ih'樟Y�d��!a�`tL�pϨ�F��W'UWQ$�t��c�i,i�M5��b=d �F����
#(��>7Z4�ě�����1|uR��.d�B��/W�G5���4"�e+��0�t�\��T�gD	�W�(!����X��o��._�iM��.��>���5��H9����"e�"쁇,���i�PWUwm$��>2h�&��s��տ�h��z1�'�
��U���u����ye9�<����ߊ�I��4b\��To��A�,�U��:�d�Ϧ&v+0�8/�]��������I�N��׈R��ј�Ƅg2��c_�n�+i��R��-Uor<����ގt�����#L��&�6F���A�zc��	��2л��p���?��� �1i>�J&�	fF+�T�S�zX(�V�X�� �f̌���׾��:�a}QS��c[ZE�A�G���Ս�V���ez����
Z�����zm�*}����i��kƊd2�k��e�U�X�('0�vj��Τ��P���η^�iȂ��Ɉ��1kȃ���fYk��I�@�Ik�{)o/?"�����r��2�C�Ef�����yކl����8�ow\g��*ȵ�����N$9ez�C�Հ_�!+�|}[�Z�wx�/q�uw��d(FQ)	ڭgn����a�iKD�rU�H�-��ΣA��d���^h^���oA�m���ؑ����%����!�=.�<�8��Qo]Wd!�rQrQP�&���^��!s���W:P��*n�gPmUqW�Py���8�XUȍ0�~�q'S�Qj��e���9#~�O�`���[�*���h䍾�j�v�<��iJ��]qk#
�]*�v��w�Bn:�9���HgOl���"����P�\.1ԕ>������Õ�ӳ��8���]�Lib�������$Ʌ�#��he]S��m�⥻{t����$�}�������X9��:�L��-�OI �������"�-u�ol�E���{��^�����X��|�Q�b5���v���_�i{W�{$O��>Jv�wA,�O���A�`;��rJ�=eט?��k�}z��� �����Wln-�Mv����W(�5y�vp��G����.i���%܏#BfaO��qy�9�Qb��i�8�p)ܛ�<�Q��2%�T����d?]��,����V��"o����Z�ю�*1���,4�"����+�����+/H^�|�s���b|駊l�0���J���?��<���7�1��3k�쐥�e${��F;�\������
��Y���ArݙT��1{�͗�]b�Q���=D|�[H����EH)ǭ�b����������z;�c� e=X�=�w't V��yf���*�|�d�a��G�c.�I�k| �%����=t�s�w���`и.2�ѷ�؆��r|���� �pJe7�����9Ŝ ��[»�0�=	(�f*ܬM'��M��o�Kѥ�q��[������>�`uy����ha��i���ԉ͎*Ԇɠ:D	����z�0�� 򎞆e��?]��ى�9V��"��M2g4�%ℇ�~!�H�!ۈ�`�ϳ��u�����wYj6EX�1�Rsp�c�����̨D���z���K��zp57
�9�8�Wb����ŀ
�8w\g�+���S��N*�͠#2�tC��ꉠ�����L�ǟ�s�-@����?�5���P`�%�mȳ2���>U���J����Ӏ�J�c�)��0�'>ƫꇥO��Z#�&�,vfqi�;�Vי1���ջN���ےAzF��V[ �$>�U]q�����{I~� ȋ��h�`0x�xh����s�E]_��Ob`[p=�g#�h=�;�	�y�&U�n��e�gh��8{�/-f����7Zf�i�
X�M�آ���~�#j�t�|�{��5��E�}��"PF�F����d���3�v_�����]�j�L��W-]��6r���ݒb�
��Pk�:�I��*�@F~ �3��
'(�}�$�1�3�����&���Ēڝz�\�����kF?��&��ްf�EU*Q�δ�Zc�H��(��U��Oz���7��`h��)i����#�q%7s�à��tr�O��R�O�0���>�/��a�:�ؾǣ������KYS��#��'�Ņ�F_�P",�����4Η�e�/� ���W���ΡK�i�nn4gܲB� �7PͿz�{*���ç�Ϙ��u�9��[�<��'�|���]�FV#�o�x+���^*���`�K��C��9������o�"�ه&����K����}����;'�#�ʭII���u��cV���}129��fL�83վ�6�E��mH���D]�ܓ����b{"PKm ��#���%�h��R�UN��=A�(�	[*�HBn�A M���E���)���@��hR���')VWG��;�bl)0�ha��v�td%�mV8||��!�2� I�k������Z,���H��{/��z�ϬN�e�]�;��2��D-�A1Z�$z���P�UYC��E��t���6ȡ��?9w�q��>�+��D0�pG�o��RCg�@��Ce��և�����b�'�Y��f�Tx�-�V�j�=PS����=K���h_�?5�t�5˖���Ѣ�k�����C7̏)"����?yE�ZA��p��l�Y�a�ς{x�[�,����n�Z�!��P8�u��"���)�Eõ��|o������e�v��(�9�����K�3^��!��T����Ĵڻ��[��iygn�����ip���E�ķ�4�0��X/��⮧�]鏚��R�����O�:�w�W��A!�܃w�	����P���T�\�1\h!���J�Qv;$g %L��1��W�8W?z!�NO�oުVjt�y�����&"�\�i�F���l(��UJ��qY�.��3�����Z{�/��`�d5����ī�o��g�����hV/���Q^���U�"��{k��v�D0�g���$�q�-Ֆ1�d=�	�����lĢ��������D(�P��ݼ2��-09-�CZ"-��)��Y(�%X�n� `�n�?�槉�4\IWlO���7�h��f�ִ�n���|��R���6G�{�`HTǢJr�تY�x*���y\)Ȥ�������vթ\%z�uhA��#����zEݣ��ץr�R,�c&�XI�zY���@�%%�z.��pC����pUN�$�'FHRę\�i�\�\���k(�*��Q� U7Y����O��?%Ѩ����/��5Qt���r�^GZ-^���YP'����ena����I8{v�D��Đ�\.�� �L; �N��Fi��o<��z�����B��9����nA���ë^���Ik-�aW͵孉�t_OkML�1�oE�O�M��H�򒈲>�I�;���4����(�k"��y�S��`�Ý�k���V��h u�9�������!oa�`�D��.�n��^��" ����K�tߡ�u���h.-�t�����ٰ�Al|C���L�U�(q@¼��`#�Y����i�9���1�8QTD�G
Ō�?�?�ח^�.�ئ\;a���~% #�P�o���.3�+] �ݷrb�_Cj��98B�����ΚEYA�4����!uڡ����DƮ�7/SB��OE�ժ�e�q�&�t����g�}�Z]�=Ul�3E�l�����r�etV�������Yи{#���
|�
Vֲ�/��pG��΄��t���j��:���ҍ�M�1����yqV׏|gX_pE$G�A>������ߤd�<��m�������$
�OiX��4+�N��	��M�S�7�YX>6�Z����]=�x�6y ���H"!p�e�K�i�`��4�Nr��p����5�A����<*�O�y��H�}O�B����u�AX@V�m�D��g�����v�a� sK@�cMb�-UG+%_h6���~��Кُp��lC��QARH�br�SG#Ic�Vq\U�|9z�O3�̮�pD�&lh
�W�kj�K�5�%Z���,L�,�65u�+����u��$E]n�H��U` �de�ՙ~
�,�3�a	턌���W����Z�����w�#���B�ܗ?��i��w{���,���ZuT����	�]�>X�������̭!���䫈����R�_�F)��%�N����)B����F��<�H��Цd��M�06�o�b��S��vp�!�\Ny��h�m(t�)yb<�J�i��g`"�N7�<���e��PJ�\���-��/,	|~�H�%���f�e�V���Q�wh0A1F�K�_1���#>��ëy����'�l�0V�u,�ox���f5����:Ҁ� �m��&zX5�]��P��j����gK� �芏t2�QPf�����K�/���,b��֖�hr��&�V��a��F
$��ږ��L����ɜ��5�rn9X� /�I�J�RsD���+��8���UU�jZď���C|c* F�{��)��io��v��zh���P�T�<Ekb�^������Vb�O��n*C#ȂO[���[ꈵ	=q�s�%̧���M�F��
/g	���{��e,��7�&�{n�p7QW&>]	jup�O���F�o�y�U���֐H�H(�f��,6�$�	���w�e��3�=�^=�d���'U��ơ����Sjb�1j�Ui}�2~�b���;�A�Z6kc��<��#��p��i�0�![��#&2��$����ԂE�x���~�э�TA|�[Э���&����t� �Z�Y��Y�B	5�vH~M]LZڢ�N���j��'\���	�ͅ�l�u7¶�q*R��R�mA��o=5�v���/|/�zrX]e��5�@�'��ݩ��.�ԏ��2Oj���2�B!�����
��?��-�*�#���e:��q���W���"�w�*ص����ʿ��I ׶ˆ�j�9�5�h��<ފ.�b�����V����S��dP�:�_\a	�L��HB-D�8�$<^½~Yڝ����9 W�Ԟjr��e�^�]���߅T��4�ʏ�V"��0��޴��#_H������ݧ��EAblʤ�R'���E�i�ւáqsi)�7z`*:��X#"�V���.�7s��;����S7�v� E� �1�Qӡe�����7�*���@���(�@db�n��J�.޹��=(��C���0�WN��t!�k��H�jY��Ϟ#��ĺ�t'�e� ���[��ڏ��^�t�MY/s�4��MT3�E�I���.|/�X%��� t����,,��S�O&�O.�p-ͻ{��✪î�Y��o3����f��aس߱��ۇ���pEu�~Gͦ$�Z�����k��NP�^�^�k�G/%zg���}���X�"T������M��!y�tD`
{1+��҈�ά�D*L���hv��J�֪O1�2���d�BS-��Nt�^]w_a��򳵔j�`'�^��٠��Tݶ$G�΋���'�&��:�-�
#r@�t�в�~u��P��E���# �E�:�_U��tL3�&;�%?e�?:ދb�Y�` B۶P�"I����?S�w����N.{�6��mM�gV\�w�P������誹��;1~.��E�����L���rB�䱨�0�",
X�8���W��t��L�ƿGœ����zSL��L�d���5�?AHP�����;��x�K��o�U�u�&^�����?����oZ/�MK&
�~�H�2�%�,o\�����!fLA��ѷ��V�����Qhp��ķ}7�������PN��`J 
Ծ�E4Nc�c"�=^�3��?+��Pe[��T�m�S\�yi����ͻ��w��̖�\x{��陆΅ߪ�`��1�����;6!j�_7hΝ�;�c~D��LL�c����3&�_|���{��S_��Dj�Cq�
�!E���� ;:+*�GA-fQ%�M]Y4F��z����2����Pg{eb��XKaY�T��xo�Aex��f��}��>�1��� ��#�$:�n]��T�s�/�w���oa�(��&��&2�����M�*��	t�"��oO���X߲K�G�����Z�!R���i� k��:��sl^����SO�=?`�z�����a��|S�|��K�U&�{����|�����Bꦛq�\͓����~Q�P��Q#���k	؎���J�h�Dͺ&<�����`-����ݵ	Љ2�cAb6�A�s׳�����t�
��e�%p-���D�1��R�ۭb9�"jNH�����Zi�}� W\_r]b��Q$���a�ڕ$]��+�a���?��&ٍ�Δ;�4����wӵMh4���?Ѐ���-��߽���x��Ts����CM�����P��b7��"�5Ш���a��� !���Fl�xU2Ť���ޛ�[1�N�a܌΃U�T�	��k�o3�Ts�R�&��4#����̦����Ն�W�K�k�v7c��*/�ށğM,����`�t����\{�	����x2Ϧ�Ģ�+�:�Bby�$���E���lr��??k�L(�5Q�XO�Yv.�⇒�n[~W�ے�҃4��;j`�^�s�it��������fE{v\vAG��$?�S��lۭ�9�r�����m��h�=��]�vV�D���P�s��0�Q'���5j��p��ᭇ��W�Tc��ö8|^�),������ J~'G���'N�}��B�V��/��6��	���L�8������95@vX��U��8��f�P 8$B��#��b���Xe�]5L���N�@��v�"�t�`M�E*&,>(��`Kr�*�����~R)�'�a�.�[\���×8��^�U��x� 	6	^�
ST�D�!�h
����Ԇ���?p�e���itv������ӏ]~�@k@+���Y���lӬ�S��j�3���~㝰�/C�8�Ƅ�Isb2Fj~gK\��<�eY ��/Kv�A��}hUZ �52_eʺ���xB�)����
/�x�Ȗ�
eˉɡ���̷zP?��	�^f��ԏ�q��<�#�v�"�B����
�Z�����J����� �)T�(-:U ��$�劍�v���,�ynyYoo�����ѐ�a/U�E��:��Y��@�;�c�P5�ս����m��U,�ｴZR1�,L�O=�T���a�L��|��o��F&��M2$x����c2u��:�O4�BʽVM�,��#xZxZ����IdAӿ#��A�w���0Kh�?�vH�@��j�����2ӕ��fNG��#��)XO����-<����~��4)Lz�@2\��&7��$��ﵑ|J{�Մ���+#�����a��#(fW��"��_���V��kD���RS��)
Y_)�Eaj]����� �4�PM�B&��x �r���v��O���Y��]�5�ZvU-��a���$�)TE{W��}����'�HD�f2S��mH�D땰�����!�"2���}�EfA�Q��d]\��Ɣ��x�9�X�F|3��	na���y[�����A�t��~++�l3�i�rpU�I�<�'�m�\�#b��ʠ<������"�$h��~3WN9��mm�ꂩPtе�R{�w������(4�������&�~E0l��O� �б/���|J��䎸��f��;jR�.KH����2BTݺѣ;?D)��D�B��A:JN�*"�����Q�5,_��,��?���sq�lD�Y��q�u��~���Q�Y_������KS3\�]��<���V���}Z�*����'�Eb��T�C�m7a��� rxj�q�[��Ԃg�< ���V=��W(kߜ���iX��T��x0'(���7�埻��� 	9y�Y�׉�\�[��U��5םG��Js�

o��l䎎*�,��B$��C9���j1[9N\�%c�0����)�9LCS}��D�im��!�ţ��^��M��2?U���m�j��1�%�A �뙄�l�pq��Ʃ'��A["b�q�u��W�!��꒣��b��b"���mR+9$�@����ƽpIC|��F��3��>��%��4��X���d���m�И�����X�yZ��c%t?ʽ�WCB��dB{��o��N�Y�z	;��c,�A��v��� �e����]��.�溆�}t�ȍfS���J�$��4X�k�gNk�1��� �3<�G{�)Ox�q���}p��ntsЄۘ���s.�&�(���7�6�%S�(4c)�tbFm��q�n����3�b�u:X�B����l�P�A!��/%����8�Tt1���2o��M�l�{άB�@��
���Koط<e58��B�� �~�/�)m��I�x��j���:��4C�@�F�)Ì��m�@Q���؍�3�.0 6�lU��Lf��|k����8dUd��D�'y]ytx�O�Vz�_���&W�_p�M���:X��ە����ڊ�+��:��O20��enp�WXN�9�g
u$�s�IﶮVtA�*�$*ɞ�Cp9s��{�K[K�e�D�ͽ4����_[%��>J��+����r�J�M�.���"����xҨ�N"�Z�Vܵ��04�$:����q��P�E5��z�^��]�J<��D�*]4������]�]�ڧ&i慎	+c'D?e�&��%�� mN/-�n��_`g�UR��H���aف5ʳ�Noi�����$���@�6P��×��,D�cr�[+\�	B
�+�������V�
�(�i1�aP���Ű��]��@f��E��a�ķ?�w]|��a��G�.���$��v}3��?%M�z��tt]��6�eC�9F}�lahx;�����p�E�\h"��ѵ�Oz ����B"gtVV7.=�����/�d�-��k��uz�)�O�\+�&�Ň0L�2/|d|�n��5")J��p��2��P���i8��7m*�3�f�,�4_����S}�DR�Y�B��Q����,6g�i=+�%91�Gm�"��4)>6�*����#	����^�|���� ����W*S���f�H�>$���ȵ�=�#�DwOܝm"�P��d�7j�Ss���0j�>���Bn]A��)v�p��3+�+�g�	�!��d�͇�8mR!QxgzwX��Z��Ns�X��o; ���b�`f�`V�(ޘ�g��}zm�S��Q��f;�]�dy4�:���'	��E���O�>7NJ�9,)@b���[��ؚyDo�<��XE`����>nd/k��Z���l�^pN��'� ��>�������C�GeWL�P#�g}m�є ��)L�w��y�j��aN�:�3�,'E��M��b��.��(OIҠ�nL�9��y>���of�%�4n�֦g��Ov�
�.���!SFt�5��iε�� ���3��`��J�b�Aɪ�����R`F�ꢍ�^<�����	��j�����y��S4�߽8K%s��zc�0���Wb�«�_a�Λ|�m��w��GF��`N͡oXǄAZ���A�Kq��A�e�A����͜	��5%�ќ��J���{�4'b�Ś�jX��w{��2ei��n��5o�ə�&��S���C�M���,�8	����k��ad�CU<Zy����#��J9)$x�M�is����.#�s�M����*�7`� �7H�H�a��~��w�:�>�T�}v_�VOP��,��n�U�\@٭��;�L{�.�`�N�w����G��N�<�����]��j:b�u�� |�S�S!���zƿ ���o�s6�/����Lri��5៽���`�����Q�h�'9m֝��O���ᠲ�H��FLk�����&k�,ʋn +�!2�m�]�3FtsO���c�产춡v���-ʈŰ,����$��n ���Z>s�Ͳ�Z'w���¹�܄�؛�%��u�iZ��Z8�|�kg��A��Nf�����A���ٽK��r���(���9�e_	�.�$T�`�[�ǩ��L���:>V�7�[�`I�vAk[�|ș�,0��)�Z���1ae5_}�´%�k�@�T5���Av��/=����S]�%�^��$ke���Ua%J-ӨR7�]��e\6�|a>�ޠ�4�a�bd���c�\����W���u�
0Q�Ӧ�[�ldm��� �/f��J���ػ��8�`���F):W��h!�:�L;:����&��zGm�cz�u�����$���DU��}<����c�6��)����$%��W1���P���q�U�==5�O���9��g�q�;��l}��?��L�?��M�}Z����aZa}uE��Oe7yL0�Ȯ��������ʤXB�����)y����G
&Y�$_���%��C�n�m��,j�4��{����*�[$�f�YO��~�$�Z����aM�f4�jF'۞! i�W*��i���.4ձ>��5�;�3�p�s��"�
�Iƺ��	�K/��N��J6 s6A��G�t��|���.^wK7��.v'6�����G7ە��]�����[L��u��<O�Ԕ�)OT �a�4�F��.k��!��xd�Vc5`�,`&;��s(IJ���aE�y"����(���
��zh��.
�z�J���~&5P_s*Vn�}�����wy�
o�nEȲ��c��=Ś��#Rå�G�Zq�5`�rb�Q&��+�̎�se)��tъ����ș�$�� �����J�*�����'�A�eȒ5�f�x�[�B�f��[ݣ3�9��r��^{��:���zW����"�in���ӓD������[ks�W�U�	���otN7�4b^ b�O�_ T-&��D��6kP���s.\$��\���
��@��+BD�hp�Mn�g�_9Y/�'+�*�fy��}6Qkv�0
��P�^8wT'Vr���H���Mq��>�"�����|�n��.;]�1�0{/y�	�Am�sA{S9r�Sz����[����}�'ҡx���֯�Tp��S�{�8W��Mh�}+\+<R<=�hC�/�n7<�>w)_o/���I�b%I� �:����K�z�p��o�$�;��?(����m
F�%&R�-�)��g�M]�)��~J��1���<�r(�0����2��G�0����+U�q˱ �͚���j,aK��4Y�rۘx��2	kƹ�~]�^�d���R���^�V�m49$ �&;�����t��I�y�%)E2�&��(�"�ЯRC��ǚ4A�y����-�>�ڒ�x�A��2e�Ǫ�R�^I�h)P�����o�,�ڽ5w5Ik?�R�Qs��7xr� /m�X�Q��Y�&�p��҅���@*����E��3��FIE�(�JAB+��	c~���)p3�����ל̈��ر��((�cP
~)�ú���wF�%��d�W�������q�p���������Ｚ�P�g���n�W�oM��d���P#ES+6�H1�ta[��� ����;�Y{	c�)IRK�d|��Ɓ����?"aۙ!��r�m�N�o�-A�����X_w}'�@�����BTI�ſLdx&6bSyJ@��:�+�!�x/0�ڄ;�S���]5mt�鋁���v�h���D3d(�K|(�P@1Z	���e�'�I�5�J���_�]�v��Ŭ�9�Ɛ��<#��a����e2!~����b9W}��#���]�-�j��4PN.Cn�l����p���D�E�ӕ����m�>�/�Qf����v#x�9�ڈ`R jGu�|�2N����T�):�/�t9~��S��L�:Cn��D�'kD *���M�� 8���v|�h	'iE���JÈ!�>��N���f���Oz���Lq�@��<���'Q�˴|d^����"G�s^�U�,P�׫0�`.��Ʊ�˂~��)�����kB�[��8 �Sf��[dEI��S������f�H/�s�&2�_S�A!%��s�1v!���F��������g xb,�G��x�zܘ���t�ޮ-�6������V�̾� C1LD��|��(�lOa�I�X9Y��S����(� ���]�	�)4(�m���{�����VP�|5��^S�PU�ܧ�%��T7I9/����h�C QAʖK�$��f�eɛ�_�ܑw����Biޤ]ue�ܬg��A9��eqc�y�����gھus&��
��_�um�k�W\���ޡ"lwv{��g�c���*�O9//�"��קj�@��?n���ȸ���05$���]O�P�{�cs�֝eeW��%����>ل̴�%kC���%~�	毡h�����mZ�'4 ��я��Ԕiae��@jsp�<-��WB�����ȹ�Wф����+����,W��������yg@���c?��Z�xqǏ{�G��f�>�S��ba0�"��c�pcBp琉u7��������S�n�z��"~!���Ϸ�{�f}�sǴ�{��%�M�1F�Ʒ����|Z�Q.��-?7
Y��Bz��7���)A-f��s}�7Jf᜜hխ��Ob�zD����p����_�?�/�7���ĭ�#�ib��4&�!�P�b�R�S�K�6���)NFt2���](YS[_�� �ʘ��?�� ��%u�[,���`�*�G�k4P�3_�E�T�ZQ����E����"0�AA�Í[��B��s�ɑ�p��6 Y��y�+"�[Jzj�j�ݭ6G�Zz?9�5���5u���=����q�_�[6J6�֝�g�b�=����uk{S�uG�=���Ll�FjC�ޤ�N�����u�5�Z��~4����t�� �7X�5^
�mj���肚�|
O��7�YG?��P����q�FCPۤ�3���h��P�I�(Y����)�gB�d�<���|�ý���T-��}�K����0m;\D�윌!�q7����n��6@����]�M?j� !AUhd ��d �^�}G��~v:�+��;�b:B!��_�R��"2�>�䏸��;U�$��ӎbG��K*`窡ސEMB)��{^ZXЛa0���c�B�\��_�wrN���+��W��� ϻ��.=��H�z�o���a�{~T$��砬c�g��7p,��_2�L	��(l#֝<�Z����qtV�����W��v��k�X��L���V�κy(Bw��!�:Ӽ�@z�k.�	�sН'���ZU��R���)�A�l�VK�
e`߇7/�1a@a���VqE8�������g�,_Lp�Am�D�s_J��p�`�����������2}Y�Ԗ5)f@AET�UT�U�����ʉ��rR��y�o璯�iG�"�L�Ƭ;(ih��?[v�����g�zy`���1nlw�y��椷��_���[�)Ζ���$k��33��#�a��D���[�g��V��Ԉ��FY�l�1��d��nA�#ۻ��f����� �����@lU���rstv�H�T>
v��P���*�i���k>�&��W�x�$������jW4��|�\P�۪'c��;#� a4u�+��^����+c���f���%�z3s;ۭic�2�MB���q�?R�LR���h������R=������k�x�t*u��ji�d��[�ȅ-�r5�|ﺉ}U��q����e( �3�a\I[��2x
3���o�?�]75a?���R\�3H�,�s���;���嬳s 8� n�+/N֩�Hz1��G��ؿ�%�z�@�2�w!��U�����Tr� ~�O�g��&�oh0�j`D��t^R .B��u��\���o=:РoS�E������״,сh��Bv�[G��WS�Q�Ξ�����s\��U�z>[����ۆ@|�u'�pۊ��Z~��{�E�[��y�ւmq�k/1��}E��CB�����	�D��s�嫯7>���83�S�FDjǗ��h���=���l2�޻?3	0n�t_mF��dXVh�1&�&����\�p�-��FE	E��� �n;�a�E	��0�>T��s���S;[��.�b�D`xC�z��P�\�-�b�$6�-��(��S�J�yE�2*�h������/�<�o��ǯ~+�T�e���
N�8�I�d��g��gS�|�R��Yx���7���O�S���[#�NP��NҀ2U�`��]�p�´P��r�����s:$m�Z�Y$�;��A�(щ6�XEP,-x(A}�f�QU2Y��&^����<���.4�|\���2��.��ՕЀ��6�S�p�#��)�[D��}~
U*v��e�X-m"��L����C ���������"G�$h��G��ݺz�Rm?�}4�k�ko*T��xx��>9��HJK`I��[ɢg����%�'(�]��t�8t���w�>j���+�>�8�ʀ��R��M�Y7丹�ع#���㹑wUE?�|����0����?�:d�Ĥ��?�z�jj?��`|��	�c#L��o͙�d|5'�@��2���c*��_!�����R݉���R$ř­*AqK�#��ۺ� �	L�O�w"�\f�~{A3��(���j1Ww��%�l7f���기.��62���I-_�U���CKҜ�/C����K��\�zu�kܲ�)����=�qm/�N��i��d���0_У�8K�, ^K�q�b����qZ�J�>������~rf��cN'cL�n_�.gM7�_JLb�a�>=�Y<N�o�zb􈗗�$l�f*����BL�8�+7܋L<I�V�ƺ��˼�廱l;�_ƳI�3U9��]�p�w�I�e�)�1���Н>�=��/�����7�:��_-+�G�;���v�tE"a�zM�����˅ua�/L&�����}�I6�U���Xܮ�	���B�zg
�I����9M�V`SN�K���]�#j������H�:�����I���"S�{?7�}Z�W��>�&Ĕ�r��]��X->ǐ��Y�!񶔡��8�0ﳋ(��Q�eF���z�� �x�yJ5��qɪ�U�B��9�j#��#�*.c}���d��G�Z VE9�#p��7kT�X���D�"y0�{�m�/j��kB���D��po�^%�9�y{�� ϼ�6sB�}@�"�!��S�T[��>�����Z���kNb_X��>�3bvsP7x$�mw��n-�~3oa�е��=|�հ)=-�+Ɋ�E��~2P=�;��2��˘	s���5��P��ҽOF̻$vQ�M���Au�(��2�B������(�Z!����X�Zײ �Q.�Ft��+�%� ������Y�)��F�� �4Z�J���_.��ā���,^�ۜ9�P�d�%�ݐm~H֎��%*&�5���޸�E���2E�֬j��I֢����JPao���u_Cg�� Y���Wn���u��hu;k,������Zh��c��P5H�h,~VdĈ�F��z���&�S�&w��y�ON)#6�|ǝ�v���	�cY���ճ@�.�-.B��&�)N�-O�u��/��=�KP<d3c],
[s�R�p�.uk�'2v��e�\'&$��q-s��z��<[:�zL?�~~t���6'�Q�k���tVXG���^3�3�,�T������Q����\��l��(�=2�2o?��֑�%u��U�,Թ����\���!zFЃ���4r���4�3����;�� ��^x�<���1n��O	<f=wWK��J��=X��A��ͧ&'��p&�q�4��姐$}�Xv�Pm���ZXR5��"_���I��Y��Q+�L�.�p�`�wV���U����w�ֻ�K��w������<ܤ:.O\�EX������IJ�#���'�]�ɆLe�P4	Sŏb�ޝ$��[�-M?󓣧���	&�?r��,�h��]�Y�8l�)8UT)>Pmۯ	�T���^k�3y�pK<��gh���w�wE��H#[��)��ѕ����o�s*�ʰ00�_� �h�6�>�����ݸ�ͱ�>��G�f7�/4��鉿��T/$�9�����%�	1bю�6�	<����Y�Q?qp��
!�0{��G��M�%ұ��m�䈍�嗶�\�Ժg�F�����`��-{�F�j�OL�n���N�\Z�r�@�.��*���j0�F�;�h�@�t*�������L�Z�xK�X�����,z��2���ɢ͠%Z��@,���(��}���S�ާM�\��A��r����Ԛ�~��oT�7Bt^+�����[ d�y5N.��0��0�����_j��a	��U��"�r`ҫ���T�"��^z�h@�O4���7���>/Ω���&�dKWq*)��#�bYh�If��u�ԤvV5�e�Ƥn�z�Eb�=��3q�섬^t#��g�n�;-�
0'��R���
ېX��r ��x7	J_���j!�G�����QM�߁�=|�9��O�R��Y���/�#d�[��	}8\���SS�H�;����؏�r_΍�Tgp5�3=OF$,��h��?���$�닄�_ܡ���e�J�N��l�Sg��[�(=�]V�pzl��G�
�\Wjق-��o���An�b��ݹ����em�M"����#��ꏄ~��8��F�,���q��vX2�a��%Ƌ~�G'8��&�q�A����2s��0	�h2zX��\E;)F<R�o�$~��}}�G�� �Se�V��p;m� \�>.O�RB��¨�B�ymX\g|�D'����!v~����!���?��+�Ì~�D0<�`v�#_LNA�h3z\�,D�cHf�����9�>�V{����i-�v2��i��u5�;�Mb\��$��Sr�	%��­\�Vߢ���"��4q��P�Ӗ����v�%0���5�?�.���ړO�"�
r�wBO���i�2V.���S5�wT��"�7�M��:�'b�>bd���_���D���OJ���'S�+吩�]�8�Y���!������>8��w4IE�@�8���i�WD#��{��o�"p�m�mo��V*�q�o*��ߣ����r]�Ҝ��aҞ��׼G�(<�Y�1��\�E�ղm�?N`m�M�.��$7t��ɘ����=b;����cp��$e�a%�v�����˂��� y�*d,����c�>f`V{�9WH�ŨQb�j��i��jZ�w��e�eD�g�|,������ƴ�H<|
Po���Sl��Ǝ�7��3�^�%Y�4�/�U�~��k�V��8����t��sh�DWB9tMOTgi��u�Fޟ��|S�Y��:�\L!��}rf������-�ִ]<S�y`��B2N�=�w�ϵt�Dh�:��74����.�[�xH?ľ8�hT��Ţ�EtOW�[9z(~�9���>�L���%v�l ��7�QG��#����,.�R5�I��-�o��wn�[?g$�,����Y�f8�x����TzW#�^\�^����y��P�����	͂��h����|r����Vn�e�n�������L$%�縺c<z8��nA����bR$d��p����T�=
h�j(�����ɬxEf��{@&�����h@��g�bL�)�te��ڙ���*K��b�A@�{ɠ���yԁ�L��1�O*�ٳ���A ����er,�S��[H�Z,_���{�D�A�`E��L$Y�T�[�q0�*��ٕ��7��:Vc������]� 4�H�V��X��YfL���d�s�?�%e�f�����-C��+��uf���|��=���qEo-�7��ɶ����w"[�yl=����%���.��L��*�j�3
�
�w7�#���[nx0ۣ������1��SRJ�&��HaK,���Gq�7� 7�%���E��4�~�@tx��1�m�X��2���L_c�lU��� 0]����.�Rya���qJ��
�O���`F!ð�,3ur�o"m��Ic�^U����-D�6�X�!�� $��<�+�R�	?�>Z^ֆߪP�e�;����ҍ7E�{&�?񮗝*������&�	?����JK��F7N�(��<%l�}����Ó��6:��k<�r�]%+RL��HG��Ô���B��ׁ6���k������t�*>����"�6s#�~��R��.��Ui�O���d(����+'��Mb"�D2-��+�R��A+2��yʝ<�����v��d�Y��B6��;-vh�������˲;�V�]:ԾP, ����4�3����ٍT�~9t�l��b���,���J���'6���ci�y�1���q3&�}!����̜sY�]�q�3l�q�[��h�¥��O�)	W���NP=������(	K g@&Y�n����@5�M&��C{"�T�t�+�ڊy�x�ld�˛�E�/2��"b�6����$D 7i�㳚�X"�U+WD�j�e�A�������-���I�~���k�wF�A� -$��2��#�g�M�U8�57���{~�ԕ�����+F�a%�N��:=δd�G&����LQ����k�����@�4�ƺ���7@4��"�vf�Q�����{�D-��a���Um�Z�\�t��8���򡀭�-y���.��*��ߤ9��?�)��6�l9<q\�3�Nz�V���������Q(\g�3�C�y��n��6?����%��2��tޖ���!ZJ��F��P�!��OwB�}���IZ{�}������7�J��jV+�p&��3m��?4�I�BAI4��u�~�;RL.�$��r΅�cш,&J*��e���	�ni�ӣ�h���#{'�+���3I��v�A���z�SAN����"��i��J� �i݊Qd�M���թ�n�|I�j��Y�����eYAǵ��C���7��>���%���'�68���D%��|����X��e�46��ل�'�˓��M���RWl�,ƝW�@QvB�E��h�f���?�	XF5��5e�F{z��Z4��{�|�ZE�*czD�&����
utx�I�BLz˟݄G"����hF��G��!4�1_�Z><�s�[7Bp.w���{���-�&�n�F�8��V����X���\C�tp{2N6�qe���X���s�	�&j��Zx�ܞ�ƇN+��%�ѿ�ʒt'�a�=�MyL�{<1<��u�tj� ��B�=>�!�ɋw���?�#�"u�8�Ey^��u�R*b�P�˭���� /�{���G��0m�_�7����BZw[��^`fյm��H���(��3*c̓��R��Y���*o)�G�r$^M�
;�ۢ>���m_��͹���}�4F� K65�v
�U���4c]l���l�޸�����'�O"布�A_!��|�AfK����/���C�Y��D��!�㝾�����,���z�_tpS���.��&bd���\��r�\�`�����*9~�.:���wF�J؁�p�e��
�!�{ ^N�(�z��SMN�3�]�3��F��_G�T`䆠�9.����Y�mӷ��"�ٯ��<	�D�����_T,�i��j�	�ya��QT�B6�M��qղ���,��(r�R������9r��&��i����4'4�h�(⹉?�'P����51U�U��x�ũŤ������8��@q�}8��|)��k=<�mu�$��oބg=�u��@H���N��$[G����]�h
���D�9�
��V�1h��:rz�zh�W?tr�8�e����1cd>+V� ��X�A)���V[>]������H4�=�Y����NIj"��=�_d�,��ϻ���%�Z�� ���§ӚЭ�<���v�qKZ�x*o�O"�{�3coa�ۂ�F�W6�,���
=�Y������jW�E�]#BXU�R1�����kUm�pb�9��ey�) 0��K���+�����-�
�]�����q�JSA���c���φO��1�@3���ƆϞsk�j_��a+N�FmG$��VO��}e>�(��'}��� �מ5�vߢ4��1
���X�G��s��rі�ջc�
�n���(
��9)8�����<׳;�S�Z�����#�į��7g;ZR'�J(�|�����SOG��ބ�Px)�J���*ox�x��V��!MW�a@M�i�&��R�b��2��`�fJ�콁��XL�^@����`Q����hjm���}���!C�I&��x���)3��O&�]�c�H�ƕ���ZrTz1��}D��*qÞGT�㸧�*��K�Z�$�WʁZ����T}�P����f�r�<E��<o���ݓ�v"�Uü\�wЫ�v&+�Y�A(�4!�����>(%�=]]�o��������V����H����9]C��-�}�.�l�
|�b�����ѐ�m<�/,�ߵ�a�m[�w�1��g�1�z#s��A�(k�����˜�p���v�*D��tbkT��pE [��P�ءᰳk���[�O��~+�7��t���t���[�r�D\?����r�=�B޸��ڥI��C�I$T_�"1~�_��Ԑ/n�2/�í��5/������?iܬ���#>�p����.xJ#���S�w�.�^fV:~��Q:�YJ�];J� �ȕ��P�Z��V�5G�%*�-3$p��̆���w�J�0�tw�n��E��n���&��L� b��&�lCbik��8^(���?�^�a؊&��Q��@T�{Q�tY����mr��4����~�lT݁��[�d7�foϱ���Ex9�Q톹�����o׉}ѣs>��&gG�yp|~ǁ�i\�t�xH?&�B �&k.�"�X�wIj����/��a�����,���B��%\�"�Ƀ��)���ƹ� ��@J%��Yؠ��<K����xu�}�p�0���Wf�歡̠���.l�u'N=���ԝ�!����lK��-a�B=�
+�w�>��A� �fw։!�d�]�a � ��{��)�����۠��֖��e�	����>g�@�*("�� ~�9MB�� �f����F�-
3�-�<���C��O�	�XQ v<Bh�@�n�/��O�MmF|I�v���&C1��qJ���Gp�{�K�z�$`#,�(A`<ⶀ��<����	��q�������͟h��Ur=����x�r�"4˭�12�x�i`�ㅒ�-�ܠ�7����"��'gy�L3$'�j�}����U�=�����K/�8�����ݴ	_��x�M}����V��0:Q�"��lh�T�䦠���7�n�|I��j����v������*�F�Z(���1�/@
�U� +�Y1fi��g�<t�i'F� ���k-�B
�h_�̡�hP�^Kd��E�W��zR"K��҈`a#SL�G���>�b���,z�+�+-�rd��c	�˜\YDreL8V"��ظL��tgj�tM&�9�˶m9�r6R!*YҔ�����a���K<��0���	��]�,�-k�7P��N�a�QΝLG�$]�)�Ԡ�#L&�#\L<!��7C���Ss��HÍ֥��`;�Ć�Q���T����I�#�Ed���噉��,�g�����!��LD������Π����i�i%&H'�ӻ$�ۄ �p��.x�g�2d��I*�-�I#��2�5�ɝл� ��$���B�S���'�.�͆�>π����3�)�p�"q�}>�l�%���ٚ;��XV�@f،�P�& �� �S��2$����_�����b���
��j����UI��,�h�)j���{�H�^��<����,�0 s�̿K)�J����>O���/���Q]���0�d��5hE��o��Dn�|�^�iw\�bB�H�>�vӮ��$��iى�'Ha�t�e�-C��L���4���v�̹SH���iKQ�E���~R �5�-S�Ũ�g���4>�=?�a.�Uޑ`u~�oB-Ǎ����ߦBf|w���CaA&깨��=
�A�agYl;�<�Gc��Wov��X:d�ȳ���e��cϖ ��ۈ����w��Q4�T�lڊ�^�Wo�5>c=�S�q��9��6���3�jkc��3Q�&ޝ��؅�> �L�&�G���E��p�C4�s���j�GZ�}Z��~�38��~�-��=0�|D���07�Tw8~)��ȑ��JM<�:x�댉U�G�N�V�Dh2>X����BY���~��-8j�'\��"�Ӊ���y�\�5ƭA�ی�c`k�&�z3@={y3�L_ĀD��-�@fop0�єQ]��]P��!�t���7<K��(G3��@B��{���(��E�-�C�NX�Pg��m��q4?<P
hs'���LJd�hc�\�,�Ȋ���̧��#�Q�������e4�7���R�R~-H*�����{Uf(����u��޴60G>�=��J�;ѦG����F-8��8ty���](G��Mn5������`��
s_7'?bw,�F+_$]8KPs	g��0���C(Or�--�_La����� m�*���U 4�x{?���0;��BM�nqz���h�K'w9�f� �f/��W���T��8����Tc"�N_%3󙶡Ȑ;7_��qZ������'�>6�;R�;��r���w;��gT�ıU�@1��I�< �����f@�l�鳉���#r���+]���`��?��[� ���L�(�P�y4�Xŧi�&8W*:@��YV`~��x�v޼t�T���(�_��`��2�וz��ڞ�"�0Q�.ѐ�����iaQS/���Бa�Uw8��!Vy��@enc&^w����S�����n�R��q��2���gץ�T8���Ct�kG���Jen,��kI
���>�c 3'�O+[����~e}�n�U��Nj;��;�u�=-&�������N�����R�Dsw)����0~t����	C�H`1ck���[�3��:l:p��S�����l���r��k�E�����o-ng��rS� G�e��A�_�\]�%H�A�����P�b�Cg(F���d!���D���kL�ш��-k�4B����+0Qx��IԢb=��l�lA�0��r�'�or� ?���Pb����Jг�mb���+�x�ST�#��Y��\�F���dH$���W� 
�(��[PE
v�$��"A�� ��t�zW�!��ة���B7�S^,��k����\پ��E��J7��īv�Fž%):P ��.k��s}Ж�B%��������.ad��&9*P�ޭ#AK:���Y���+�'V��l]dΛX?�����0��[99� 1���ı�}`��c�Iv��yT���Q��@�����3�Ӳw=��=�{�l:1Md�j�����͵"VX��Bh�̎%c��y�A�֝��h>:�2����aMN��V���c�0a�DٓoP��=��Y�%\B�*���T���1�a8$�_����ze�͈����:	�͞'�wx�~g�Ha-Z�-�r50���eB����e�bt^��;��x.V>7��e��J��l1��MH��#+�[�AQ<���Ļ\��#��=5�STY�}�;����GjiQ�4q��|��ƃ��!݃�#�Q�xX�W���M�/��^{�cM8�p#$�{ 9�(�ળ���Y1x��W�o��e�����)����1ޱ�4|U �.�u%��Kz��j/�"#�Y��][~��,�9 [Ņ���:�
tj�Xh'5=����9�%C��Y�'�M�I|.p�<�8`L=�/�9��ي|A-���:����u�udC{*� �3��4�fPF^&}�/��f�p*=\�R%�6����zKP)G���vl��̮���Ŷ0�|z�^���,��B�t:��t�Q`9�s5Z*4�Q��3J�Y$���k����F��Ь����d�]�e2{s��b���nO۩�Ee
D��O�[��� ��š�o�@�JI�HK��W���K��'
c: �j���2$$r���	�x�}��QFg��r� OyA������-$Y-�8�t	�c��@6�;R���玌�a��T\�Sﵷ%��WcT�\� �o5W�"�g%^+��ěP���'p ��fiR���ۙ�'`�k��-�Ѷy���!pW�V�:/�!�1�s�q��E����AZwdd%�rbr�̓�������c��6�%Ɯ�u���X`'N����b��nj�g��[~��`1���q�:�d�1�%��8��h{z�kVF8�=��Tu?��1�=�06��3[�@�#+��e��)��f d�H��1�ޚ�zo����WK;L1���Wq�SU���Y�15�� �&!�X~0%Ӄ�F:L�F�(aub��D��ؑ�p��3'Q��I�<3�ݏb#>����-����m���m�2��|;n��ծ�%9Y~��"�r��:��u�/��$�t�CO�:�<���6s�����"H���L)��Ҋ�0��k4	Mb��&=���N]��?�f���у��ߏʽ���V¶��`�ol�a#)*�\�+�9�c�#.���g9CD&�41���^d��rG}�.������S-����#Y(�s^�S��\H8�)Ɗ��iq�%����M�3ݩS�6����j�e�L�1з�_�g��RzTw�Aȃ���@$�	�̙[���.+nR�N)������}@����5]�f	����J�Q�K�9�f�%j�N>YŁ��OUH�MS�+-�Tog-���4;
)�mJf�~-P�|�A<����]ʚ����^���G��xT1"��tuJ7Xb�G^A8m��ė�?��z�%�$�������G &�i�/��qfz�&�!�oq������bQv����̒$��D�-��=h�uaNXU%�i��o7��޾�XF�S���~�;Q�e��Up^�(�q
}O4�V���������t�1%�j�3#^}McS�C�6f�$<
ۅ����������p��6�$�c�gP<Ϋ�d���o�o�F�-�x}}�����2�`��� ��u�k�ux4kZ�Ǘwj�-[��6�������y�ٚ�����hԞ��ܫ�EcYF��"��1���F�J��7e��uPT��E�p��\w!�s�ӑ�zՓ}45ZX"M�f�e�1���91:�d��h�[�����7�T6پ[�>���E�d�W���VΡ	wœ��D�\'J�7ko<^������]f3�̴���&���Y3���Y��c�<7	i�m�L1�dҠ�VcbjF�����s�%3!�I#�0(��N�G�1-En� L��=��j�6��à�BqgPWvX��Ǯ�"�[���R���Y,X���
slAe��KV���Vl\������z�)"��P�{�v�f�a%��hx���i����@T�ʷ'�v��m�W�����L�<����œ�u̡�G��G)��7��IK[�0�=f���,��5(���$!/tȾ�ܪG��%�H�KD|�i7 ?�6q^�.S�s��٦_����g�h���1��:��l���C��l�{5��b�L<m\Ć\�3V�_�ݬ�����^%&��$�Y�㏰p~W�����ۥd��/��L�wp�_���E��T��>���x=��Y��IHK��\QՇ�)e���KhG8��"m
`H��X��C�(�5<�[`S'�\��p~�Tզ޻1��q��싫U�Y��VPe#|�B�_���Q�o������
�Y�W
�I2_�Ol,5�p�$2�~
��4|���_��҆��41t :��tMB����Tk���[~�Y3����MƄ�L�/1(��< ����u�^���m��d�Ƒ;��S����j��r��%s�V�K�
�'@�lĤ���!��u���Y�7�$��r���!�����|.a�oJ��י�kc
H��U��`��8!�Q�XV���nz��@*C�[ۙH6��ה5�Uܦ�-����|:�Ė���`����)'Ӵ�.���t�N
�ӵ�P��M�t�I�X��J�(�h�2p���?�h���f��MD��-�)l�\��1�JW)��۩�"mó8���T��)�5X�1��8�P`���Kq �R��k>}�1~+)�Y�f��Q{{2�<]���2p�m�ݩꀞ,�C8��j͓���u�=7���Jr/=0l!Y2��$Ns"Ú������Lbˀ���=U�&�N`���<�#�؄َ��%���'H�:#���ǲ7�̼$T�O�5we���Wc��w�y8�Y��f&+*!K�>A�a+4������	��|�I������3�Β| ��w���LvD�ߚ$��RYbM$�!�̲�*k������������"���F�7�WI���y:A�B�g�a�q���ߔ6P71�D��ϔRup���35\9I����0Wy �X�x�������9B��:�K�3g�*�g���_.Z��]�/����I�������)��i��
��p��̌|+�X����lp�fy�T&�lv!��Vx&Ŀ=�?������wp�'pl$\G-8w���e�vnxH*y?�,�Q}��FQ��(�oH��Au��*�A�{f��Ť��?���i�w�v;��
�㦺�^aQ�����4�7��̂ݳ�}��(ه:@�0D��W<W �֞��;�U��"P2J��֥�H#��5��Ye�v-H����<t0J�X�����#� �Ge;�܋n��@�R�*i_п��� "4�mc�H%��M�`�i��y�l���(��P�Pƫ���w��/�gWs$n6�<��/����(�O�C(Z� �B9��N	��70f��b�r�S ��UHV�E2�3x�,��ƾVȟ�����l������6/�y���O�}��
9�����>�j�.\�%��<@#N���~�"$q��?���h�`��Xf]�J\w�+wQ����T��U���S&�I�:�=�_�"��,%�\k�Ce�:�7�tzG�����xC�S,���0W?�+n���J��<\�E���á�Ǣ�;�j���S�]��e+o����'3� 
IP���wg��G��X�ނ�V6�{�}�*G*�TG�Ь�}A�	�|G9�թ�f��e�cc�#����>���źYlI�s�7�a>�;�G$&�d`�9R��Ì�-5f\}EIt�a�Q`?^����e���Hw�����H��dZ�Hq�Vk5��\�ApQ>�t+��
�24�O�o��$�t�)��|�T�m��hs��'U�3w�s<ݼoAH6[>��!.��h���D����1ۏ��M�����N9��}��=�y�@��
i��\3�r��z]q��sD�e��9x���b��+{&S��E�>M��S�@���!�f��M����u�q���z�D0�=�rf���Q�|JI���)��;(_��ൟK
~r�-,��Jh���/;z�ץ��Vx�m��KYK�P�՗�̇C�i��b�!(���?(�Y#� .���ђO���1]!/�巄�Q,VRp�R�ޱ���+����J��uq�:�o.?���@*J��iY�Ҵg����Y�]���}x����1�3P>ɗ"�k��1�/󎓘����6\�m���Ey��Wpi�����k�<x��ɳ�]�F�K��#�����v������0=�8����- �W��d��I�F�uy!���0ikh�x�ֳ��vw�=:Ճ: �"HB,8O��݆��=���\3�N���Oh���↔�O@*� �� �uz�C��^?�)z��lVbCgfv�һ-D�,p󧪬୊fP=A��o�i�WoK�88O|�M���(\p��UA���ș#r��چ�0��R�Q�Q�Q[TY��6��ǊX:C����|h�\�Sgq���BV�?�@?x�D6	Ǎ/AX�cS���fŁsf�CS�Q�jcS:���6�ܤ/�"�Q.�{k������*��fU����g��ySi�X�AAe�|�(��{��?�0}��+3P��0����6N҉!�{�Q��qn?b4�_�Y�Kh<K�{�!��z��
�)5���k��(̀y�P$��F��rl2�CbĈw��:]�Ne/��a�7��e�7|���~�n\</�O��z��ˊ+%��FL}:ח�i C �-]�X�.:�ӽ�Ȫk|��	�z���W�%v��⫰�6�:~8,��>0��i�E�%]��:׻5�s����F�a���M��V��e�PBbR��~y ��gb�o�#���
a����i/�Oy:-P�0)���iq���լH�v	��]�tTg�����6���Whw��OD	J5��dփ���m ��n�'��.(UR�ٝ{�f(���$�m�Q��]E�\�	�|th�'ko�������e���̬��d,�5W�� i���!�jD�V�0!��3�t�.�jv�-O��O�2JU����"�d��Zշd���-�ϊ�~S�P�d@<m�,L����%�e�U��`~4$��C�w�*�L�@'�M���<�Qs~�s����V�G�?T��s�zzp����6Jl���>��8�O#��M}%��m�T@Q�g/ŉ���5L�T9[ qf��%ڲ�p��\���m`�S׏�~pU�i�%���X���2����ֵ�d�Z���`ぇ�����i�^6L��Q�r�IZq[�}rq���|���9~R�\kIϊ���lp�d��/4O���A�[��M7��� C���?(ב�*[��Rc�bvq��������|p��,̋� Bs�S6�B�|�+r��jLu��	ܡ��W��\��+5��W��
S��(
$���ggb�|���c3��f(:��7%��GV��+ ;]�[���(�Y�$?8e��O����4��^�E��<�?su����S�莣��Yb˾�c��ܟjRQV��$-Қ��6�aC��h$��Y�(*��k�B��4���������m���Iڀ�P���Vs���7��_��+�)k�u4�k��0��1窒~�q�7�p)�i������GPcE=��!�ET���__��-0����H�W�����<d��|=!����}��&�~\ �9�������sY;u��u�х���>�B�dUw$IR��`���TF�s-`"V^�A:&�v��p$F����v�_P�4����>Mv��A̛B���j�)�t�S}
5��6"�2�������+a�7�P��ΆF�eN�RI�$`�9E,.�[&܊ ��8� �Ux-����ge=֏�fHn���Z����VX^bnz����=�~�������F�lh���ų��B�̇� ϱ�ڣ��\Z4�y�t���%��{z9B2�2r���9�X<�����F�h��<�� @�aoRּԎ;CУ1�PXO,���#K����F�����E���y�u��Pl	��>6lCHc�3�"&*�c�	�ć+lVd[%/.)_��X�ޞ�����݅L�^m��L�
Bi�{�Dd��P����O@�[k�l���nd��Wu"�Ҧ�P��9aR?��L}��`\19�4~N�C��JZڈ[&H3��qMn7���kW
2<<]�b�8�c�|/*G'\�sF�
p�e��;���g��oa�G* a��3M�t����sN��<��,p ؒ�|�����co��|�=�/��EԢy�	yz1�$������!�V'��'/1 ��#�l
������ɛ!L=����Ċ��*V��⪓m�넽��<<��Oj�mmL���jd yޯ��N��u"�O*�Ћ��2 ]K�d�.22��C�:��DiO�n�Ҵ,_*/^W��S�e��B�5�䪨�zD��<��'�xcm�I�D@�����Y�j^I��~>��1`/�VJN;~ �4
�a���&�؈u������UA���-q��{��V:�?K���ؙ�6�/�E�wGzs��^�����>�quŔ�͌t��B��"�Oe�Ϫ�	6��%����8L��j�N�N�#k!�/,�6l��v���7r:͗ҏ�*���{�w@�r�Ak��l��;PvuHuNdd�d\x���OL���]Ef%���f����7o�&���/PJ?�7�����������0��B☌�ϥ����L~�Ӗ]{�@�ɭB�	��R\�Ʒ�H�J�u{��rbY�S$wJ)ǽ�G�{&��1y��8�ʖhߨ@]���GH�p�W�&�[�f,�Ni���U�M��#��!�&�D������������Ǆ�adg�:���#jn�{y�����9E���x�(8�R9nw�̥BV�܆�D�7(��SM�F.���n��%q��}��;��39�l�F��x����~+K0�}����e���܇"��0�b�	�eyIC��#_c-�ñ���^Qe����SnK��)|��v��2T�d� 5ߢ��O'����Ce�	(A`���H#��
(}�K���d�O��QW3�C��n,��,! '7AE<��G閰��3?v��~o�Ϋ�d��<�#Sw����q*���eu�a�������0R�� ��	���i�7{�#}��Tg���I�l`x!�|x���/�|�՗ݯ6�iT�Ӈ|!��j2_�e���p�HᵓO��֝y1����%M�/<_Cy�t
���f��<�Ͽ�wX>\��R0�#�K��b���)��{��	\R�n�>J4��`� �c<�'�x�_�ۡ�Q�xǷrAï9Ӭ�S��`�)p�+��N68Jm&��&D�
[�w��/̀v8�nE�r�#��c� ��Zk����Yl��ܱ��X��8���#�y>��l��\n�ͥ�?C�oyNU�%��	�ϢDK�.��gƓ��wP��	�p�/�a+�i)R����J��_	8YrF�Dhفr��^��s�fW�㬕�&u��jJ�J�IW@��L��Oo���0�"��rsm+�A��t�p:E(.�R�h<���oճ,Z�f���ѣ�	�����y���H}WsT�a6:I�P�0����������ʄA�I�K ��,ｺ@��&��p�o�H�d�d?h?47��IoQ۹�~)=��.A�L]�n�'̂���P<������L�ۼ�����S�S�l��[�gyx,�"L��*��?,�я���I�(��l7R`��d/��֌U@.)j��7���:�1���F���Y���1�Ew��0�RO�n/�A�SƍP���i;��G8�&���q�ͬ0B:î�]�&^�xr�h����=���.b�2Y�ݞ
.�5��?����p���{��Ie8�^�jꩄ�J�YWҿ��\VL�
Q�9��0M֦6��v%�{ �U>Ǯ��J_l1��.���= 34|T��:�5 �=�}�ĹX�}��ӂhL3������Ӎ�:�b��n��*˘�\b1G iT��l�o`� �*X0�Tz���
TѨ�fqB��)�ϭO��hv<��|����I_�X�P&gJ)�ȫ� s��o��תd��|�:��y�Y�ڦ<�|qk�����D�"Sx�H,��]<[� �q�\͢�{�O~�t��H��W�Hbn��D���ש9i
K����7�dR�uc��
?�i��G�g`�_��0>;�$N��@��	�=_����9�@��`���ݔ�N��^�g�,xZF7}�]ыж-��+\��{.�7�F a[:iI���u"�'�tݢJ1}�u��Qj�����T�	�U��Ejm�ٻ��o�n��F��~>2�q{��ss5`�r����;���쬚ǻ�6��ڦ<tKX�O��p�y�oq��+���텍����>8u�(y�n/���/�{#2V�����1�~����w�]��Iw����@�"l�C3�dyOf�3H֣��$��/�M�-���f۶
�]ŭ�8l��Uʄtl��L�ղ�	h���foB�Dwt8�Z�s����G�+;v�5>V"���*�Z���Mfi��U[R�������4��M�+�U1��$4�=�%Su��]8'�79�?��� Ŝ�{���ݍ8������lJI�-���bHuT��5�ݕ&k���e��񻼪���9�� �%��|N̤@�Ou���=	����.m�k��� []�d[S��oŦ���V���,ҧ��&T}-Ն�t$�$��ڍ�S�eTa�Vq�p:������"���H�P����{]@9Vj�#�ߑ�*�fz� I�.�Eɑε�p)�ծ�J8�!jx �-+�0l��o[�L���4��4�Q��L�@�Y�%�w�����0%lJ��J�*nCF��!E��E 8���y�^��z|�0ޖ��������)�r�Y{�t�y�5@�X�c���[�pT�mD9�q�+Ě���r^�N���P�狄%/46���i0g��~5ATQ�����)�2!�sC�2��"�뉴s���u���7��Ou��q� jۛyt�B��M�0�~�t�׷E]P�$ų�;�gY����M���G��K��:[5��vX�[=��t�lQTg����������j��2k5Z��t<��ÏQ��7 �y{�ځk.�c�U:��?�Hͻt��p��m��eZ#H�'��H\�3�S��p�E��rXo)=:;�u�u�I~����,�����h
���O���jB��G$_Q�Tx,�	މ[�
����ѥw�؃$��PIw+/>%��]aZ�)�9��ݵ���v]Y8G�r�VF>���AY��}o����<i�tZ�r��%A�&ޭX��B+�-K�B.���-q��� e���l��5�����?��$`K.�"W,��S�GW��V�ss��W�Ҡ;)
�L����l5�=����,��m��^��fZ�]����$�jN��Z�sc�i���]�?̿&�E�����ܧ�0 �&pdZ�"��(u���1��P��n�6,���Y�j�*���#t_1��^�Tܑu��j�V�;���TZ����Q��VXFw�=�ځ_�>�s�?��+�������-�M�ű����l�|�,
��(�#�:�����w��lC��S��=f<`Zߖ,q�W+�;U��,i*/j'
^�1il&��}A���e?ã���l�B�w�AS�5�!�Wo�_���&ˍ[䒐8~�7;��Px}(�8�Ӓ�d:�-* l���	W�����&x��H�sg>�;o%g������";W[��j�6#��};ܺ�~�r��9�z;�t�?�
�9춬Vb����*�, :�]�nA?G'����U��J��uX"Q�v����Gn��7C2���q��ƠA1&"M��΀�K��1Pʠ4����]���8���8��!8��X֙a:���w)zNY�;"EUE��ӻ��g�\aj��T�B��*> �0 ֲ-�<��ڽ��P#�1л�X���`$�jj��F�1���Nz&4�vd�H��⫉�ыL,Q��ƀ���8��V V9֯1�J_������Gd٣؏e�
Q��2�4#E(周x����������A�]��oN�R���,�]9�a>�����ܤ������jd�ł��:ih2W6
p���[�
e��<��b�l�]�K~��y���B�Nf�������_*I<+�l<@�X�(W�:PH�KP�NIc)�O>f��W����n�)�b���vB�P�	��Z�P#��^H�	�Skj��l��B]�"��^zWn=!�{�Rj��Tl/[�Q��D���)�wjm�1���,��@���0�U7�?c@��Q�؉�"s�/qwpul7G[� is��CE�Hv�� ����/�i:��J���M�"�<9��BӤ�Lp���v���!����y��z&�������)���¼��A��5��7�����ۃ�g�w�њ��b$�J����U�������������P�$Q��q�Rͱ/	Dk�$F&�61ԇ��|��Ĥu�^4ϱ��V���V���	#�:�W��w~�����d�78�),s> ��57�+���2�vc��?���:��V���ژ������G�2$��s�V+!�=3W~O�"����Mꭈy!�%٥Wmς��Bl>@�N�~����e}T�k'8�:/�"������B�R��Q���y��m�/�2�h�`j6��7痺q<�֠�f�w9�r���"s�V$������%Le�_�kp�C#G��C�hg�վU�%���8�b�"3\�B^�p�ohΨ9-#�6m^�¯L�`���@V2��)��1R��S{�6�a��C5�$���J�.	�D1�.���>�c�^K�9�3�\gԭ����C�x�J�����D�!��q�%�p���-8��ɸ��L�1�HQ~?ٛW��:ϼ
���'gU��N�q�␦BH}7t�6��<��g'�k� �a_ɟ�h>�JC�nU�J��8b�|VJDb�yj�`����MW��ty�%�h�V9D��7ヹ;m�/���D�_��]��������LKW��̆Th��aC�y�#[�+ڊ�WP�hj�� 
h[:��'�W�(k)�`�x�c����S�#+��q��KGG�e�3�y�ۛ14�b�m���w@r�����0 \�D�}��q�~�;����~�â����Z
������8��jQI2�@w�zRwExL�66L1{��;��K6gMF<�i�(�^2dDB���bX2��KB�,VS�5��d4�6⮔���P:��Ke[������ݜx�A��[��h\�h�y�x_E��xr�D��oM:ktE
����!%[����̟��Q�}ܩZ��fNc>�����kJZ�`#aJq��s��RkT�a�t��0�:�4J�uY������/���=�����" h��R<��l)����<N�DF�;���|�/{�|�� ��\M�Ah�ˁ������A^	��+���8�L�gi��Q��=����32�F��s�vM]u��Ic����u�C!�|�	�4Y�RF3XU�P2+Q�J�������=6���uO���Ǚ���[➥�����P4Զ#/)t|rI�"%�H��y��bR�r鍾&)�$e���V	�iD�@H���F댐Y�E{?�Qo|�����A�j�B)���� �ra��r��؆��Zr���bcDPa���M�ɘ�Pg�(�pvE���o-I����S�����)����eik�CUq���Z�P���܇��gV�%ڃ�z�w��u
�a���Q,Y��j��
!rX�=�>��q�3A.~����9��t@c��M��������ƴ��Q�4�������� �x-���Gb/X��&��O�6��˜���C9!��r,�1��۹�9	g�XKz�'���W�W8��,��տ�9�:o��S�uXY{��G�쾉�@@/��_��<�cb>	:�$��f� �Fi*�� [9�� ��S)3Cܠew!|��Di��l�e ��p�kӜ�U����cT0~0=������KE�X�q����D�^��7�pA�U�<:U�._�h����A��QxS��A���n�7�	�U��u	�#~��Q��I�綽b���􁋚0�:��9f��q|��,֍���Z`��m.��U�I(U�����o�_Kت8x'?_m��(>�������(B���K{�q�LN�Ŭ:�c�G�1W5�ߦ^�kei�� �O�1wNўw����Em��2L��,���!˩�~�����7�c\�P4�}ʊ_u�."F��\{�Ԗm�DP�o����Q?���.�hzpɪ"G�Ϊ0`;ͱ��o0�$�k�[��af�T�-i'@�>Ʃ���!�<H!I��`	�M'8j�A�j�~���OY���t�0�ǽ�f|wرDq���jX<�5�K�:�v�p@�ЈY��#�R}��ˋP]���A �����)�uh<��h(��G\�ҷ����}��53�(�vlG�����Yv[ع|&b��I=��b_{�/U{�A8�ψ�X_7Bd�V��:8�'F����ܞ�t��ˡ�.mf��RD�����J����N�П�i	BBq�L��o%l�x��X/p=�� 6��D٦��ʪ{s��=�|�����MEC,h��/^m�]L��p�!�qP5y����y��#�� j5��3ц��A�p�\J�B��b�����օ���)���9���>V��azJ�?U;�5��[�����,�J�.3
��4_@`�f��|��'���Yi�0q�y����	�l�E5��Ǔ� OϽ7\�:����]��,�ϢL@��Ae�������m��ip��`���j��]��m�{�:_��`XCG���ܻ;T�������n@[�)�,��&_�¶��6���e`���Ч8�(l��Mt���/T�kZ�9G�P@c���l���vG+���˭�p�ۮy\�F��U:O�͸�S~L�{tG���`�gN��_�O�<~��bA����xfc��1]��_� 3Mb�i�axI�hO8J���I�{���;��4���o�
�(�6�`ܚ)�Mb�,W)Wǯ��`���Gq6Q��/�g>ìn�� I���؇�q�w���g]�����Y%Ph��1�_J�� O�ڳJ��j�3m�X@��?�����R�l�G�"
�fX{RAx��	:P�ݏ���z��XÅ(�P������%��̐�#�/������XCK*ʻ��M��t�-~��8M��ed��O�D"��i�̲ArC
eH@1%�K"�n��2���'WBXY��F8L���-}BM9E!	p^�ۘ�h��߫?s(�\�;D�i��q�K�Hb7>\���kg(��hb[�+���1�]^zZ����q���-ZL�Y\�a��_@�r_k&�E��K��銊4��71�_�����G�!�0�0ܔ�����U+��=�����Ss)���z�$F,�W�-��ʻ2�H��4�%ih #�PO��X?K���?^�{N�^>R����`���ξ�J&��f�*ź"=�2[+��L�@bea�b��YP�"/�pB���f"��
+{��Q{]� �ޕB���QO�Bjs����~�lH�E3夡_y{fWo}� ��ɶ�P	�M�.��z��_��i�r��5_�O�e�ǘ�2@��BC.1�OF�:�;S�D�M�V�j ����3��������l0�}lV��݄�Ts��(K�ɪT9�FZ�~��}\��Z�W����?��'��s�5�w t߶ؽ�2��d�azv���Sn��)�G�ų�I{���� S�>*u��r�@-Wvta5"�]:I?�}��Vm�J� ��4�z��	�D���fP�ա��V�����[�b����O^ ��(Ǚ@5)R�]P}�&�	ꕁ.ԩ����8��&-�����1�����
X�>D72^����	|�e��ո+�D`����ǧI�E�/��ȝd���1� [���X���L=\��d�nM1�0E�d����Q)�1{�a�e����\O��\���q����P��\լR��Ll�H�v�.9���͢���m�FK�Yr�5="���aTI�+��+c���ƚ�)ɱqێqgwӛ���nWËe��_�	3���=�k�Q&���u�-����ش���dLB�S�F���+r@�� ��$���@��5lt��KYW�m�)�U�;�骴�D�F�ßv��p�4�Kﲖ";G<V�;��GX���>��D#(�#��V\٘k�d%D&�@%~��h�s�l%���`��tX�,3?�c�3C>X).X/��=���)Sx�|��I�Y������#�~'x��L��[d����F�܋XO�tx� <����^\�FN>�6��i/�e�<�b��t��1+[� �PIFo\�.�
=c�P����2Pم��$��,�n�3�.� |��T���W�/(�/����e̶̐�\	2�l���DS��=&[�<���j��/�',���fhؚ�n�[���F4Ú��X�4�dABŐ?yE�L�@����3�C��PHT2�hF�eoR�� )p1�v9���,�9b����������-G����y�3����κ�jy��XXԤhc��C#�6p~r��&Ϡe���tC2LVx���k��L�I�n�1����R�)�,��8�Wl�H BU�֠�r5s�'�!ge:#����M��8�bV]�5�,�h3��n|4.��Ś0�r��Gк_:���Nr-���>��(nM9���'���|���YVo}�`}Kyϻ�b{(1 T�I�4��d <*wu��|�{u�3ǒ�t�\����{LW���z��B��/�@��ACQ[����R�f�4���ioVWMoK��46����t�� �6����W�EX$��i.]����������Z}Ovm�Q~��tS	���#Iܥ�(��
�E	<g��:�h݀7�-ʥ �/��O
��Ԇ�Y���䠸����r����w/W����1�Z5�����q)��9,��i�����NZ�@k��A�+����V��NL�=ɡ�^��`�*�����=Usa���O��})��TG�����=�r���|n!?f)�.��]^�;�f���6�z#7��`�a�U!��<E�.AYIA�5~��s��A9��3��:�֩��|��|�����"�ޢbS�.����`^��m�]؇�E�ÿ�
���J�(�{����HC���D���vZ�8�e��B&��o{�yq�X�G\=�m�7�pՕ/�_Zj�:�$csnn�qh5]�R�-'<��1(��]�yo�>=֘ ��ҽ�>]�=�lg�X+Q�oo=.��:�௑y��1�_*m��b��pC�7�(�3k�� >��������;�m���s�\D��\�z�k��0$?\}�S���~��&���ϸ�X���5�[��%��E;�A3�Kb����<�ڠ��P7߻��_��Ś8\)2�n;4,Q���Q�>�ܿ!@Cq��O�B��Zo�O�$�"��S�(��d����R�ǅ3����>i�x�a�u��R��X )C�r��0�=����v��:���zr DU�`&���b���j�c� kH�
>R�j�C����*O�+�Շ�����	Ӣ|�ֵI	{�u"��ᕄ��Vc�q:�6`\l�P� �}N�i���Hwd��Y�5Z��f�ʧ�G 5s:��-�8���u�hּ-��e�$�'�;��[�KP�����m�j���_㱂��jp�찥����(�j�z�|�a�mh� f��Zb�Ӡ`Yc�&<܇�hˣ�Γ�ш~ *��wR^7����`k
i�������y��>�U�͆J��R�����fX*T��ד��	T
�� mʺ�{��8P�(4�hD�Fa!�\0��e����h���@#�%��i���.kf�R�Fk��S̤y>�[�89.���^%e2�2B��9d_m��~������5G�|�H�(��%�kS��	�8�0Wo����}B����W�4k>.��]C4V;�k��Q)Q2�-�O����
c�Ȼ���> ��=s�uK��U�q�X&�A	p�#u2���,9�碰p�l%zߎ���fGoR!�_4p��߉$�J��#�5�S��B����a\�۔hւ��3���{n䮅��Z��s�(�x�����Vuc{\�C��r���N�x�H���V�)N�
��6�\��z�ܸ+���0�C��4.�A�V��A"E��*D��f()��v��s����6"f�W�m>�~9���C�.al�6��&��&��R���
�JxQ��	9� �m�+4���"�Ӣ���I�0�����jd,�M��fޠ����?�+o��	v�,�޴�r�Y�"�PJxBB�'sҋT+�ߞ���.�}�:6����5����E�!�.���������1�V↹� i�=ֵ�yu�����78�?��zӬ�2Vr�����:G��������0|�������;R��vV�1�j�8���o�g���S�3�P�ATx��tDv���Kl^2��,[Ep7m$�@�
|�A՚)� A��J�0�ӷ�� �.��;#���'�~ӆ�*�4�֒���=׊ĬƧġh�o�K�qh�3�Z�w��Z�H���"��>��ڷ˳�����Gk�ʉҸ�w�K��ݻ+���/�^c��x1��:�ӡI�w-O�h/�9��:��v� ��Xn��ߚ��>v=��f�5$��9ʕF:_$���$����v}2�}l�~h�x wm{JݪF���~���2��:b,�Pw���tLj��t\��v�m4���3W����ʤ�K�倻�qM_�z�Y#�Kѥ1�_^�|�=����}��� �E5�D:���ȇV�>�0I��>(��K�*0����ي���,Q�=. =o:��3��:����&�F�E���x8�*ӊ���6�^9�P�I�k0�{#0T��z�՘� ��p-Hk@:�r'���K��I��^�M��ٗS�V��<��p�%������s4R+P��6UHԦ<3jEw�tl&!������|>�����DÀ�⎺��>kf�?4p��WH�p.�B{�����v����$���]���iwƤ
�c֮*[  �� �h	�珎��p�꒻nL���,�����r�W��Ъ���
A���8e��������H!��-�\� �tD���9�Yd1��x������ʡ(Ia���!�w>�����#-�n�)<�B�~���������e�}a��d��ɐ��X_N���ǠCIA4�Ox?H˺�\��żuF*� Ў��uDz ��{�qf�-��5,��)�r�[�{ʸ̥1e�T�r �x<�{�q[�Fdb�dv&8ZFeV�������u2�K�=�ńJ��`�|
�O?LӬ�m Ǟ����5��q�}�u�{��mj�2�懘ZR<�/�lT@���~fݒ#���h�* �F�\�O�=�{���k��#��{�'�4�6���.CͰ�/��.��V:{f7������nzwm"��	^�}��hЬz���F�l~g>o,a {��4�5�Ĭ��
\*�4~��]�~���qa��ms&�4p�1� /$}+�+��rq�����a8�0�sRљ�t�o��R�uCg�{7ڢ+�ڋ�<�?Ba#�@�4k U�,�!�={���Ƿ��*!�hֿ��]��:�s�B���U 4a�ɧ���0#�"y>	v
�5��`��7�� a�o�>*y�<��6�NÿLn ���<�C�z�� ��e������5<�q���iz኷AN��t��#���u�r�{��?����h�c'"��6�,�ٜ|�?5+{���� (���"��=N�Ϊ��Nci҆�|�j�F�F`��I�8����Aq�����0�Ƴf��^�߿��Wy� ��W���h�u�4�*ɦ$I�	��~�/4�"|�"�\P�+��]S>�J#~�b�fSV'UM�㡡��v���`/Й�ɩa��ޞx�J�JJ�8f�#�+I��o�WH6'qtO�|����7�h�@5�A:Hj�R���b����~T�8�����Z���S-L�7��s����OT�2h�[�1B{ɪ}�����5!��Qc	 �B蓺�sǢ�m�ڸ��J�EA�&�6�]k�i��x��;ViuʜwVS-蝅��$�^�V�R"�"�5X�6l�3i�+�b4c#�1� �-�x� �u��ׁE�A��-Qs�g�)�-<̚J��)?���ٛ[�K�� Y%�qh�ɷ��H5�;ml�.���X��M���G����x���{+
���ao�v�2��No�����`��4����z���	��,y�۵M�Éځ�(ѐؐ׷�+)4<H��O���a) ������v��=� :�B.����'��9-�!�c;��餅��c�k.-4�@��C��h
��X��s��)�WZ%�W��Ҹ��Yc$�\J��Ո����;9��}���q�{R��%�c#c�kri�v%��嘯�o����6���ߎ4H�k������[�uڳ��IG%zKw?���/�a�=��>Ũ�n>�	��XKk��� 1t`B�J�<�q�� P��Ow����ؠ�r���Tg���x��eU�{<��;�`����~����SY�$6��6/����Y�i"� {��hOq9�,�o��i<y2~�L����*�Fֱ7�xe�@r+�Y��K�:0P�YL���l^W�@��8�-�.b�`5�-#z?���DON4ǵ�Q�(�8�t�a>�c�z��?i�|����ZFZWv��{�'z������^1�pZ�"�B�K� ����3���h1�i%F�^͕o�`��
h��U��F�i�tS⋋=t�R����:�D��&��?��u���h(�S��i��#�鵢ޕV��)Cmf�+i>���T�Hg�3��y ��V���ШwH������v{�9<�i/B&�uff�Kұ|Ta2e�k}�8T1�.��NE��IhdJ|�)�,�n�;����0/a��z��&���E��q���N��R{�\_�����f�R��j��W_ޣZ!�噞Iԇ`\9l�� r���Xo�����%�m�J��	p^����'��f�1��� Q�y�\����[R�Z��z�)�F��شDQ2�p�@�n���1��������N�LzX�N�6���O`�ʖ*v?\ 6��4����|��o%�T��
���](-��I�B�����:Ny���Ns\���!+H��|4e��O��F��c�~�"�����_-�e�2�H�Pb ���Ky����@��'����{��O̬ ����I$���.���}�l��J8��3�R����GqޚHԚ_��.�m�C4r�
G8�;0l���7�b���}o����w9������T���B�+9���3�s���%��j�rH"6�D(�����Ĵ8�5ݧ)��s�&���dH�D:�,�)�|�i^R�"Ƞ#�?�6��e:h	dx���M���ede�,泡{έj�Kx���ߛX���#����Rn��~7ڬ�a�EG ͏Έ
�]��|}��������~��-Kg�#@���R�ư�J|K[�=�d�ƪ�U��M^�����n&�}���x̻t����a
���ܰJ���\��� B�\s������d"�)	�����U��ސ[�� jq�$��MB,�b�T�~�g�c���<&B�+��C���;�ٳ�$����k���p���$H&8xTp2�>Z�SS[���Hƒ�H�x�8#�t͵ȉ�9gF�ha�[���\-}���s������y���+}J�P1��*ؕC��o�5|#��0|I�	� ��є'TBu��ΝR������;��3����l���/ݘ��w�;�4ҾO�63�$F:/)aI�l���[RN�,2$�y,;��
��X��#n�A�����]�(
��3*�9�]\�@�3�E�u��a����4L�br�r_��7roY�g-���4��(�*�E#
�XB�]�i����Żm���47���R���,謶f���0P4r�虝l��P��B�����ʪy];�\���`N�"^�	���F�*A$"Ղ��S���tq��DB;.�N�ȴ��_Mo8�v14��ѶN}��*�fz��v�L����)����~l�7��I��w�2�WF�o��4�͌�3�<����9���?��>��?<?30����T�ڭRK<.׼\���1�.�[�l���/� <>��#
��4鏚D�y�b�x���_�v�!{�����o���h�`9��Q�zܷ��` ������6�����Qi�>"@*�� -z.�a.�l��Y���!E���q0��f�2H�.{𼅭iRxA��l^/.�2�!	o�������A�OR�L�;e�Y��4���},���W>T�
�t�P=��"e�`�����d�Z��0$z�H�c����}m�wa���ʀ�/_q(���A��Z�Lt{���t�8�e����y��Q��6si[4,���]ÙqBi.lY�Ս� &�͌��V�зDz�ELc���D�职�/�xFG/�ރ�>9�T#��G��M�a�0��Gs�t���Ҳfϔ8�'<��e �� �������WU��[����m	8��s�,z�d(�#~}���IpZ�@} ���֊�܂�������္c�+�ځ\L���D���öZ����#l�<�Z����P�����r�(�!����mgƿ��3��-W��3�sN��З�$o����6�t ��!|�5i���/vxagȇ]�'���BHi �^�V��@!��Ȇ��U?���=:��!�U(�G&��ק��=5�w�:ם �i'�Kt@J��e�鏳�㒲�ˍ�U�� ����or�"�jM���hO ��G�S�۟�Oۺ������Oڞ���C�a �έ��~g��!���	�D�+��Eg�)ahh&��ru��7��^"En�^��ͣ1���/�����Ib�%��^�ũ�S��]z����D�ލ�*E���=�� 0o�������oջ�Mdt3���Yjڿ̊)����J�AË��,\�"m�&�H�)�f;?�j��Lo1����V)ʺ��+0o����N�{
�1�U�B1�f0���~��V�F�zB���a�?�23����we �gt���+I[ۅ�"��u��j�Tη1��[���=�H`'��J���\b�sZ	�C��%` p�>QNō8!��̟���5{跛�ia���\۩a���>����;J�u��MpT�Ƨs�\n��A3\��|F�' y
@��u T06p���L����$�O��B2��Dͷ���8���^p�"��Uvl.����*�>��R��n(����\pj9��[d�;��)/�+^d*�
F�����{��,J��n�ӷ5�6$���K�@$����	o$Z�F�$&0]�����t{��6p�/-^�h��R{�<�g�o��"�^rԝ�B�g5M�[�8�Y?���F��4IGӁ\�*>Qg����~��N	B"r�گ���!!#����«�a���;?E�2�����VV� "��3k����X��R�������:�J*Ug!�QW-���N:�	�a�f�>�����'��\�zD��,K��e�����!������Q��{ǽ|�#>R <�D��[�����{�`�l^��Q��ߎV"�YIC�T�[[�1�Ȩ_q��- ,.��*�c �)ґy�z+|�x��<ʺ��A<!����)�EU���Y-��b9�c-�1=Q��.Ό~m,�{r�*��C�t�b������D{� j~�j�j9��9!-�O��	�rD3jy�I�p�c�S�e�
�h�ǟL6Fi��1�jo+1W힝��5k�9��u��g �0��ȯBɺ(7�;�0��~������#u@�;Wk���:�Z� CG��^ x���ψ��5��[��r, 1p9 �WE�;�i��W����u�#:��wC	��o$TG��3�K����q&w��R�c.ڞZ�M�dk���٨%���l�����0��d�:v@����;�ľ��C�T��12�P�K�k���Hر8�i�/R�u�3D}_�Ηh�]����T�1�� �&��t2n�!oYK�+�3+ܟ��?=���ؽ���(��n�y9}fg1G�"�PA��\{��}hik�/���^\��U,@sb$��zޒfO�v�r7o��� {����@A�.�
��7�C%�Bp���y,z��O��]l�L ��Tm2��α]��Ј�����
J�� 8x1;��EW��OV�l!�)j��� pV�	�:��H�� 4�8XKbP��8#=Ɏ���W�܌�J. ���9m��s:_�>?����(���&�*%E� ��}/2�0R��>qY��I�<77�Y��N�Txi+����&�L�����׉O�D�h�e��._�����/��R�/��;�kW��r��&�6��ֵg�O=	^O,�L∎���f[�BA��v���
�wGBUe����CKJ'p��c_,^���)Z&���k:���ceD%}�>i��P?���o�_����9�Ϧ�	s���j�֖�f����5���bPg)��3=�,��6�=��������&F���w�ؑAL!�T��X��>)z>�&���W<��v�H�l�'^>�w̡�*�4��=w[�$<S��bp�����d��Eٹ�m	u�rth�u�R\�?�Cg������G>�+�n��qyɘ0��6;׷n5����/�p�3��BJa^Ɔ�>G+B\~4�X��o�ǔy���7�"���$un�}S|���?t�����%w�	�H�`?�wj�����C��*�:����R������ʕy�ى;��i�$�О0h�͓R͖�����aW[/�)�q�si����5����v�d��B�2,g0󎉯����bI^U7c�]�d��/����L7�M)S����4yO
4a�g�	B�^��3�Ecݚ�x�Ef�IaDҮ�S%����Dx��Op�ˏ�8N$5��Ι��ӊ��ҧ�u�r�]�x�「��,*�9����F�/�4��S�aY#)�$8Z
�2`ff���ʞ��C��H�"�ee��C�����%�1�.�Da?q{�@��u�,���ִz�I�D��&G[6G������C�� �M�O9B�q:��f(�HE,:����_M\���������=���sh�?b1I���F�n���oGam��Ŋ<H�kـ�%�����U,�(4!o�1"|p�l�}�cA�V�j\��F��fg��K���X�s"R��Sx I^$�
�T�ɂ�a��{]�����r��4��ř�AҐ9k��hή�����?jo{Q-�寙=���H�V����1�T���c�H�Q&[1'v�E�x��{�e�����v����Z���w�t� ��+'� MT�q��iQ9[�j�`�=%�����l&����4sn����,�>q�Ϫ;��:�h��GÇ���v�v��^L�o����Ժ�Eu��zq����U�B�q�$m743��P�,8v�C���Y���8�GRw�v��^t��,h)�Ug���&�]?	��%��b���ҠCw���fQ��-wy:�L6T�@֝u]s�`8�)�"%| ���J�'(�*h[�r+�e7	�p.��4½IT�躚�%��gSߑ:4���K��gX:���f�+
:o|!.�j��[($�I�2&{�Œ�#$飼�-����(��3;��ÔmH�A�45��t�/�_s�����^�:5{_�Z,8�~�h*j�(�iT�Y_��iÊOf��	�/����/��a���_�6�v83��R����$ij���2�$�{[X"`-���oh�!���c�n�*A��U�`H&LŁK;�G�Tw񥌒��C/4.O�'�S׈�d�����D#�>X���}��*�U�%���:>s,�/�É:�T�u`,�>p�k�Y�DF-.SƵ�d4���UMٷ��o�v#� >D�uk��u_پ�7=�Z�̶���C�0cA�,��WR�{Z	b�����B�v�� V�`R�=�p:��Ul2�F�,w^���V$�!�%wY���,���w+�^G�-��y���o1�b{)�D�r���Z�.F��p��bv^����6f�@d{_�jG~L�p"�HvZbrj�n���ɫ��������z�c��܇(+���)��XF�&/�ˡWca6��A����HE%�݁��M�#��gAgjY�1r͓IJ�L���)O8+[6[�l�N�"Gw�ѳ��
'�3�p�u`=�ڙB�EGg��k�G�)��r�P�[�2ۙ� �C��&�i�	��+W�b��`׾�w_9?:n�V�Dޮ�(>=�!�$r�}�^���\K?3G�A�Q3(�`�lhw1��t��W$�	����'��^�J�36��c��ѦN바ξ��s�Q�~��66��RNm�@(�xD�T|���%E��1�ȍw��`U�ҙ��M'�z�y��S� �E�w��u}��W%�q�����M5F������zL7��������
��u\d��@�I�9HA�V��t���G�rR��e�x��`�T��3o�������#Gk:\g�ny���ыe��9������PS!:�hȵ_"�`��ܤ*[�n}���4����MsG��Bs��ҡ��$K]z���F�`U��ւ�@)��1��A�9���T5�DL�U�4^Ȗ��Ka�#��4�ل�
�Ce�L|�cF<m�ɱZ�Fɹk��x\F�:x����,�rf�赙>c�o�O>燕-C�I?��x��-M���._�0ec���f�p_�Y��܁_�i����|�)\����ھ�wSy[��%}7).pgg�o��j"�	n����Z0<�Hл�ݚ��4��/��63G�k��~Ɨ��6�M7��rS0�i<�T6��ߵj���jQ�:��f/X�Իie���5��Gz�-�꒒�N��@�s7����mq��Ho�z����d�Z��v˪�C��5��a�b� ��3d[��h<���q͸���R�9}���D�%<~�+k�к�8$f�n]����F���'�^t�8�,�\>
c9��W���
�܂J�Ϲ4�{�� 쎯9��:]g�M����`���_�ĵ]B�u��}L��9�$M��!��d
���y0��O����~�b�=����G����q9f�vC�3�IgX�*�T=����:�e ��v���W�vk���]�*��Kں���������0%T��@�5�x���X
-HMk���-r�2�<���sͬ��lZ�r{ �=�H��!�t���f6��zAE�Y�T�ܕ��$�L^��IB��}H�'�ԡ�����g�7�{@���L��a&a�m��@�E����4���|��5���:�ݒI�B83�	���8�V�_'M�+��E�m�_^֙h���~�W�c����8���ܵC�/�R��'�
9b� B�k�L�7���<����y͝e+�g��{Y�i���hg��c~�<v���C�Z���B�tvb�ӡH
��uV訷��J����Ǧ������r��3[� �����S�q�A2V��9�]#sk���(+���&���0���1����Ac��S_j���[����������J�k9�2���f�V*$�Cs͙,��p���i�Lp�S���+	�B�H.�����Z�ub/Y������!��p�*����C��
��5�à{Ŷ�ޮ.�7��O��ZjO+��V��=<yZ(��d� �� 8a�^�}�d���)$E ����4���j�A2 ף/���W�⯞<��z�s3�DX��D���Qe#��s��3��y��C��i <��ȣ�Ip��X�g�H�H��ߚ�`�E�)�&:d�0=�sMYr��q������2��?��W��.��P���=�z�ZMS��v�S�1�m�m��э~�Ը�`˒�po���v�y��/�g��f�З�郡pufl�����h�-�=X�>Vk�����70�K�8�؞ ����x���`fM�
�L*��K��c�}�'�4��V�B^�;z�z�s�]X�'�����_Pɲ��@�r������4��z�aPT)I�Pk�ք�k�>����~у��#�x)0��j�.i���B��a7k(;aƺ���쟍�h�(�l�̆��D���
FM��*�s����S���ё�Ƭ��e�{��ϦEa���`Va!6�&���0���,qo�_Nr���% l���{��~��i1�i�O6��D8�
t=�g�ٛ2��nܡ��oR������%�?�W�0�_UnI��aG��
��h
�m?�q�RYYuKL��}\}������-�/��u�ŗ�46\O�B�u=s,��D	�@V��m=��a`�
q��f��dWJ�K3r`�m�4
�f
B�9�1�
_[ǿ]�G�u,`�`yL��c���/��.�Z�V�,�V6��l�.�	�7{�g>e".���C~tc�ו�g�:�M��HFT��
�h������	>kZ��h�|�X�6�(�HO^��ag���Ô�!�ٖ��y$C���y�����o��Μf���W�G�u4�|&�hTo�>	D��
=�zd� Dh'���T����3�?���Fmu��7���`/���0o�ó�@�+��+�"Fy��%��)����go�7�b]�j����0Iw��9p��A(��}f;�bҼ����$(L5��ʖ��:?��ҏ#������h,b��"�%�j���t��U��;*��	�cq�p�r��mc?��SKu��9o�����z��C�.,	�҃a��8�$��T��Q��*Ř���1�JӨ̐��m�=���T0��AW���H�����c����Lj�*k��;�`|�n�h��Y��?DW���o#��z7�	6bumu6�|,�N�4V۱ .���,�� �8Ek�=}���\�f�z����ug1��7,忑2Da�兤Zg�9���s܀(�`ye�.z��'�7t���Pdmm��ZCl$Ɛ��L�>�au.� �I�U���.~td�w��#bi]u}��b��ls�s��n!��jxNR�0۾37A��FP^�'�@#�=&���Vx��̮��%�*o�}�I|��d�3��%`���b%�n@5���R
��sɦ�j�5�y����;fW�§缟���sP۠Kk���1����*�k_Х3�W���y��Ű>��˔	��,r���/����J��ӷ8z^rnt`,6�튋�*TR�uKz,[�z���CKϴ<�8oE
a<_!�3�;����}��U�Ix�^����@�u1��˳��|��W��E�Gi��wJ*Z~�4h�����H�B���9]S�M��QsS��~v��/"�!D�k`iHL��'t�|[����8�
�t~H�qn��#GJ^(A�8Q>̆���$?DX�{a�w��5�c`B/][_G$�is�������a-�yG��+����� p�}}]n�	�fiW�Q�J�9v��Kjv��!l��r��땬��I�hs��%���$	#(���$��Υ���v�`�ن��TIB��~�[�g��x~�����B��I��a(���:�[�k����ނd�Gɤ��*d�yI���0c��=���.3s�|��j�,��L`�� �côہ�d����Bz�,��HX�ȠJ�~�t��7���c����tR4����%������:5�x����U����b�DF������vƢ��}׺�b�'
����L�Z�؞�]gcP1'��u�KC9�[{Q��ndv���|�i��l���tT�Xe:J�u!	1�����hC��K����W�ucWW*�(9��!@;W�uQ�4� ��j�����052��ܔ"?�ڰa�,(����҇7��f����(���L��E�>�ֶRB0xs0���ڇ���"���=���ѣ!Lx�?�����֚k��a�c��B��o�isa��2�`�5k�}ni��d*pE2�%�ĝ�/��k�J~�2k��x?+e�"�>�P֣�S��{J���y.�ً�\m?#�iD`�� �ï?{�Vȿ*�3+J��Y�4L�$ʝsq�Q����s�eX�!�4E�(OI��wV�^���4��+[�#
��R�o�����Z�-�/�{������-"�y�jL�����U���[\�Yt�)6����S�A��_�/��P���u���(�C�6�	^�����¦��݌џ�=b����ոb��k�e��*S�]�"�eN���a� :��ڳF&�xE�X��%��Y84���@��\ˋ��Z�e��1�y�7�W�6��zk��̰�S\�/���0b+�� �40fz=�z|b�v�Qh�
DIn�2��óU��(Y��p���+�5��z(#�J��'�^ƧFl-f��Y)�@�s�Y��Y�c�	P����D�UY<*6�v�{��	)�/\Ｄ}-�d�Nr��U����a)ŻNe/?��M�&#x�go��������N��8��,�No�c4�Mw����G�J�1H;��:��爩����[�YEw����V[�p��*T�x�1�+w���GTMF����~xs��=;��f�7�!���s�%�]�/�f���u<�
v]�h !81��5 �59�������ׅ�I��]R�H��2�w��D�
����?K����ч��ù~�o��B@� .�#͍�VO�(#�3P��ㆉ%�\����h���TT�R��̘�"0H��ca�؃���|����U1<Vm�O?��eH������}���F!SU� �Y��=̚9�\�l��3Oa�������;�W���#U���5��FdĖ~��+��R�����d����[\ܻ_��KeL?+6S�6ұl
��?�Z�J����5*��#�=���NU{3���gB>�����@�������Q!t5 ��%��8��H˵䨚+~��	!��n1b��	E0bo��U˦`�i�����߬��5��q���'~�T���	���7Už�YBd����� �V�m�`J�p'�6��rڻY&��i�:�M�V~��H�L�GI�Ʒ�������c�2ëQ0�������S��\��A�ٺ�O�LK���G��i�A�˽^q���$�"��t�����-AC!���ӈ�Ҹ���v;��T�n�{�mz@5pLE6*ؗ��v�eM��|��3�T�f_a��x��s���m3�)՛㤺U�L�r���w�5�ɦX�� ���:q���n�TË�\���)l��s��M"?�s8�ei��2j|��:����UU�m���q�@Vs%��-���ހ�KK��]�C��M
B+���I��'5��`t� a��oؓ�����Ѩ���O�tlH�X"�	�|v�m���P�h�=G�y�W_���t�ߍ�����1�)���7�>)������\N��c���6�1�,S�/��F��X/2.II5�=��ק˨����=�,�+N茑l�G��Vv���wqH-l�`��ِ��^�u�S�NhD��K��1*���#�	��W���I�n�N�siI�/�ItH�_A'0�g�]I	�;��j��&V��b��J��N�(\��0%����w�v'H���mh�y������3�.��߹#Cʸ1�A(������
\ې�m#�K�2�9�,w�,�B������ T�َTd������<*F�|}6�3��ȡV�����y��)��@�G����6G�0$a;����B��_!��^�i�Ϛ}*l�H����[��n\s*����Ƽ<&������Q1���{O�RI��|�Nt�D�3�ǧBu�t�ى��R��C�wI�2w��c�kz��
�$��ےr���r�������˜bM�>�!Oo���4!4]q/d҅��Q��ظ&�u��T+����!<� [�?��G�Q�W~��hT�$�Ѵd�ޟV7fa|���t�l>����ZP��á�wd��ㅿKb�02���"ڋ�OPu숀"G��E��%��Er��g����)���T�ŏ�\���ˀy�3�$�V��Ǫ����wa�-'�~1�-I�Wq����a��3w:�O+Ry�o�M&�!���J���"X����3���2V��vZ��V2�̼|�3�5�u�&��߄�-�-�A��l6t������[\q���Z,Eܺ70~i���>l跲�֓ˊ�������ьx�t�a�󟈼ȉo�z��`_�K��$�a) )�|�V��)�:�zt?WSOGs��Tz���0A�}����,m�	ѓ �z�c����&h�%v����J��[.�òs�_s�&���S���QS �P�1�([w.̂-W^�yV��+%�D�G�@y���$�E4CUǮ���Y��� ���w����˫e���z�Հ§�������~
�E���Y������(e��Ņ��{BWB�@ܣ�s�E�M��̒��h���G&Д�iY!��a\ψ�.�W�*�q.�%�=��MH؇��
�p�q��V���6��O�P������V���׾�F��/�����-��"��S������f���~���bʓ]�Wd�X<?v�Y�ώ�/c˵T-@����\�~n�ON�!��������m��so�eS�)�><M���W���4�y-m�$f�DK):.gD�(�$(R* ��s��R��S�x��)uʁ��1�x�	��Q�Oj���������a��k`��q&o$�y�5��Ĉ�U0�Y+ڪLu�1۪�߯mC]�u�Rx�a�bwD7�	U�"'_O@�@���l�+=���NoS�VD��f�-�q�j�!�Zq�a��֗��8o�͓i`���{1�YB�:x�%b���˒\�Wuϰ�'�X#���L�h��J�n�D��}0��$n
��9I>�*Ry?SY!75t	��2Y�����@H��Obue[�ǅum��1�Eu�����D���,�KߗJJT�{�RHM����^F~r��
�싾&��!�[`�#eY1���*��X� �f���X�'���艧�*g|+�R�����5�d�X��Y�J�"�&J�h��ۃ#�c�֏[���/������4}�[�BBMNf�=���/\���l\d#>��kE'�J����%ժ���X��}��A���?[����Jh;n����~1=ZZHw(��"\j��'[d���j��+Z������jo+_ڟSv�����Rш�;�Ͱ� ?�'0�-�'����=�qAÕL� �����GBZ��8�S�7�����$�V��пN�7��H����Шm�O�Q:�c�����<������+�hz��̉Ԭ�C�)Մ1c����	�����\�x���9��U68Zb�9o���}G.��+0�*���i(���z~]w�)��(��S���$TD���5�ӑ8_��^b+�p_?���qM��k��V	���|ܳ�	ڕ��ҫ.�{�Ǘȧ��U䱇�����Ȕ�p;�)�1������񣼑��/KMӧq��� ��)�}yfr��g��!g��-0
&Z7K����3���7��y��S<]of��Q����f�-�,z��U%I�~�<2��"�	q�So���a��iB=O���F4ή<����������/���2����o���֮��/ߒc������Ш� ;"������p|2��@��p�P�����y`��\!N��[�VQ3/�`��tm�3z�LH���������ݛi-.�F��ڳ�2Ϟ�vn	��ݑ���^pB��cre5��m`(��6���A⾳)-����K m��@PՎ�5k���(���� ��b��\Ԫ���D�WR�'�J�08�B�y �j"�`�/=��~{����#�>���x�ś?I�@�%ԓ���)�����y�?���<����G�k	L�wE-�G�F���[�xh4��|%����U�;�z�ȼ[A�\�
���V��T���%�6CU_5"�Ĳ��'�G��^���8}l�|�_g�_2��a3o�D=����qq"wToz5W��H":���t�����wF������8��Ú��ol�09�g��IG��R��HѲ��܁-��;\n	��;B�όR�x�=��؇�*o,��8c��+e�K�2�?ѵE�0I�!�8�n̑`��Ԟws=ך��5�* �,Akg���s�����T�����[t'(��~m���+8��/���^,ߣ�Ehp����}C�WftNɊ�6�v.�������F��N����X`p��P�G;�O���w;��JCټ�E��P�Lkq`�xH�a��N��*U����w�Ū/Jbue:w���G\'�JHsh�=\�^\{��e��EvyNG�+a{��n1k�J�+"�Ƌ���y��T�������)���]͢�m�>���ڿ�k���'Т�&�Uv��y�ʌ�S
z|8��ј9�<��������DʹAHt��Tx�ɢg��#EL�k�`��e���Q1rn��Z��}��_�Yk'���$.ۊt!���*)���+:����"�w��(�1K�M���~z��niʣ���x[�<���]M�3��&�@L���:��>�v�A}��YHju��J|��F���� ��h44���5zr]-qW��@�����wY:i�ϤY�q(�R]i�H��n�Q��J/C ��.�f�$��a��dѣ )
F���4M��\u�Gѩ{�]�����'��1�xa��E�@>ZH/��.�q�Ɵz��^_��Q#�,''�V�313w�#Ic���q���s�xԮ�F�8����G�ᑞU�-��f�2d�y ��^M]���6I���Aԋ��Fg�Q/��b9����8 �'�OK��C�ć�H����m������
��d�d�iw�A���#�n�1�pO���M�Z�\�\ޯd�$��[V�t]w�&�B��.��N0<36���E�"�����\�p`{�~J�C�b�&���=�<_��1�V��	Wǰ@@q4@�4@m�h�z@\�K&�,䤅�>׉����XJ����5�I��,�CH:�;�st�"��q�� �5����䓺�0;HRm7����u�4ol:���J�W�ר���.kJ�f[�ܨ�
ܹo� !�	v����j�o��fM�d;�d��ಊ^�-+S o�E�����a���P���An�0��~7M�Ӣ���	i�=._��MG/�T��o&�\��U��"�g���e���*{�X�p�9.�"�^�A�}:�c�7�Y[��`�t]�d�b�-�k��)���fn2�vJ��^A��jq����?�k� !L�!�==�4Z�;�����j��[l^_���©��v����Ի�������ԃE��|����A���I�k����͸��L�ul���ܟ�1��p�U}�y	���O�~��� ���m,"��Mx#�PH@�힤�)�+;"�ռ�;M\Y���4��bl�
:�Wdw��B����xw��i��"@_�$B�������W%
��AXc�a��&=#e�ri��ڲ(j�4u+�r����gql֐�\�X�m6Peƶ �12���h�i0~���N��J4�����P��$3���m�b5#h]�\j�B0v�v�YMD��V2�ғ���
�'�:�^��8�9�U4�g-��
y��U�Y��	������.zO�^���q��A���67C��1%�0:[�E"M+�Z��k1=-!�~yg�L%,�����S�z2_ʠ:0��z��Ac�;�PY�Xp���J,�s}��PXG�<��E�Ճ~��!�.���iSC(<�t}��[2zv#�,oL�r���v_��B����#|�D���di>�+s�� �8C���䳋_��'���{*d��5�P0q�]#O���߸pv������0ؽDY���p=Ww�"b�b#,,(�1�a1�?�{�;���$�n�C��F���Y�������'��Z���B�;~�wJ'�9F̑wL2�;b�a�Q���0f��BE_&G]���g�.��^%�ʍ��\��/��bk�n�����?����@�ً��8����[) Tn:�Q�͕Q�ɮ����T0�ʬ �*E�Z��d��ӈ���}"�v���\�g�B��uZ	{��QU²y";N�E������h�c�7� e�M��ci���M�2P)�vu�c�7��ވl���y��á��xfh�v7��Hz����0��х	<�m��#��P�,������`�������.M���(�>e䊬����[��*\�1�ns*u���"��Q����[C@�Dti�qM���~���H�7�؟녯A��n�]vc<�,B�.h��y(��#�b��5Ch�Ŷ���0E��}�ҜBA\sK�P�iJ�L��D��W���[kp�$���