��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�۞����h��wdIv��ta���HO��CF��8�wL��-�CY�{f�VM�*7KKo2�Bۥ�rF}�+M\���b��򽉫������_Z!sC�"T�Z>�����b1���f�9f�^щ�X�lD�� �	1��:u�u�R���Q�9�Bz=�Tj:��U�+���G���:���:ն�f.��L��2�����i&��j�C+7!@�P3iѪS�Vrt�fA��>M=���>c���s���`�X4�Ñ:,�90J~&`p�N��A��Xg3�8$�Rn���nf��o�w��&3���� �1��� 	c�v���:��k�D�W���~<=ʄr�S�De�6�q��^�]~�㙲�Q�饲�0���(f�ࠅ��Zb���.B��Y긒�->`�j!����1*�i�p/�_fB}�A}�83��V�m �ҭ���ֻr/���*Ȇ1Dº�	�=��*�?N~�9��<_f����>$����TsRCm^ա�^6�V�r��y�Yej��1&nbUT5�-g��xIΚ�\X��*�i(eV��d���~ ��~�1�A1\�$�s�������3I��f+�����z����+���8���!�Nv|�|�be�Ww#êN�
��P7�7f��,K��~+	N�b4�x�����X�6�V�Q�p����x�H��V>��n��,nn��{�=���T5�{��@��.I���.�51�Е@���8���X�ś��HȲL��v1�tX��9m��Jӛ���#-٩m~��ǒ�����?�����n�]�[�L���nrG9~Ǚ��m	X6j�W��d6�QQm�-lջ���"��+�ln⠠�?����]��F~��
������+v.0ɘ&Qm�C@��$�k��Y��m.D��.g��(L���w�$b�Q�aCJ7��3?�5;��3�@ڍ�ɾ�S r�V�W#h��?C3y�W6[%�:��L}w�0ې
U:F���/�Xd��#r��hLǕ��]u4�k���
��=���D�4n������6��COR��A�⺤�ߌh�`@�ݳ�~z��[������M&�Eg_��p�h��_�+M ��FW�9�:�����t�N�����T<��p��OJ���ۣ�~��ߐ�u���"uBv��F7y�\ضW��>nƒ���Gp�T�C�/� ��?b�����
Y� 5_3�<=-)^ή� ����@;�xȚ m��Ny�<`���U�0��S�:3��V�fo�m�|�	i%Y��Zd��b%DZ�^�M=z���ڀN���:�,o3�Z�}��ދ%��� �Y���ZPOɃԠ ��O�	����ntR���J3�GAJ����jZ���E�����<�Xי�5.qо�0�ѵ
S�R�?[��G��Of�R18h8X����a��Y: �G��ĸF0E�Ř�E�BX^_L;���] �j,L��,���J?�{�3K$��4��v>�y̟��󬕭�&�g#𰨀�E��K9D�*fۏ��M#��5[٘n�V��#�C��=\>�b���ĉ��eg$p<�����P`rQ�kOX������ZjE�K���j���_G$�ɡ�ʅޢ�|%S*��]t$����aJ��_����+�_S���˯��7�P���3r���r�Ep��7<.���Ӆ�RK6��Q$n�G�tM�(чڿ��AtXn��j�쉎�Gva�	��c!Ld1y��|yS�J@��E`�Q�0㇌
�������$J���l(�N�@���ʴx�~ʓ��,
9��e�J�m�����������b4�nƫw�m�-���|�F����Pl��E����!�|�Gے�ʉ��f�����ff��^�I�nfՃ�]��g��c��� ��$��}d�F7�.)y�x`Zf�}��g�2:O c��X;��m��0Ӽ}�Q:A������HN�2~��)Cd;�����2
ʱ��`�~���l#�!���u[`U[���1�!Os�dL��1���2?=��Ņ?4�(����xr�����+gVv}���8B�'8��W�{����#NTN�AX�r���2,��8�C��lQ%63��:G��vp���*�$:`Y.(g��`Eox:����^����%��;m�6Q�>�*"��ʳ˹���K��o�+Of�p/��>������O�����=�pifαU�FZ̚����f65� ��z�s=�((�s$���J�_�C�,���,��ޫ�2Ɋj鿭� `*QZ*���#\�r>���k]��F�d��cF�L�Gի�a�(m^�~�(5ŋS����8$�=��~5!\�-�v��� �C���l!F��E�W}p�����aK���-G�
�3x�mW������~����lQ�C}S��3�t�mW���f�i(nC@8�bE]�"�|��aW
&�aC�N��?Y�%D��:�O�=�ܒ�0;/g��h����`C!�d'�X��lK�����teSa&�8����~J�.D��J�Pםi	�����Fwh9���̰�َC���_w7�2�C�c�='��o$�j�����&(�	$o8XPV�=�ĺ�x �ڵ�FA�5������X�|�l��v���|�b"�J�͑��������4m������ݏ�'�~9�8�߭0�bS3:�� ��m��~'��pđNV�0hB���"5
�n1�,��qs��