��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��NV�3j��PS[�_p�8_\|d�w��JZr�<�Bql�����!*'8��K����Bߏ�ύwvcc���%$d@N"���/.�����ib�Lˉ#�N�:��|b&��)0}�@���`|Fۯ�n~H�|��`/>:���e��se/ớa��[��=��RFb��n���*���9fH&-�I���s�]�lmz�rz���O0�%��q�q3�Њt�;-�ϊfk5�1�1������@��tF;a�Ծy��!D?���H�zҫFw�7%tHXs+��z����fX��R��V�y(������$|V����\�2��O�w�5���T����&1���9n�1m��A��k�}$���V�(@�1c�ƈ52�b�ف(J3�)�|\��/�Y-u~Ϭ�h4��Af�n��S�leQ-��&���5$��S�:er uӀ�\�U�q="�m6(��5���Z%�J��c���zo�{j@��=@��)�Y�?&��}�~^ ~z�m�ndi���+R�۾�D�1FIg]��<�O��ua��A`3�]s���u]���%sF�px�w�ʕ^���0��ٗ�@�� �Sf_G^Yk{�*�����k3rzs��ok9\�>�>�@Ze*R/�vI?_�:0�w��g5���)�P3��1������,k2�A�[|����-�"+�@�/��J�I�����$Ҟ��I�*A��#�g�k,鿏�?U�L����Bbc�а{<��|b/$�'欥�x���nĴɐa��#�5�nW!��L �H1��QV��]����Hy_/#��8��K�bl�޼ˀA&�܇�opwW��0T�4������l���+DM%9�m��}"ݎ����-�}����1�5C����b�B�{��8C�]z��ͣ�i��7~��������L�^��O��-N�6�Ǝj�R�@��ހЏҟ�o����}����")6�3��e���z#v��{Z��g^�Mo�|y�³)�-!mfI ��q��u���&���?uW���&ǉ�yF��."inb�	� &�Cf���ر���܋�[����-�T�x*�֫�p( �(l�Ԟ�n�U��^�7ZK���do=�>�!�	-��GT�	�N`���f�Q�'��;��l6�:q����F���H*��+�]2����nI릡S
k�6%{y�h�Was�GLɥlWr1�Y�34Ԡ�����a�����2����h �i�8/}C�֎e]����K���<��>�h�)J� LR��1B�ҩ���`�^�?���Bd92	$'�w�D.�j�tr��ז�}��;�����/R�ɣݎ1�zY�=�@�2;�	���i����U/�v*�]�.{�[�=�n�J[Uc7hZ�;�;+V����@�Y�	a~ �O��#��+�N�xyҰ����n�f�uB6���]M���WZ����v+q����_�,�����R���FD��V��0�%�>��Q�"�O�,��S�����	(�vc*F��'��A�7�J�М����x5;jYn����~�}�*��g�U��i��&sUq��@���N�kv���D"E��P�l�n:S+����a�	TX�J�\�}(v��P/@�O�Bq���W|~�cX� c��H��앲�������8��sR��y������'m�`�֖��M�{���A���`/9C���Z �25x��%���%QO�v�h�<z=*\y�cۊ4�J�e5Ĭ�������-�3b" �s'~❀s9i��P]b��=��Ρ�f��]�Pa��QV�M���ff5j���}-����8�����'D_b2��pd�gP�㿠�bq��8eD�*�j����M��7b�\8�� nw3-���2<8$���3�DN)No��Z�H�\�P��,Uu/+.�ޫ�΃����02������%wQ����NHV��U��8("S�� ���\�`<�9O�7�*�E\��)�BV��N��򶰽�E��X��4�M��ڎ-�nȤ|/������ql�b��6����,:����˘(�|�2�y:	�����|��"�S�VB�_���./ltpaC �T��d��8�(��
���g +�^
/F�`Aj:��
l/PM�A�&vP�<��t"��}���0,�}�6͔�a�9�|�ڞ�9e�9o8�Cf�Mp��� La`�Y�sPz�OwzO���e:j�i;�(��3߾ ��?��Hk-7⏁����;@���l50�|}{�~�.��~x
�1q�u-���^��]��~��Nl��a �Z#�q�5�\��`��1����q0$z�{�W9���:�j����D�{�dH���k������A�0mX?��� v�&����������.#t W�{�@�0WX���N�����6�ō��D�;���6ɶ
����y�J�޾?�gq�/�<W*�;tlĖ�(ET@I���{�|4����!�9��۽���r(��0�TF�=l��<_�"(3�����K���"*g>}���4W����o��;�E�]!*<u�|A�'����!�ձ~�^!���H>�|���|��>ߙ�}����-�R9�U��.	�cNM�l�p�#쐖"؝V��L�h�sb�r��2��#�3�=�4�ΐ�l�%VjL���(�Z\����5�"���n� n�Ƌ{>Ħ)�#�2��+�@��N�������TT������
m+ 	ot(]C�Mw���ҽ4�ڀ��挄~ޓ	�+�:f:G�F���;�Ȏ�Q���k�V����YO�s��@�z���4�&�FT��}�h�ݡ��N�Z�f��7���#R�����Pn�,u��%�7(���&+���ۤ�Q�LT#\� ��B�+�~�<�&�YrX��a�ԫ��H#ua0 �20H��b��fFi�$���k(L`��->��"���}�S�!�VI�<*dp��w�U-G�wxv���3�	����q�-e&�s��?�ڒ��a~��n�^�g&^�;��k�����lz���|��z�l6Z�@�d������=�����#��˱rΪl��OF���2ɦn	hgno}���� ��AM_�$ӱ;���b!פi��2����tUwpg�d����]4��2?�Q�0.]�ͻ��'�C�+/{#���?�4l��>��bI�^oȃE�[2�����N������6ݵ/��P���|�Ǯ�����;U����iD�O��,+��b�R��%���奺�?����,"� }_��Ȭ+�X�C�C}��~��pn��@��|�)��vNБ���h߱��<��1���C�����ꕼ�Ȅ��!gԙ�mA`Ѐ�\M<�����&0$��I�8*�OD�Bᔷ\o:a����	F���a>4�>��l���ً�呫�iV�wb�;�K�ZCw��X\�{f�28+��є�`p�ו�]u����!�6(_�[����i���l՟�����&�߿��) jL�W뽙�����PatS���;��cf��ᒲv?�$�C����B]��Kw����o32��+M��/�6���G�� �GH�T������R�G������lQ�;r��{�����	hZ�d��9��gb�AMt�D��h�_�Ȏ��C�䩲�t=E2��E�i�@a��Ķx��6��s�T]t�g�r�;�%��4�ڝ��m.���J���y`LSWc���L�^A�yPt�zbx�֋����k3`- ���1�]T?���3�X���<�M<S�����0�A��f���m��$U#�路��߮͐9�=]a? ����	��V����]zkK��!kàv5>R����j�M��)�ȏ`EB�H�e;A�J�_����d����UI��d�J��n�7I�u�S]t^O;J�kr��:q(gs��������߭x��#P��;�Έb��`�5�n;������N�Z/�V6�j&���y�W�胝q(�3�����A�ط�T� mC�i��|6�Y�k��O�K�S���a���<�z�JA
�皺h�ݐ�/*{S�cW0$�<�Qd-�c�Ibq:�غ�V��x #�\���`s��x�Jb]�Xr"��-�g\|D�鮵) �������so&}�h���~����ݒH0���s9��۰�y�ŀt�<�,OpYs�_��e��C j^o]^�6k�>QS�i{"N/�ߪ��˯*Ւ�w�OfA���)V��|�%}U҂�?Q��ە��a$�4�?�-�}7��oషAry�ծ��"�0^�`l�W���`q��
�Y���*n\�����b�ٲ�5�o_k*W�VJ����2T$��T�ĩsҞh����1&�jQ�9�t�Ot����1��g��y?ڂ�-���̊T�d��5���ߋG�u���gr�����0aK}��@[`��CCQ�m@�����n$b��ut��a�H$�<w?8w,�!w�$<��4������/��bt������:��,m
�<�y*�0�9�e���部�c�6�O��|>J���Ǖ�A�����o{�G\����{�#HK!�_1p���G����%����/��y�
Ň �8���e�M#Q�1ϓi�������;e����I�N���~s��R� J��ԛ�yT&�.��Ӗ��!R�y�ޝX�c;H�-;vi�6���A����_cE!D��w}�ۥN�d?����(�i�6�1��#�! h��1��n�&^s[<��,m����}[������qd�s��SƐ:�� �Jp�aof����\j�'���k�ު9���-�_�����d�s��#�d�V�'j�\�ւoȔ:�fRF���;�lV\gmJ�5���l�W3%�v��4M.W�{��0�������G S����(m΄l�B����@p}��%c\�L�@$������0�(@�wꍤ��y��1���z;��~'��t�D�b�w�bvFD��`�dO�t�n�B����n�S�o.L��ۮr��e�b��a{~�T�ѷ�e����r�a2��+Q�\Z_(wz��U
�F�f�����������`���;��%�O��z�M��=ba�Rx�a���AзͲ�.j�=B&���z̻<Jg��p5h��/S�`�O�6��K_M�4~�F��7Ub�C��P"�j��&u[x�L@f���n�A�Q�ZۛG%p���0a�P �Mk�Ѡn��20�VL-�'�����V� ��.��]6��'ŌH�Q�3tMw*��_�����Il�7K�	��F,L;�a�
��խ��M] ��-1푱�m����.�ڒR�)V�sw��0i *x����!z�ĊK��$�q�X}���_C�?kd2Yns��b;�����7���6!(���콻�MQ-�Ǚ�I��c�eV��%&���N_"�y��ɴ̢�{��CrD�{��ݔ3�vbOX�_k��V��9���|�*ݗ��k��}�ڱ`���aC��<6� 0�;�_I�Q��S��2��Y�F�\	��{[�O��X&F�	���Xٺ;��-�ǭ���`����\^�6	�)��D��~[��D�Rn�v���-�}�|z5����߄���˭����D_�#�ȣ�s�c)�����v�Jb�Bg�-�s&�b|E5�!I��4cQ�95�~��ΗtF�l�V.��<$��:M;^' Փ�#]	���'�!�Ӷ�Y��9�o��
����
x���ꁶ�E�c��T����U�����7h,@��G\)�ޞ����o�Ӯ�6�7�;��Mt N�̔��[�X޼�o�rUw��S+WH3u�{����/�);97�?5�z���%����GQ�o&���!H9�A�EN��
��)?�xv�=���E����W��ϯ���%�r��k��yZ���M��K^�J�����|ue����TC�b�����s�i�$�n��U��/D[�9��w�It!V�Md�e�|LN���t M2빵6j��*�Z�7�]�N8�e{.p�j���[K��U)�(���=��|(��q�	1�w�~�[Tk8%[��)���f�#mͱ p���Jc=����%���N�ݛ�%=}�w�����՟�x��c�$o/[q��^q5������x��T=ws;�-��U�3#`��z�k,6q0��l~�,�.���h�k�����}�{�4�1�$_�)O�Vޮ�n�M~o�dy4,z�#M�Fۂ�pq�y�[�����3 p�'.t>�.�Ԇ�b�U`T-a� �~���U���i 0����� C����C���6y'9)g��׭�;�U�9MP,�u�I~�Y��i&@��� ,`�����m��H�W�=�0g��O�m�fL�_ߊ0���H�SClp�G��
���#�־�:A�e��[ 	
�>XF�)M',�q)G��������y���R%4i�Ss�3K�}[�4��O���K7��1�����ץ�-*�p���ijL�BH��Ʋ����df&��Ȳy��Ka�!��O����|䖾��4��\Lfdv�Y����]V��<!y�}7'W,+^���)o���C���3�e�|�#,�i����q�`Y�1�g˗�bd��Vt��yr��nťQ�	a�c��S3�@d��1�A���ɣ�T�'XoҊ�]��H��P�{ ����W� ��ި��B=�P9���f�x�`D�n��!���1N5p�gѹ	3�-8�s.ͶP�og�A4������ZS�;VB���G��۬4��D���A�E�D��ꃿz�qu�?�%6���D�X�pd�˷VB����Gű����a�q1A���b��#��JXX�i�,"�pےکt)��,|�U�\��2W� �W��oO�L�@���Ƭ}���`�Rd�[�SX����{�H�a�8I�2}��GƤZ~����}m�������3Fg���Kנ-���v��N�
<���GQ��a�p��0g�3ajO�WgYS���8�HW[W�k$s|��;�WuG:�~a߸�r���+��^}V>.yĕ�w�G�WW�W���ؚ"v��s0]qt�(�xYQ���'}��l8��F�8���(��|�B)!�9x^GD�Z�0��D���$rd�gy$t�Ҡк�ꖤ�n۾�<%��[���2�T����^#ka�e89�G�K[�PK2uI�R2-Dw�㒌i��.�.-�1��z�� �����~��0�|D��_T|��,��VW�'����@V����F��V��(�I|��(0��5T�{��AL������S#��ҷ.݅����ȌR���;��������bFxZ�V�c<fvhV�{>��8K�bdmT��VH�$��f	������bu��c"����j�b7�|[C�+~[kQ�|�n!�>��#z6���T�n���N�&���n8�2�۶(�Sn"����{<�Zz�)H��2u���0Af��}�{�&I�/�mB��=\ ��(���12�cԜ]c�vE�a7���i��I�7����3d9j�K�R�k���}�H�<�,��{�Ƿ`^��0K*q��K�f	��c���H��b"D�,f�X	���I�;K�ڌw�؍�{�&�r!Qø��"]є�,u�^���b���@�@iB�E"�J���x�.5��;(��b@-�YP����G{H��H���Obg~��$`ɂ��Y�W�8�m��&*���>���o�V`�zV�;�~���N�P����"&������B�oY�gq����!�)��.GG�<oK]4'
�νR�;�~�Ǧ�':Ę��o�6��de�*�{:��7\�<�#u:-?�)���͵W�0#����}\��.�Y��H?ڍ����fI��Y|��8��e����z�'�{ X����<ib����{�Ef�]&�V"��-O����p��,
�Q_����k�=-\Q�Fp�pa������o�#�q���������Q`�`����f���E�G(hB.d��v
m*�ȲvG���T�W��9��G��Z���o{s�Ʋ�6c��\�������r��ƥ�Ŏ��n�V�3�9H�]Cn�1sդ�VH�qS��W�� ���#=$%��*F��,~�G�������´�v��
 ��w~�h�$�� ��>#�1��9f45ث�����0<l}M��1h��\�6�\�Tr�z����{��wbٰ�Isr�N��Z��ɐt""�QǠ}tSM�	'jvq ��[u �/��Zq+�4�;b�Qx��@�r'O.�6M�[U˞��-�x�C~s�u������s-���`�S�q����.��/GBKs��U��ܸ�����1��C�B�d�"�K�FY�a����ݘ
o��V���8 �2V<��>�T�2F���X7��[�ދa˗��S5Ѷ�~X�x�at4[<NS�=m�M�w�(B��âoHo-�\�Ɓ��}i^jZ_�E��}3��@&YaJn:�V>ɚ�Q���sd��Cر�iG��W��DBaC���~�}�V&��X�n��fCS��5w��;�rz���9C���Y-��+�\�0k1�eK*$�F>!H��TI�K[�q:/1F�����r+��]}��W}�SYs&���Z�ْ7x=���F�ۊ���}��F���/8W1�1�}�Z�2��KV��N�2\��3��wHсr��A7�sΛ����AS�3�˂�m��W�8��^Zm�t��b�	f���ؘ��o�mm�A+�̚��r ҂�[/�,X��3�oH3~����D��*Uw�.\�b�2�����䱋���n�+�\c�b�S�x��;L4�s����������~�/T��SQ�$/I�$~�����Л��*� #���3kj,�����h��-��WEb��-���w�����"�$壩���o�J�c�^�p����X.t����';��� ۳�b�E���sP���!%������p�j����~	�$kq(��SN�e^�e�;69d���Y�8l�ƢDY(g�L�QX��YW59�ߖ����+�2�2���#��ۗ- Wh{�$)����Vn
*�ȅ�r�}#�8(ns��
��m�Z��`&F7�:���@XD�������n+��ahr��������s~[+�Ӗ8��t��˂�1���'c�7�T�����a���<1�<%>��Î�^����Y%wR�Iͨ�9��y���s[�&LY�kG��ͼ��QE񁊐���7MaiTt�H[�G�o#�{�1�̲�x�?���(�Ϡ���E!��a��ٞ�%=�r�ݺ0��1�."&�Wྈr.����I#�u�e ���5$��P���~|u{���ؤm[��/��^��M���Y7���&)��s�hx��?����7o���-D�����Z�:߫��oV�סxy�K%���s�N��ƽԫK�%+�%�5)�� �a�#��
�����׭h�s֖�B��&���kE�����DH�P�<�o[t�J���K�0oP�5�91����%���=�;��a�.�ھ�sG~�&Z�,��ɱV���0� �!���;�o��`̎��-�0?{��`���|�����$@Z�:3�]A�����[�I`��*���a�Ӊd��Rn�u������l$�Z|��Z��?�Y��ѻ
pb��ɛᚔ�V����wd���������L��b��������tH�c#hH�T�<�,_`���e����Bx3x�G�S��U����E���oH|�h��FܷzǸ�P�щ���}yeGO`vf��&ǑHO���@
� �Z�p����e[05��a��5f��Z�IL���,R����0k�����3k#mIk��&Q��+�𰄢���� f�׋��{lq�Mը�,���,���3�'�/����-:I�waH7Q!$��$�9���v����]�%��'g��s#t�?%�=�a�a��o�1�w&���j�,�lҮ��c̫�@�U���aP�����5�
�\֗�"R�����sEƆ�WJ>]��h��.�L������i��s'q��*6 ���S�e�1i�qZDB=�G*����s�����z��2ܵ�'�3c��枥� eT�h|�7��O�2��&t�FI�G���XH�Ֆ����}"Ϲ�l�rB�� i )pR���(I�/-&}.`�vT����6���|y�CP��d4�Ui���Alg�½.+�����F��Ά����ؗG3E!�yEOz��-I4Ġ�;0��_���Z��^ж4S��a<���4z�v;yݰF��x4���5a|]�A�xw�m���*�4Z�Zl��"ǀ�59�;��7մv.)�{��m]m��-�a��p�Q!���^|�:ԃ������{J�}����Ew��F��H�=���������FW�e� Vݺz�1k�_�~6�kMݺ�0��.�:A��=1�[7�2@�����GUceҚrd�H<�i�3���0m�6 ��ȬJ�I����(�c8J�#0��3]��,r��*�;{ߴ�ف�xݺkTl��1���E�f�~�I��b���J�J��JI /�?�����A�N��#�&RM�^���]*G��7F�N�\��F����[Ѐ�B|ˣ��?�Sŋ5������H�I��8�����L�?0�z[ķ|M��	���b��nn���㭕x�D���Ζa|�U�|�T�9��u$q�m�p�[�Q~}��g ��e�g�<���F{zU�)*�y�Kl���S�$*��<qh=�8�G�5i&T��=_e��/�#cX�P����&��p�������P�A�ָ��4�u����i=Q���D�Pb��.��Q|7�ϼ�7?{5�ҁ����Y��`3$�l�����hf�L���h�ܣ	B7[569L����7�2���?�/���[�8n/�{�*~�����z�������7�l���IO����$�/�*O�n�._�w� 1
hP� �M���:J��U	��o^���$����5�_�����?׫�6w�Um��;u���)>���o�!�8�e�#�Ȅ/�X4Fp��~�����2�)�좯��L��	-�WcĹ{ ZӶ2�$��%/��曃���ZOL� ��f O=�!��s� Ps�$c��4�w��q$ީ�Fb��X����|�w7d&~_7�sy���/�@/�������<S3�p�Ҵ���$G��@[�����s %DJ!Sz�9�%� `�=�˃vHN��Ư�q����-�WI3��pz���74�~fVS��m|���؉�	n��nt?�>HҲYm CXMC���+�~�k0�,�Hd��.1��i>�0�u����ҌU�6��ˑp���Wȡ�+� �1b�-�|��N��4�H>��@������`�e�й0��TY�8J�S����T��ԏ���������!YC�*k!�י��D�� G�o@�
ݢ�^�g�/k�Qq"<&��.�V���Z�j��Z��H�%�����<�t-H#P� [%�|�Xn��˓�UL��k�+8❊��Z��u��Y����F:dz��Z���9�9��<p�z��ʉ�C?�f�F!�(B�����l7��=Z�q������|V�)M���e�#8��Z��~#<��ΓJ��V�")�~�$���cޞ�;����]u\dk��n���6��Stip��S.�.����T�\jl�N�F�p*Ļ���8B/<���w��Տ�_�㤋�)���3�*���x��l�e̍˔D{+���<DB���R�-EnՆ�#2�C����U���s�jI��-/�e���J��.�Q-ʗ?�qb��c���s�ceD�9�B��h�F�"09�Ic`�S��/�0P�S�D��?��4ϩR�:j��|�Ϡ'�`o<����d�
= /vg3�_V9���U��|5�b��|�� H�#��|�p��E�7��\Cx��d�n����� �ӣ�89�(�lީ
���ZYݐq�P���k	@#������8�.�������'~Oj%��� ��}z�i��t7���I��!$�\�N�(X^��w�/�l1��I�o@l�R�}ĕ53'���ih�WN�9�|��
Z��F���{b:��+ӱ����5
k~I���zۺ~�c��-�ϗ��˸�p�LF=�P�'�>-��͟R�ƒ5:<��76�	\�0���9NaLx�C�=`E��j���"��ԩ���@\fM����ޚ�LBM0[";`_\&)��#%̟/�*��<>\�D��G�����eU2��ݯ�G+L���bo�Q�M�kYe�󴤢o�g�����Mt0��rY��	|�sӿ����=4�a+��bT�� "�Mn�$�"R"�Z����<�#���o���X�+�O���4�l��Q7�%��g�'�ݼN�F���H"z@0���X�+$�C�|����C�I��R��掭h0
Qٻ� ��{b�v /A�.�Y����0�0�r���|�og��yj�J�ٕ���^��Ax�F���Ͱ6�s�m-Z�/"�A�� ��L2�N���J�~Ytq;G�7N�u]�͏��.��zƥ�BN�E�G��|_�vc�++Tjo�	�;��h
�5hިE�[g�:�C ,���o��K �sP�b�)F٘/|z��&�y7jX�M�L	��`���H�r�l���t����r�zIs�Yt��z�-��:��쩣a��-��*J�CK2�FYM���'�������6"�*�f/]���	���E������F`ŀn�+W=U�������6��!�d��cB�#l��Ďkc��C~#[��NĆ�����6Q��i�Y��,����X��m�s�Vu��]�Ī�`��S#��XD�˵�wL��)4�����ى�� ��g)<`S�.#�Q�A��֠�|�|{���;N����Wt5O)/ߝI�+u��Qň���STK��=��lq���ˎ�(K2;M$B����ѯ�`+�DBx���	YЩ�P�k*�|�@1��?b��mM:�-�3`i7>Ǖ��f0G0Iޡ_�@�{��}��*�G����{�1��5Ԕ���fV�:�>Р$�n�W�
_�t�M��2]	
�~+����'�P1����9�����z
�bd�&�2�ң�R�\�&�s= "r
�����^# �/���i�����L}L8����}����յ��&�\���q�(y�ҧS�q� ��=��::z.U�V��Fb�=t�Q��Q)\>��x<|8���OajN����x8����y�'|1Ľ-���)X�%Jq�5jҼ���Bt�PC�Q~�x��O���@����kYf��*��8U�����7	�aV�f�cn�ģK�ى�z��Z�����P���d�Gv��!���{Cy(��g�e���y�����{ �"+��f�?���ťǸ���~؉x|�3:�{�5��,��9�Ch��E��C�W��K�{��c���x��5����i�J�Z�3�KE�NYve�GͿ��t��\{��'(����ܗ�m'��r�_4����1D��9�,��Ձ�G�)
�[^�gB;���M�q����EB<ؓi}���*���}��(Pf�QO(rᐩ.�D��1����.�""@na�1f����~Y �]�� ]�Q���t:��XCu۽�u�ܤC�����`pX����#Z��W���gP�����|����z�S��K��I����&Y-�c^$B���a2�1hj��<;�#`�	�6c����~���A�K�4�͑g�"�����!/����f	L�S�J�Ύ�CwLE7����H3��S��w�Y����D�����H*u�5��v}?5~��eBA*lWX�-&mQh���l\uFh��m�{��тl6s�N���iqA;��R���1ȤG���I����Y�����L��6�b�3"���lf$�O��jy�?���h_�5��5c�u��Z@�}��A9�0bDۄ0��a���`�QU>��-߯l�h��䂝�bB�=y5�1h a��*�+C�9�a)�2����WU�X���{5pԘ&z~�Y����W�C/�.�������V9|���XхM,��x@��	��_Lb'KBvK҈�����C.��ʛIL
g_��m7d�`�ɑ>,���w�+lێ	F�n
����乼��]}���d���|����o��'�[��K��_"��nW��m��S8�M���s� 2q�(��-�_� Z���*���U��
��&�*��Uqnu^���eÏb�'�>6����rD)�FA�M,~,h��"o8�⦠yW�-��Q�0�~A!(����
���T���&6CB��$�#3Q�pm���+�2�L\���t��,=A!���T���i�
��c�٨�p��Q�}%W���1�Qo��d����d�A1���;��^Z8�*X���Ҩ�|]:���NȌͫ+ �W��S�ێ=(��q�Rk�ͪ)�x5��̓]�?�i,f��^���d�B9�2y�]5�����"�l~73�!6?/h��:]�
�Z�����v�
��-���
ĥ�Ǹ���񈨋���gwܬ�����`4b�Ke��0�li�IӅp���b������ x�qw?h��/�t��x�ٺ7�G�����|��dJ,]~'
�eSM����</�+�p����#��^�3tQ�03����#���a����w��9	���kcϒ�h���6���m�o�~���Q�i���o��Wy�IӁf��)�K5%�jɷ�?�L8Q$����0�8ul?�hz����xKmoI�B�j��]<��8�p�^#���ۘ�L�n�9��Y)J���U0'�q �-��y"b�Vf��]ާ�l��n���tY�8kV��$vo���Ƭz0<B����k�?�8�3ZzՔ9�ψ�5�gAa���g^0zsH,��7�_���Y:�%mK�r0�v���HW�k��LB�����̿���k�"��R�pG�[��o�}��4ɛt�(��Z*�F�9������u*�aݽ�U^�uQ��v����­僒B����[y�`g.A�@2���nM�jK=���b*�:�@J˸��bE���H2YV�͘�-��z�Vt��9O/���~�R�߮��L{bk�S�u\G�&�c_C�cjZ9�X��q�F�#A@��K�,d(v��=˦+�ĕ��/�=�,ږ�o�	�Uܖ�S�(��v)[�*�=`�o�����e�!����]�(؟�,D=�����#D9� ��_���,�p
@1~�Aɓ��f�>�����	���ҷK�~}��ޱ��ϕ9�V^O����i�|�B������qc��hb�aQ�,/x��5;>�Z6z��W;�����I�t�j�t8��8�s748��_@wA3%�P��(}�8C������%&�^����/ȱ�a�~�h�H`�B�]�v���8� ��o#1�$ŜtC��.�����=�s\ϝI]�-�t��0�LѠ�7KJR"�Oz����%�����!$����!��%<p�0��.vB���e��������8=�1������<��H���lY��SR
4��Ze�!ig"�v�xA��7y�,r"�Qփ�&r��!�!�lU�̐�ak��#PO#�����7�$����_0��YX�QY������7enqefZ?[�Q
;h��dr0���+�ϧ\ �:�x��#��t6�ی���}����CR��u��ecx��H���jq	�H�a�2H�/��^��#���D�
�<��)n��Z�:�&��}.�%�¸#^����Q#�Qڣ�3����}�XK	@�%a㲟 ��6~��c���0���y��pV���u���x>{�,�ܨik��13�WBk�j�5�Bcp�J��0�^�C�(z*��#�]�!g���eJIr�A�rno�n��B��?j�ef��J�f!Q�_�I[*��T��@zu�4Y؟{�fO���c�h &�l�>���\5́��Q<,}�(h�JRW�!�� ��?"��]�C09ώ7B,�4������t��'~��n�U������	�7�`�WD���$}�WFӌ���ʘ��9�@gQ��Z1K0ң�m+��)���nY�'oĹߏ��dcȐ�Kg�6�Ih�ѡ�7��(1��p���[�:��V5l)�t�^��������Օr~�NA����2^s�K�d����Nw1����9�-J7h��,`�v8�/E�i|
�2�ĥ�C# "��+RIp~����~\t���u�N۾�Ӷ0��8��s��`9�]YN�Re���6�h ��M�T
�Z��e֐�X��ު�Ҫ������{����(A�wS�X��d?<�T�4P{�1�OC�I��i0g���&���_�҇�8j��ڸCR�c	cQR]������	gL�;�� �F�,���]��]|���S;�3��hgI�U-�c�En��5#�������% ���vp���[̆;f�8�
i�6Kynו�=N?-���W4"Z��"���o3�U�Q�z�ZW>�O������nx���D��!��]�1c:��\��'�{KY��=����a�N�X��g }?u��R�XyC)1u$��о�&���
�;�*=TT�VL*B��C˔��N��?�#�(�ȸq{;?�W Z	r��v���T\���u�	��I�B� ~����̪ұ����05\řG�= �@�)!c�Ϟ������6k&��iV�T�_��-��;$����.[�`��M}��[u���I+=�dqu�l흣�p&�=._A��=�^�D������_*nb�&�~ٟ	)B�{���n���'Eb�0�".A;6l;���pY���+��R��C�6��δ��c$��Ryj;�FǩXx3�z�3x>M���Ȥ;��&,a�!m���S�~�dn�;��|#X���}ݾ�sQ�#�T�7O��v
1�w� K�W:=LΞ
�G���;w�-gc~vʐF�0��O6�st�!,퀦�_+�wo�Ͷ��VA���I5p��={c��ݺ��N�{2�љD�$�����Se��	����	��� *��Nz�5$T'6�p�^i=�i?�z1%��"�����،�nJ��%�w�Xu��4~�k8m���W��+�c��<IB1�2R�=	�؎q v�r�����R�A$����u4kHb,��P�a�9z���U�]ꣶ�1Ѕ�;YeF�6~���z�E������@UzT��-k��RS{U,0fb*�����eHy!pf
�=�/�ë���!�]K��l�3J��b8�/D�yf;7��K}+��b����S>���ZjL�y��r��/���3��.��Aϼ�jIqv��_P�0T
#�/n�> ZP��u��B���B.�F�wWZ(��
��b�iigj+l�{	����w5L�n <�����59�U!����s������,�*�T.��E���+吇�@���A�����?U���o��zq�A&D)z�T��XO����O�?�U�0��9U��� b���ͅt���p���`=s֝�J�5�
��Cω�J��V]4�j�B�&b���?�GE����U8���;��A����L�����k'y�	�O�N��>u�1��\mj&��eDHɌ��"{��X�<i���Xq�HY���i!a���j����ȥ�*�W-�k=�~D��m��?��l%\�x��%y���K��e���ߜ\�%��*A�Pv���!�.%牻'�0����"�x�)`im=u(ְ�@I����Fu�6�T���S;�$��f���>_�N���#W�n�i}JM$z��2�d/3>��9ȴ�({�����{�v�ABv�[�F0�1��Kׂ��)���_�]��L��H�\���:���Fp�{��ݼ��Ҩ�5����:��-_ys{yTg"wT2��37���>T>>� �3h�]�&�7 l(�f�v�8�<��)^�$Q7�d��W>��F�;��e`������s��]?r*=L+�'njw�\��g(�sa��c}J�����N���#(w�.���G";��Y ��D�]�M� �ᓧ������?�.k����X�?=|�oc�p�i:��7q�,� �g�f�8%�,őT爫	g�c���B	�U�g�u]�HG_�Е�B��>.>�?�n#}�dסl�!�TB�g�J������)~$5�����c�S��{���^�ߏ��F�ܤ�{�@е���h�6���OF���ճn^��sp�7f0��"���:]G��]�v}*�R��s��[n�g�{lF��f%��±p_w��C�P-fb�B�aa���P3�S��p�3�����J~90�h��+�Қ,��Qh�wu>��}��'�(��hs�`�4S�z3��):#/QW���q�]Y1��;�E^�j֓ȯ*���/Ԣ�W1���K���*t�Ϋ�Ǣ(���J2ԋ)Q�}���;���/We�GIGf������y�d�-3ҹ5�h����$^tT`@ ���tRJ3���[W��P��a�|�\@�a?��tL����b�>�Δ��2%�A�M%�=�hT�c����Y�xl���n%�T�/b���1K��,��v�Z��~��c8�z���8�v����{ql;b����}�WhF�BH|1��8�����̝�*9���/�6�6�z[��y�Z�@=c^��g���y�t�9m"`�y�h���� +ؑ�#J0%�܀[�hy�Nk����x|&ƊZ�e�s��Y���@z5"�s��x9�j�¡��C�f})��~^u���f�&Y�Dw�v���K������.��8�\�O?��}�Xq�j����no���C�H��lY���*�.S��"��#��Ҩ�GT�X�+��٬}ks���Yv
���i�N*i�Z��\���@"J�X��u_���=���t�;�]^�'Zf3#������N%&zG�m�v�'F��,\�B�������`��o�o��4���0�'9_+�Mp{i�cv���?\���IJ|ࢄ��,��ˌN��Ǵ� ������Z�)Y�{v�=v�V,�)��4,���P��-�����x���(�����bW�=�t�����/.�W����'a]����Ѧu��a�HV�y���`r�@�^�B�H/��� �ޖ���[.����}љ蹻�6�w��Ĕ���A��2����C���:��>oC�Ε���9��k�y���$�����Q���{�0-c�pq@�����ػ��_a��0#Pm4°)�K�)R�L�=�����_`�{�5��Y�K�ΐ1qu���`-��lx��&7BJ�� �4�nI�smeŏ��`��K���}�Y�Q8O�������欢�bo�t��W('
4+�{������p;�1�n��J�=ɐ]��G�����"d[���	xs��;�4Vt�S9���) h��$S�ns��2ETġ ���F,e����p�/B�@;��0�	�#���kf|�ʶ�*,
�L����|˟��#3|a�!c�u�H3���x8��b.��M�$��}���N �g-����~����n8���Ҳ[Ph���K�m�p�[bY�����F" {,A�
��,s�!.Y#˿H/���g��D+k`=f,y����Ҏ������U���oԷ��e�xI��ʸ趩�Yg��f@Ը�f�%
q�&�.��v̺T%���L�)*��<�~5@���#�`^�.�U�9�@�T=k�]�-Ħ�a&aG��U�î�����o�s!ee�0�����j
�3ާ<BޡÛ�^��
�����u�.����D�jR�/p[�w���{��_w��}�h܌�:�Tf�&���R�_.��ɍ���1�s�����c8:?�?Uz	!�ݧ�)9�ݟE]	�2bg�,�C�.^L���1،���x�6=x堇j(nٽ���ltf�Y���'}��T��[b[�8h8�=�9K�\-!X�`b7�7"5����J���H:_�w��J��u2p��l�`�Xh:4sy����
6p��t�5��zC�yu�[DcA�u�ڸ|N�{��uʲk�D�;Hzj��b��G{l,�¼P����^�y?��2@�Y���]�3m꧈E�"K�l�h��_����89|4�O�-!bT��6$L�!w�Z�&���673�Ճ_�8��K�v���2��W�������� �t�� 5�U���;N=�?kuk`[Z���aB�A�z{��|�J�:�
FIV��g���.��P'Ft��h�.������@�p[����Xx.�#��J�.~c��������S�zߗ����cm���R��� ��B`;J����N�@�̰ˈY�����&�w;��x%q�C�J��.	�TB&[Ř�a�q��l�$�I�y�+EFM���k$%���r#ů�k{;�H=����A��X�R��X0p�<q���J����!Z�ǩ_�ϭ-��Ru����զ�f�p�0FF��h9�.�	�-�|�L¨t9�H���Նp�8�}7���;��'��D�0���On�&��՝t���$o�m6�Y�.O�L���\�	�Z桰�����<����c�94gﰤ�s���R��uD�D�]��j��r�Q9޷x������2���{�n��R�u�� ��OUӧY�d�săK��L�Ђ�e���M@�d����ڃ�.��p�=���}�L��"��
�FD�8P��4 [�(w����W���V=?(��,N
��T��yL9Ys�5f�|���jv�Ɣ�i��R�:������f1T�Y�u���?�y�0p��r�2YL�5�'��vb 8�>u��-Eνt��Lz3��p˷�5DT.��+Gg#�j/}�������{�p,��"B��UN!�0�ai�)S���ZR���3-�r��O���,N	B��ǿpz�,�X�V���x���Y�q�ϒ������Smj|�.EKݖAp�N�uz����z������k`|Ʊ���V��:<���K�ǆ�_Vz<(�)Q�"3}#��g�}&q��N��i���3#�2�`O*m��?�kn�*��������A�Ǌ��*�yx٬�����r�:�:̳��R_>V#����j��3��dav`�n�>��x.�r�Q>�,r���T8�:����n���S��Ml�"J���=��z��-�8[�����c=��(�2�([�&�4�Nn�Qw���GUoI<% �JE;�[ו_�޳�,�[��qǯ8�O���XG���7��KQy�ĭl�L�=�[�d�>�Eg�מKA�G�
�3d�3@*f�L'Gܤ����-1�)K)?�JO���30��^�/�qeI����&m�x\"�lp��bc�Vv�=�M��^8K����Z,Bn�H��F[����5�A'�o�zM8�NM�ĚƉ!M�X��i���{�,�0z�j�R &��ǐ�a*��s��䎳(v"��Z-8�"Ǯ�'2��YV�ʠ�ۗ`��ݕ��l"���N�����Q5��w/۞3��}�b���!h��)�Pm�YQ`8���B�ީ�N�Ch�jwy[oǢ/t~È��ﶨXK�@�9k�����}��dvV��:��N�-�3&� ���m��'/� Dx�6CSl�F]��"�Mk�����Jr��w��K��P�
�������dT���4
��(R��:;X`�&s���.�ճ��5z9�>"!"�ݣ�u;l7�㰡t�f��_լ�vn�zث����7O�$��HM K��+���o *��W���W�~�N��!֫�waGT�i��~�X��6�C�Q2�k��/�e/Et��c�Y��(�z �9��7*�кE��1te�T�X��!��>0M*��%pH��);3�7�z��<�m��K z��8x��a	v����c��6�P���Z�\F4� �[�GqM7�\��;g�3JI=�RND3�B�]�u��s�ʙhRsh�}w�\�������	P`��`�+�!���Ł�diT�'2J�l%�C��+kZ�X�9x��)|�����:[D0�4�h���}A���
!�f�oKH;���ng��V�`D�?Wb#^Vi��NE���i�p�6�p�w���u�"�x:��;��讈�D� GA���5�||1QO������3`���K��%�U��6��*��"��B��bB��C�-:�SZ����n!��ߘ�C�u��RF
�z|+��AR#'�y5��$6�D�4X� J����3=,�2�/���s�W��z0� /C)�JiE����O�{" Ӱ�����eyJ@��N�Q�3g��#h%+�G�2�5ٚy���ޠ{x��E�y�E24��v����2�� �}|����,�u:�a/�HN4��{Г�כ�O@d�!��x9��<���S�D�񛆄�E�E�^4c�eF ���0#(�!�!�פ�E���1���u�s�p��Z�:���F_����Yj�(X|����ٹ����*���濍'��u�����˲)ʎ>�Xq��Vfk1E�F�-�C�=:/S*S}�����������RH���Dǜz��Jt��v~��R�+�9I�.Te7��T�/��p�� �j�"m0K�e��a�=%�K
>��������N���<�h�(�ռS95EVY���q%�"��A+{:͗(7��nB�2��y~<f��U���,p[����ðt-�2X#�����']�T������%p0���}�P��'u84��JV(�T���p�)z�ǃ���j6�%a;��
)�X�8ٯI�.����`�JQQڀ)����¤���6I^�^/c?I��)��&e�\p%^�ӋGdzi#��c>�J��hh����R�@������t�;`$��/ȵy�U�0$�l�'�3Lf�1~�^�T)Ka�=��p��8��<��:#+��VOI.I�yǝW;Oő6Ѯ��<N��_�v���Ű��/�ۚ���U):���H�L��m�3l��<,�N���k'(ā ?����7��<�$]dQ�è9Ô���8>�=���$�ַ�$Cq1�����4�8C�8W�,�m���]����Ȍ���	����F�țjK�횷!�ٔ���f��N0���^*ÜR�Ϥ0퓹�el�Wp��a�i����+�� M��g��6�I�#w,�1�>���]���s�����E�S*G�֋�]kӨk�Y�\�b�"�T����|v��*IS�i�����W��}4cK��G}����<}��+�ؼ{��u�v�qFT4Zl�@ݔ:�[��g5�B&��iަ�ɟ��.5]����s����$�j:_#Ё�A�-n�۲)�U{�2�2�HNi���?U�e���G�G̻U,k6
��rVC#�_F@b7:	�$�u��8�ݐe`�!ރ����Xލ�[H{����ĩ��P#�����ߊ�[�̚v���\�p\�c���������-l>4�a4�eI�%�
�f����Wl0��2Z�l#�Ui+_�lM�R��Ё��e���|�z� �TJl���\:37r*�P,tNJ�4. S4Xy]��i���mZYП���B�=��K�0Dٕ;�.fPG{K�ze;p���ӓ5-���Tt����Fcy&'�M"���pAcm]�[
�����zaD�E�~HA* gO���E�>JGm���B� "{Y���*F�Wh���)$ʝ�Yq�l�O�ٗ;��p��+�^ۀ��l?�ܠ�����.�x��ue�������R)V�_�pT�8��j%A�7�m`^��!��O+�}SA�s���#�jyA��h)���+��	���D�y�[������&zohݞS;��9>�����6��|�&1htޞ��l�'�x/O�w0��>>�q	�} (U����?�֖��!����Hl>��*�em����e/4$�Q��~���^4e�՚͢��8
F��W����ʥ��!f�τ�GN�V���kU������O�O�A��#v��P,�4yyK���<�K��1f���������ld��5�T+j%�!Ӝ�U+����U����x3Z�0���}�rq�`pq��RJo_X�Xj�
Vv!�a� Ж+��5��;'o�Yz��C�qf�FR�0��Aׇj�׳��2&��́����	�)�:�d����������'�DP]TṖ&	��\V�pa:p������: ��8�~	���� �<��Ⱦ��c}�Mͨ��Y�7H����5��BBe^��'�1�m�� �u�'�Q�M%{��⏼Ú%b)��G#X[
���A��]�֯M���֬@�&N���RI�Q����#�8��M}���[q��Fry�s���1ٞ��/�m�clk��ѫjI�Ed�:P���X_��n,�kD)3G���N	��ۮC�r��꘻C1��T���/�K�q��l*��L�ߜ��Ų9��P/���z����jM�����FNU
E��9bkj�.`[��58���/��ˏ�v��:+�I�hͦd�\�h�Qk���r��7�h6�Է|���n���W[��� �o��еu���N��nh5y�Æ�<��%�>��3��Pt�o*��ujAW�<3h8��=�X�.#����?�DZ)5ƹ_�N=y�^��F��	C���h����9�E��ECu�+��9rO�����l�AO�VH;�J��h���[�,Z���U!Op�*O�9G�QH�_q���NV���*�<�򽌼kѓ���Ы�j4 ʂU,|L�ok�c�d��4w�xg�ڨ¯PV:n/��b����Z%���MȾ��i�Wo��k+�V�����R,��|E4=�g�/8��4Z^�:��z�et�nh�^$�W6D�W,O�`�#ʿ$;7���h�e���C�_�j�}�����m�;���Ja�9�i&!o�ƈ�I�&�l�T���T��~IF��f���%����į�M���i��EPNT�P�d�XYu'E���n���э�{1����P%2b���K
���"�h�E��IJ*=�[ۃ��PeƊ���"�a������8̭H�=��*e��:{��w�e����;v5Ya�A�Qv��c@Om�D�l��Ŧ6�۰��9�H1���oi��ܵ2�%O	��G�����,�YIF�*M�A��W���ս��Wf5a{�i�"�7���l����a�n�&���Q�D�?H!��n�1�-ޚ4���g|R�@�Ԍ��s�=K�C@Rn��Y�[���� e�����fX�,,�Hцe�2�F�hc.mH���O4�h6j2O������z���3��i`�I#a�+c`]�$9��cu�����)�`��.��!a�A�1��&����L^�_�e�WL��+��H`�ihY׼r��,�n�&i+�۬.�fJ��S3"�IO"(��D�}0��/�+��i�9	m�D$PHO��B5)˃ߎ���	]�f�h#ڄ����ϱֲà^���I���)\K|y�vz��P �K�g/���-Θdωчܱf��gd��.>/b3�9�:�0ő1��F�j�}�q92������N�5����F�3)U� E ���m:2�uS�,�Á0ϡ|砺���� �=�l��j�vǅ�ў�r ?$��\E+��Z�o����_���ei``-����̫J�$�`�64����H�#ꑞ������AX;F��!�Ŋ��@�Q���Gcu��b�T���RBn��3L��v����~�Gi�uUO
jj ���0��nt���s���6�o!ֵT���d�F�Dk=�������5T��j;X�?����
��9tb��O?�����<�y�.$���}?>1��I"r�3��k����4��C�U_�;mM�b=h&0+{k?��h72�Q %��š宽��O��;�b���]<��N*4YQ�'���p����}�g�HP��p��9qǦ�dhY�y:*T�� �G}p���j^�b)���r��cw,`�QW��w(@��I��׍M�	��t�}�GBȮ���%e?���7���yd)�2;�(��D^n��׼=�j��/Iy�F(���)�.B����jYh�d�js��#�t���\T��b�_ۨ��6����W�ܟ����L�IГ2�u{�l͆rAfRi�r�n�{�I�Yx�>�,�r��O�&V9j� XYx�+2?XQ"��V��p;�t
k ��A��
�8n���A���O�bBR���{ m�|��tVgx3y�j�8Y�#�(���uh�MX�
_���b�����~wD��%gZ��&�$����b=U7 �虬Ov��QL�
�xF��lh4�#�>yH�����|y��z`�=������w˷8D��DPV`;%�/�ղNf,)�HT6�F�����JYmq�w=S��'e|��Ru�F��G�ˑDg�r��:���PO��P���)+��A/��_���Ji�'���n��Zq;��{BeGO�ס�0��+�������Y�&63z_ZA��~��_`���Ko�d�ru��<�l��@g��l~��<��ڸm'=��]
G��'������y���?��q&�17��� ��ԧ!J�5��]�7X%i(!~b�~����L��Y�<�?yN:��D������ 0ا]�,UK��Ռؒ�Q��Kȣ�I>�	xw�Jl.6��X�{�(	U=W͢���i�"�v^�.�H�(.T���;�j�ָd�=&s�~҆h����2Y���$i�U��C-�^��q��(������9��l+���l;���PY5��\R���?&><��F;Ô���LJX��6�Օ Y��	���L'|��[�����MmUcኚ��;�t$m�=tҏ��F�Ln���l����(�,��/�ըY�HW�_�]&��őH���?��+��Wd�l8hr�����q7���칠��w��}�Zg���/z�PV��q��R�ݯ�ϊi*�
!�4��;��
��sm�E��q�ԣ2I�G������nC8��7���+I�: B��,+j~�ם�J]�킘��rkp[ ���Yi��Q�[�+9���,Y�i 4D����5}���w�~��t��P�
 ��6�B9�(��0�1�~D�-V��ɗ2.�f�>R8O(vr�č0�6z���Cf=K��U$��T�%�8���.��nf�h���p�]�4p����("LQ���nW�������=@J;�M�ȭ�\hxs�8���x5��_+ZW�`I����/8�+v�IX��ɐ������^wF�1����\��i�60�S�ڜE�}� ��`u� �Y�ݒ~�Ubi�Z��z��A#�у4�w
#���u�=ԍ5Crm�7�R�Ab���.,���i�|H]BIt�_(nL){`�D�A-���S�*�
�Q��k��o6x�$�=V'r����hࡑkN�+�1����'kw#Wur>�m]�%��w�6T$��E����9�8�Q� e�=�\۪)/V>�n��j5�
�j��X���L7B�M��Q�N{MI6�����7qU//K���d�~#:|̓�-uGܭOW���|R�5��$�)��&�	��P��=��Y0Q��<��r:ju�ӟO�4�Zn��1�d4�H�#SǙ���e�-j,Y�h�~|��5.��ep���"Z�?"�c��UpN�;[:!���`���~������yy��u�����b���Ϩ�\���i^��ʽϟU�$��|7mz/��σ�2�Y�v���=���KS��P�|�]�a�}�K�e� ����%���M�����D.Z�B���$O���Aů�������s߈B]���k]�f�� ������[lcn��
]F�	S]��=�|o� �_r�?�p3c��C>��u��u�6+�� �ܑ�I{�k��������/�L8
R� ��u��w�p��A�g�F�T#F���S����IN���q.^Ms�[0 e���v��|��ͦJ���W?��Tk�%�&����IF��_Ìlo�h鳖U�Z�@jz �J@��}ׯL����X����È���	+�l6�Z��b?�E<<T���q�0ϡE���J�+kkvJǖL8�ǹ��?b.5V�+��I��Jm���K�>n"�S2���2Dx�]櫢��oב�.#h]�K�"5�x	F?SK>���HǎGV��З��U��5�\`��d�j0���XF�X^�.}����Ǣ��6 F�(�]�9�>1�F�gP��M헫yR�\�-rPTs:ģ��.(贏�P͈�PE�
`L���W�|0�;!�@�øJQR�^6�#�!u�r�?)
+�_�t��Þ�A�\����*b�G�z�{d<���ֵ��ɥ	��__�6����� �	����֡� ��]n�j����Z,�yZG��p'���9�>����殺WӚv]���8͜�U��+�P��S��$b�6m`�D�4P
�8%�����8�O��F��Χ`[0����;C,fӫ��-�D.Z������3�E���9�^ț��Kr�7�Y����k���&Q�p�C��ko���sߝ%9)�q�ɡ�}%���K�#R��B7�c��Ge� ��xL�5ux�Xs+�<� ��~�(��P	�6SЖ���8�5��(�,`q�l�b��t��)Ej*�dx
�qbA�0�� ��]�!kivK���"�U�y��K�l��q�4�C���g6��-���;�}�E)&/Y��ZP+�T�pa�%�&}��J�����vɑr��fFv5�� [ݍ��)<g����	�$����$�V���d��}L�����D뭿������kE�j �"���C�U��,v�:��9����,��l��1�����K����Y�G�2���p��� cgi�`Q�9|��e�+��,������``q����dY�4#�\�T����
��]�8X��c�>h�RH��^?n�i5�p�Z��\�V,��dm+�j#�3��Jl��7���"U�" �e���h��/�k�R�xT��4��v�`�bx�m�u��h��JP��J1
4�n����@f���B���ofI�/���&��k*�,H���M�]&���x
�-d�@D�7�qȐ�/�+y��뮲|�z���zkr�M[�NF����r6���>�'��!azL�N ��������
�"��Bߜ$������,�Ť� �e�C�3��1���ť��RĽ�I	��L~�y�~}S%�	٬2m�{3�`F<C-��1� �&�{ƌ.��p�d`5rۭ�Qv��}�_�tG��f�rQ��U"s����J6����/��4X=�wj���rr�2H��ߋx���:`��]�F"v�en����l��4�:H�q���6]���
[a{�F"�Ɠ���G�L��
��_����I?��:��*��oN���I�P�}l饭�v��/q����..�jfʭ��+ͫ;""�By���E�.|���6M�[�l�:Eo}��������?�?F<��\T)��M�HQ�Gf�s΢�Y0���lL.���>)8E���Y��	����;���9	���r���+T�Y�K�.cTy�G��d'�o'��bk�*�d�6�9����Y�KH�����_`�q���5cO7)n�������Y���?M�J����s"{5c`�1�CB,mKcQZ�qd#3���Ü��]>gW��c uV�H���}�����( Ԛm�P��v/��i�4����:��rcG��o��]~a>9k>	+LbY��a�̆L��P�@����c�1��3��>)V'7��ν��||�5��d��FÕ�j�+3wG�Uy��v�sq2�o�q��ncI[�,F�N�f�j���[��BU�_�9�@�Sgde���R�kM\�71���ǃ�2OX��/& �Dp�/��WQ�)ϱ*��ň��Vٔ?�k՚[���.�~Uރ�G��#��C�?m2tx3�.t�I��`��T7�%���j7���]�7�]`���>EP�D8འVT�ٷ�e62*��8�s&0��f�e�mY�ϟ�$PQ���Gi|�H�!��C3�Ɔ3��^Cm),�Pk�����23t��سt�&H50��.�0���z�(m�������8X������|��+�U��jԲ�t��}�S/l����$5�ڸJYn�\��$1a��c67��X�'�U��I"��>��Ɠ���z���5~p;�(3���m� 8N c�l�깪�C�y��RyS�{��:�9z��	.d�e�+���
��e(�]�z~���ָP��z�����d�dZ8��mZf����<f��;ʆ`M�*�c]�2��!�! @v��{��֟::�/cܓ��c&��y�^̈́ـ]�o�G3�u�Ѩ���|/	�T5 [GF��2�Kl�<o�D\����8�,�pM�f��%�e��p�וt�>��4���K��J'�,Д�Ñ8��2��A�^�����?x�Ր#IǂU�.��� ��-N7�1 ��N���{a�!����=݈>�"��N����77�09 /1]	�#�իr"�&�R�E��}���Yz"��,���J��u�ɛ'�/r6��x�Ǿ�H[\���ߒ�]؁N�w��5k�r5A���[�]�`$�C�#Eӟ�GL�jM��^j����>DS�6v/_�g�,l�M��q����~���@嵇:���8���A}x��<恌�����+	'Bv���rz%E0��`w�QuŠ��C��x��0M���S;i�-���`�]�����{u_��
^Vq]d2�i:��1�bIVn!
��r�-B������%��Dֻ%D�S�p�4ǽ�0�ỹo��<��3-E���@8�i�(&�r=~�;�3t9HuQ��ܰX��q��j��u`E~���bw�YA`Yk�"������FTjf�l�wП�4EΟ��t�%�">���5e�~Gξ ��w]���Z��㧺@�?�cX��Q^�T2�2���Q�U�Y$l�hM^ͼyw�e�De��i��(�|�ԵŔ���|��f�6!^�ץ �Bf�l���ٹ���9b�|�RنWݰ���M3��� <|^�쌧uss{s���eR�u%��1F�ȧ�a ͮ�����.���G���`�Z8Z��3�iOϲ��[_O\���TdՅ�T)��t���Gc��۴��18(|L����(H��y�@B���U����� �<��ș�fl��V�O����Q���+�F��B��g���W���ÉT� ���i~��O���B��v�u���μk����>�1R=$�4WB��7 g�Й� {�<��>�X���8�s��=��[��B24�[E���1�����C7�A����H��y���)��ύ G�^�*��k���������a��E*��X���T9�F�}&I��oW�h�N�m��!ə-q�f�J6�%�ީr��Am䓠G��X=8�c���I2��P�_�,\�N{*ǝH\ό�(�M����B�ShyZ�{�s�K���~+��kD
��|<$��'�ĤF2�RFt:G�R]>:�	�:��;��;ȡ�$EF9�A�.&�lX��͡�lD 	!�����z���ɻ�"%�D�lhX��n��]-0�G��|S�g}��c;gЧ�#p|��"-S��<�M���|���ؚR���a����f1�7��1�\�y��t���1���}�if_q�7���G���>;�DX��:�����R��s�KM;�u��Q�fo��+	q�
��*uϽ֗����&A�2� a�K���}/+.� ��x@B!���M�P���i��=���4��Q0�TëOZX�J,u2�նR����l#�õ]Ou����f�������y%7�0�Eat�Z�!���BI����T��7�QG��qe��q6�wJ�KR����<����T��̰�E�Ӡ>���x��K�c���|�;	��{�|zނ�	rɴ�7��� B���el�Y���y͛/�<�-r�B���ˤ�o��A諟��7� ;�˗�"%�O�H������ho٦�Ϣ�r272.��>
�[���si�P#+��c�U&�;�w���jR|�xQ#A�u�U���ֆ���7;kd/��lI���S��~ʮ �tjm,�(�"�\�k�,EE��,���7�}�euk���MR�<E!̢���0����O�s��{�Y�����飆W�C�(Y ��F�Ki0�yGP[�@�H�L��?����qZ�+ ��DPp���-��? �� ���h(	����j磚�U�	ּ���gve;$
��׶�@�iҕ�m��%���!^ Ŵ�X�8|;k�ua�:�����[K`Z1#�o�>
��@��3���4:�4�.�8ۅ3���!�U"ߠ��yp����!��;DE��]É��tDu���ȿN�H,���e�Y�I�~��|����x�D�NP�g�;ə_�AXO��i�D��70;?C�IFBݑ Ϗ�]�ٸ~�p�.S��F?���Nsv 9�3r^�`#��Sk�Tv��?Wn�}DL��8,E�t2x'��5(��bq�)���l$O�����+��5�v�ɶO��R��wS����2p�PE	����9a,Z�j�e5���̵A���M�$8�Ըm�(�1�|��%0�L.*���6��3����0_`.t3؟��!�\g��Ro�͡N������	��z�c����I�+>�ܫx*|i���{j,��X��M*�G������\l̺�f�)8FEj5��6���h��S��jC!r	�g�Ѱ��I;ҵ��H��Q�l�(���BAn�O��f��q�a�KԦ�t�9��jW��눉HR�Hv�A��#t�[*h:�� ɡu�?�rz
T����QvПCԑlW��bH����c�B�>�/-K�x!8gl��О!զK}jי�n��)�SG3&��<{��l*��2ۊ�5SJ������演�q��C9)�n��\dd���`����Ճ4�� ���-0�)9k�X~V�V͆+7�v��+�}�<��x��E���Ә������pRi{��jq�����+�֗��Uk�v7�Fj3?n�B݅���d���u@�����k�tN/��,k�F��7ˊdP9�q�g����O�S#
Z���xp���.́����(��AN��3���Jj\��]�,�q�?�9�=�Ʃ�)r����b��ej1md�����Sz�:���k��R=$y�	�G����UQYtr�	� �zP;Q��	0~J�+�r"�p�?���7�?��E���'��X�5$�l����)\���Z�����'��ZL΁�]x&�|�&��n��ĩ��,�h�
�"C���RT�+�h�i��D��/��X^y"G�Vֆ���5���G�(�%
3�G-S���X��{AetR3$��fTJ��E]@��u�c�G��M����57�PW�w�/5���-�`fu���a�'�Bf� -'�QBQ��w3)�
�%�����]��i����Gٽ'4:4:M:��V1�Gw�l�����*1d�nG�2�ӾW�֗��Y��)��+�P�_`���#�l�����wN���wk�]��B" ���ݑ��pgQo�6޷οg��1���Fd@���K;�/��Hf���Gw^�ת�X��s�㝻����#��T��R:L6���><�� q)�����wc`����K����7���d�o��J�%b�X�k�1��m>�l𱶥2�p��Y�
�n8'�W�3�*�H�o_���n'%N���O���*�6��4��~�A.3��&�z51�{D�Md>@i�X])DK��L����3I�$kZ,��V�h�e��f�dg�^�������ۙ��(�d3���̟��(�E6���`�7?�^�v��52ҥ�M���Q��r�N���yN4�c�""�����1��L:��M��f�ΥL�,`
	fz�e\�*��� �
�؋ի�ҽ���iСfJ&4��*Hߑ��q���E,����I�$+w���]��ƈIc���Ԓ�$;lW�g�R�?+��ݪ�m��#��U����iWa�p���c���벟�/��w��b#�K^����8q��'
Ƃ����h�`l�aS�WQw'�篑��]�$�(��@�	�J$7��PLQ��f�t_�d�ټ�Q�/���"���%�Ҿ�S���q�x�3�]1�[���?J�J�ӹ��r�O���� C�<��C�f�&�b6A�e(�zIq4fB�cV/�������N'�/���L&�5��Ŋ�����x��� ahkB�v�m�������(��V|��:?�KgaHBD�F�t�a��Sn�t�������B��$T��"P�F��a�Ó���"�#���r��4B"��UR������[?s7A��o���f^s����H^�~	�����5W���P6���|� C�Z��{�w.h-�����d�t^����`�a��D�4�V�f����N)K	p��m�Ͼ�e�v_�-�^2r/�C���)�L��yQ>����O+�e":>����ϗx��z8~bs���,Bj$Э$�.����`����<�B?�^�}��d��A�XxwXA=��uyz��ԯ��b���i�o�I6��_����(�J9:�AS���U�Z!�� 	���V����O��&M���ގPW7g�=�M���Zs�^��qw�5�H����eOj�!:�DdJ@ڢ��b3��~����V��X�(󁎋���Z��j��)��e��˱{o�^�q���S�#��J�_�HA��	HG�'5]5ٷ�oQ�\�g!1fM������[c���C�/���뮫a����z�(�ZG��*�vr,OBUq�V8hu����$�ΰ���Z��[��������r��U�8��y�hz8��P�U��T@�3�'{�+�q�#DDAˍT���_���|�A%7����O~?w����k�7�ʈ�kK?Ӑ.Q�)R���L��幧��hk�e4���^9Y6�b8��N�gח�e;L��>|7z���+r��þ������
|�{i�h��'V��m�҇�|l�B3����U]()���4!��^��y7��]��D������/�&"WU�]�WTU���b�jd%�#��v3f��Ix{��s*�Λ\&������,c<�2��}q�Z~���rg�t�w�22�w7h�"�M�g�C�9���7�e;`��y̤o@\}?�Pw��� �"�a����O4�5\Ք�6���s�nne���n]Gf�-���Y�Ei!��J��\75�s��s�yU5��������vԩ�"������/��..Ԃ쉱��O�	`+�]�Qᝉ����ν$QI�Kc1���2�?.rʤ���'Ez&�UJ�ȕ�Sd�3�}Q�N�C����I�*�_QO��)��n�d��jm�%fxb��1�wBg�OH�a��BE7�Y�Zb��IDr�J�x��h]��U�I�,h|h3�2C݆:5 �"Ǭ�{�'d]V[c�f�T^�-�����a����ɬ�@鲍� 3�Nɧ�W�����ReԸ�΂��%$I'>&�����N�ޒ5.��}��,]�XO�+�^�T7���R��UM�䨲�|ǁ��GiY �^ �R�7��Aܲ_~ĝOC�XEں%r�J�m}*�	����)�(HF�A�?}�ŗ��Iȓ�_��#q�9cFx�j0֋�or N���k]%�
�P'���v�*�c��6Q΀��*H��U�����Phl<�&�l��l�
f�[���Vz�CC��Q��o?�.��3��9�p��EمR5fM39��3⍄�n*_�	RJ�46� ��W�V����cp�)h��-C{�WƄ,����!)ah������RC=��A�@�x��U����f�G�z���GǊT�xb_��wl7�ygq�����5���a�A����8�p��v¨=�:�ں�i�8���z%`��ͮ~�\�A��H��jf��-v���~_��� ���ΈA��ڼ>�j'��[��#ZX���GNbˠL��d��j���Y��d7t)��4�z��B����cn��B��l@w7)�'\i�����CU��ˈK2�}�̠�d���_�M]�k���L}����Į �T.�JAu���<�����=N��^R$,�Қ��'yKQ&�bFjrۅ`���`c��|���߀)	�U�Y��M��}��G��R��dp�������J��qM�&��j��t��T�!���htʫB���й�'lC�Iw;�,��Ɓ��&�x����A��.縴*!����g	*0�C7��]��{�*��g˰X�9�;��͡��Ʉ1�s�kU��L	w������*F3�j�F�s�[Nć#��/��Z��9�UV���S%�F�v��[�|�\ɗ�>&�گ$r�\���Zr���-$�2�7��d�QW�6��s�[L��'R�S��T����:�sNN�}kn������J'��L�#�֏��+����j)K��ܙ�D�(8�E�����f]y喃��D�����8���r�4�#�Z��kEf�X�\x�z2�T��Y����� W�W)��ОȪ������o�Զ�~���69d+�	��aЦ�LgvČ�^��H#u2��(4��ER��GO4s]�Ί%iVl���ܫ��]�1���h����h���A\#N} EO�����w���{�ߵk��qb��[J$�!$�Z���6����=�rS���'�(>t�+���L?���W�_�-E̕O���߁i�
���d\�䳾�;�n���k����׈���~��ʄu=��m�K�D���[�D�n�IR�\>��ţi��"Ul�&��1�ŝ���z7�[Q��qV����TDݡ!�����T�C�M�/V��m���\b"K8֫��X��Lqv��S�.ZU����4����!��^�H}Ma�
�I��	v8�{����+9!�2��Tnn��X��Wac��8ʹ��)���1O���j��1��5��W��Khx�Z��+�#�9���BMx�t�s�Vf���@ ϖ�ōS5����'f����u�yQ�~J�΅J��z��\4�D!
G8~b�������S2w]XX����ݻ>ܶ<̰�ѓ�R^�D'c%�Qm�,�\./��~b�QP*��PO����س�u�d�1]�ǫ� '�jf���N�u�ѡ��sHk�$ٹo"��K�4cZ���3�)AX������e̖	~�ò}�;�e�I�N7��Z`�x���� Rp�&_vR���jktg��e�]A$1R
�;�=�>��靼�4d�팢��d��]>����
�Aiٮ�����?Fal[L������ͬ{�ʒ�fS>.���XS=�kl���2�1����-���� ����U��+�PT.}dJΚ��8����@p$]�e�p �%��ڍg��������x�]Z���6��'ʯ��X���Q'����k��Gb�a��F���a뽰�a���L�i0�.=a��=�$o�"'���8T��^Xf٤�e`�DuDwr�m��&�ݾ�y�&��w\U�̩)U�!�0�m��H��,0��n����,�����#C�vtmZ;�æ�;�����ݑ{,0c�o�Pr�&��L�i��+�/���}�ƹb�B� ���<q/� R�-2p�l%�x��a4[{�=�����ڛ�7/�fz��+�'����ޒV�-�r�Ω�<��0O��=�2�'}�(�;��`��W��c]*@��a@���hH��b�_꼰>@:!G�XQ��wZ�rctK���V����t~󱬛4��4��K���a}��ǻ8q	��!�刂Œ�b}� q�ij�{�q��:K>Y<~���γ�g䖷����I���
�S�3|��*>}��Ih9�;���D3��nu�/P{PC�h����/���W�ug��?��"�I����lO�hm��T��x�Ӈ7'�ID|a��r@�w��wB&[/K�,;8n��D{�sؤ�x)�l��9ѻi�����H����H�W��>��F�5�Ol��糺���܇��zZ���-���[9*�L���%#��9ˊ#�>�ԥ�퉔茓��|��q��q�&#OU�X�[ �:��D�vtd�	�Pa���DA�wv�3Q�Y��k�dM�e\e�㒘�q�y��²}��t�y����`1�����P��o�W����V�� �g�lx�&db)�!�u2��&M��<��B+�!��g��H�]�u;��_�J|��}f/,�%M�T��!�O����"[\�qK�%Ռ�Da!���{*�q2e�;.8���Y&��S^wğL���/�U1Խ�����ho�'�.�S-����m���{~�eߊ� Vtq�^	/ι��/6��&�IȷU���**��,�|�Äc=BP�]��8Y�^҆d��e�u@���"7 �O8��n����f�����vEZ ����Dt܀5�W/�wF����zN���mE��K�>���#��fAT���.{�w��V�Ʋ�83D���Yh���Ll���	�5e�g�B�S��̘�^�7���)�<�po��r��Z�#�^��;)��
~�kZ<6�:ד5������rf\�o��ҟhc=���(�"I�������=���ܱ��s,���ߍ��/�e�F!�o���9�����b`��&F��V��I��򢮌F���5s��"'��Wg��)�{�8$a�z�\�.)@x���������5{�kSA���c�<���Ě��'��;%�dd݊aA�_�py«}ѯ�9K�9�s߾��$iC���Oઍ�㓸�X2��M��H�-�A��y�"� �t��dp�h�b!�0uW8�W���������z� �:q���n/�@�N�xԺ���X^�R�!f�z�E�j?����y�v��Jpꓹ��젾��tԋ�$��D[��w�"X����y�vlz��!1�����TDg}���1��"��Zy��_��3|���<3�!�ᄠ֑�����
���wI�� ���(4ko!m0a��1|J4���J?��+&�T6nK0��i�o�ܝ	v�`S���uoF�]!(<���P�)����Uc}��]٣Jm�0�� �ʬm�񻄤*I��I��n��xX~ ҵ�9��N�qJ+D�h׎0���DG��{(�tK�g�P�~c�=Hd��M��	����S���s��)jC}����?#�"á��h�\ߺ:[�H��g�7����+�sr�]D�ٚ��K�����eζ�^�ˣ$V��3�<����_��+���4���n؝O�h������p�Pw4���X��cL��vf�ѹ������̃o�h-1�>=R�`v��s��zUpb��h����J��������@�������4�*I
[w��\�յ�����F/��7��w��B54�<��cf�%��8�h�]��^�o�{��-�D�m�B_[2�e�Z�p~� �k-�-9�nC�)��ɹ"e{>����KyБ�2�ƹ��tWp�&��N�Z��
�
c���?z��[d�voFp"P��]�Ƹ�7V�3�ߞ��,=��20�J�}��4e��c�ʁ�����S�k5X/0��������H�c>��.�U�J!�B�O֓WMi�{8U�B�/bl���MoEJ���T��t���O�H��ˇ�9;9M �xa9Ţ���E,�l�/[f�zG�����Ĕ�Y�Xi��4Cf�3Հ�L�u�vI3O����x$��.N'��;�-7/Y�v�1ëN���\��rL9NW<������c:∙�{GSH?g� �>�_�+�'�s�֚u�fҽgU�=�v�R
h����"���WA�j��9nä�Oz~��"��5�5U��(��Iү��$k��r�"�z�&eӿq���}�v@�2%AQ|�����F^���[�&y�����:Nw8B�W̽�������"�዆ϭ_�.�"�d�
�J�gg.�4Gp��?�Ö��vk�w�����c�|X|a���_�#_I�����o�]����%�ρ�U)�
��Dv4��9A��@]D
6g/؃�J���������8��Did�c��B�2:<"��fZF�_N�($�W�|�6Vm�a��j�6WN�s��3#k_�H���|�PRf�ll.�M7Gބwx����i&
{��tęZ,��T˴=	��,��_���'AW/���X�lik;'��#�N#�~�4�[����4�3��� -��lB�G��N�y?:X�ޢ�5s�v/I��i;��h�
hED�i�[d�m�:�45K�̒9�כ��#�ct��qCQ���42$�;2{��9d��g�%�$F$��������W]O��E��3Lh���_m�,*��' ���Q;3�u��u�RؕI�,��_LP�#���Up�7ki�E饌�r#��0��Sk4	_�)e��nB�Y��i�!���	���Ɯz��j.�6�F��r"�/���qq�Ǯ�DPm	��œ�߲n�����Q��Ox��j$+%,�(u(�y�P���P,D�7�t>������;Е��SO��=��t�J�v7pH��T��C��'���N�VÉ]��=���Z8eg�K8A�Bb����NL��񏝎��pPeU�w�B�r�w�9�px��>#�C��C\^��Q.z��>��[�Sow��`lp���m@�����B�E�@Q]���:i���TT�HU��ێ4=)�o�Y��G8��vo���8��C�ms���OՎ�
��k�t̞	�5�d�x]��w�;NɌSn 7b�?��x+��Y�w�����kA���{��RD���0�U��ǂ�B!)��Ć	G���T�5e��(w�qڻ}�Rt��39��Vcj����Q�*����ԯ�9p#f&�`�&��@T[�*��q�q�2[y`����n�OL�ݲ�Z1�/��>�#�f�"4�`@}<���d	|�	u����iŏ&(�y`��m	��jPy�^A������}�M�-�1\4�m�OD�/0���h����@��O�)>���!CVZ�(� �#|� �����>}!1>d�Į���n�S�`��c/#��W�^�0w����
�s���ԓ������p��o/���p*��Ϯ��T1ط�E76|��2��4� ��;�֔�c�]��ʬH���x�䚆��Nsf_lߙ�9�
��wb��ȴݰa������-�9�����I2����(a���+�x�Z��@N�e}0�$䲄(U�}�I�$V8�mXF

�!6�iB��~ ���!�N�N�����,��*�l��?����^��}��!w�tL�TPD�[@���,�&^��b���uA1��;�,Wj�qݦ5��!(�~+��w��>�e�/˿��Ǥ�o�[B��K��Ub�����6���������@�f�]�f�Nx�cp�Y2˄�d����XU�e��cDe��H"_i������+�\��Y�Y E.�ʑ(���Z�$�G��� �,�͋n~�d�!�����Z�e��Wc�
�$ #�:�H�/c�`�q5t>Q�J�O"x��*H�f��ƿ��gީ����V����(�r� w���������E�a�	r2��ˎ�/�c�ɧ��3.%w�
��Gnuٍ޸��E>�%�`iۀ�MO�����9���ES]KɃ��C%�rU���SAo؂�u+�x���W���|/&���� �uX1R�)�ÿص��%��9�S�Z��Xyy/�E9Zַ1'0�$�h���ǟ���k!�:�$V\�~��L�_����l��Y�
�lmTyo���o�l��������I  �e �V������=��&Q�?�n�Q�{N��%���;V\��{ē� @�U�J"ETa.��%������J��8�c������j�_s��#�)8$}�y�Aw�QT!b�o��`��\(c�ιy^�	ךg�*T���W5.4�H(����%^��?2R_�ų����cL�J�s��k�+?�׿�@ ~:��ޙ-�[�E1!���p��J�1� t/G:^ �s���eW�����b�̀i����H���4���f����}g�����S��E��u��K����MRX�%��l��/9�����.�����'C�����>8^�m����0�D'�|��/W��Wf��+�~�}3�(�r����';)��jw"[��0��Tg����L3U�l���c������_�7��V�6	puG�ŐP`�UHy]i������P��k�X��is�\�h<t��G�My0��)I�e����%/�u~_�o�Ѣ���62�٘/��ռ��>}��b�����}yY4;�f3F�mm�;� f���QaYW��3+��0�����e����,����{�������>�J[L��!�P#遛ʐ�١�eu� MXӮ�j��k�u�ԓ���S7�;�4�!-;��P�>���Y�����O���Lq��>y���(6B,��Tm��1�Q�u!Q�{.�!�1Mp���]Dp�`�q�0��g3����-����M������قi}Bz'����AB"�M3J���� 3	$N���&J�n!��:�uX[��W^C�B����̗�(��gq	k�4a<�5�{?�6�� ����PM"j�`P��=�T�Uc����~m�WՍ�@!���L0:���?+�P��𬯩���?�?�'�1�՟c4X4�����Rn�����Av樫s�8*��b_$�����s���HZ�|���Q�RTW]����E�_8��m�z�W�}mP�J�C�� �nIi��o�L�R�Ǌg�0��n�`G���[e�9R��u�S*k@Xӧf�W[�� �a^ӽ"�_-�-)�3|[��Ft&�cx��h��hU����&���u���5U�h��p��!��Q+��ȁ�LY_����[���+����!�(���?��w�>MpN jBјe����,��ΌXS
���5@JĘ�--�V�����;MPA+\PJd���:���(�olS�=�>��H� J�Vt]d�|�Y�1Ҙ-B�Z�c)�T�ϹUH�@�E���S�*��.�d�I����njr���d�T����)5W=M� ��t��(q~Q�g���(8�˩�V���Ejp4ŷ��N���Nd.�L��P�=|EM=�rfb� Q�S�>J��C�-BU��y�����6�8x��o����j����P|U]6*�D-�8�)t�`�������=7u(R�qJ�^7��W�ڋ.	���mFn@|L����h"�4��q�*�E�����D�T��˪̇ݏ�z���%�e�t(��4�S�/)����L��tpH��Y����Wd��	�����x�� ZJ�ִl�Ԓ��{ϒx!����*��ۜv�}����T�/��%S�����(��W2�P�Xv���<�t��h���x��~r������]���[ҍc���VL�?F�*5���]!�4�,�5Wr3�c�1Y뿴��'~V���|`��ZM������┃�)ub*t�k7O�)[�mPya.�uI��*j��0����m_Q�$G�(Li%�.uA6#�F���ߦa>���6|�4m��/ٌ�'����A�j��~3�C��Uf0+,/�D�輐�#�7`�J9�M�ya��� � �N��,r1'�鈅J�k6��m9V�9�{�ź=���x|JQ���񮍴����Ϝa�Fʢ2AZ��=��=
��yY3�a����K�`�зF��w��"{-�4*��/&qUDJu�c�ejF�ɘ��!�i�v	=����FhD�]��r�
�1�vc�B�dک`_���1��8%�;�o��Ƶ#��l]M�(�8�2;}�{�ֶ+_1�Mɖ�)�}?�L�ʭG����g��7��p)��KԊ���p��ZLO�N@;���>�F��!��mݟH�Qv:�d��[�
/*�;?m�/��?�����G^�3����/����Be,|`�ۯ�
"�_�����`��O����|��2�7�E}�Y�y�2�.��h��-��t�rc�/{��x��Zp����v��¦G/n.3��,�v���wЭ�T�6P��c,��D�@̀ղ�r�M�N��+ef�}���l���a�X����'F:�t5��CK��H�D��յ�qӖ~
�MC-�.������'�09����c��V�P5����t~=Fx���iF��mH�<W��<�4g��1����g����*D ��jmҫ^�9��Ƹ��(�\U��乶���˔��AQ0A@"'%�:��p)}bM�����r�E�5NH�G�z�ḍؼ>��%Q."
l�	�[x@9�0C7q��G�b/o��
���mz�;�sF�]vJqy�h�kd�����T�b�k�k%�s��鵊C�YOܶ����Ok�y���vit|��\�S{O3!j�p�2��9�*�U{-����܎���Md�����[~#��ehg�t�yX���IZMBi%�0 ���rZ��v�)��]��m�8��%�}�}fT�ۨv&Z�NZ|4�BN5�����'ńB
�}�|�,2+4䎕W�m�+C>��e�0�u�`����T��DaX� ���m�Z��q9�����Brw�E�� ��9�݉��Q���N^�;��;��]5L�s�N|�N�4Q��c�9��,��ns�驀7�L��k�:�Y�M��j�R't T�"�J]�X�G,�R���
�>���`��q%�M�#����7"���Ȭ�	�\^rq��;,�J�蘹q�8��i_�cδ� L���	�R�3#��/�?>}a��A�M�S�w�(M�;fA=h�B����U�=SRm�g�L�6��nz�(XТ$�ˢw�'�]g�`�@���Ơ|
�>�����T��Ӻ�ş�v4�� �3}�ΚU��=��Syxt�!���IZ�6���Z�W���ې�e���O�M�����ў@�Ș�V#��R�@�3��	�3���UIuos�o�M�m*u�g����_F�$����z����^)��Y��0�.B�(�;}��CP
���]��r�Z�����F�5�8��]r~��o�;r�cH8}a�2�FZ祏��%�/�ŝ[C'e/0ɧ/�vjҮ�ܳ(��~P+l�=�A*	`��A�Φ�A,:F!�WR���7WVgQK���Τ,O:�ٗ��D�"���"󍷎�Q�8sz7���2����l�zt��k.NB�r������C,�h�㮌"t%TH�Y��~��9ڗ=�/|PP����1o������'����>�p��]��gRA��D��������I���~ƥ�HJh��L�ik��I�$M.�� ��g��;|	Cdg��y��R~�xǑ���]n�vcjD?�֤N��VZz�]3��pEstXb���~��_�u�X�)�L+ݙ�i�P�Vr)1�@}��z�3!��,h���I��w;OR�������\@���ؾ���1�Ԏ :O�k�i�a5��%�����Z.U��j[.��e��e�j&`�%����( �
�Wg�ym��'�c~�T�l����.@�na9��3Ӎ�dPtN�m���c�IZ1 e� �y�|p������RhQT��I��ӷ��)���!H4ʒS��e�v|�h�5XO�%�KS�f���wϹ�p_��@���+�,�P�ڇ�60����jP�� -o�%�Rl�vfCJ�%��e,��J-���Ie�*	�����cj��7v�� ����
����#�n�2	��(�"�2��R<ڽN��@�@��M�R��>R.wUWK�B�3I�مںx9<0׆�X$�a�bxE��K֮�H�@������ &b�}c��6�RL{��?���L�ę��Kqq������Tm}�A�`"���� ���_Xm��a���,�k�~F�8f~14������A���"�������rAZ�ޔ�����!���]�Y�����iAM��g�Y�.숤���{0�".��:
��w�����y�D=6��� j���0��4ʜ��x;�kuuؾЊq7)���,�RշL�?	T���[�S
cp�xlC:Ľ�j^i�P9������Aϳ���(���`�ۅ���/k�-4���Ŧd������֥�;��Hז�ޯ�8?s\V��s�*u�#7�R�i#������ه3�4TAa�&-����5�Ҍ�d!2�;�'�&f�V
��2K`ym�_�w6�Yxw�k�(㾑r�5�΋���I��tȗ�:Td��wu; ~��fR�[�3�;Mt�{R��6�m�"]b�|E��\r
b�� ���l��Zy��e�k��&sm�/��T{YE�ET�~>:&W}(g��PG�4�#��X���dYP�
!ւ��#d��ɟ.�0l���?(�!aYi���!P���Ѧ�La^B�;���lPqmCPl���E�k(���o��|Dh�7{a,:��r�Ί�§��h,(��:�H����P�[��@�q��Y�ug�]�5r����P�X\����_b��Ϛ� ��)�:d;���e�_L�����ڽ�wa�<nw�p��nAɿ�y������h��|�}��5H�'�?�.%�5�2_:�u��͚ݮJ�3=����0IDJ���{w�����je��K+*��u+0B���C	�-*��{��%��ݸ��(y�j�C�@��U��jhܼf�}����~g7�mx�� :��V�<Hf����#���t�C9� �`�_%OAM�GyY��k��]���BwVAsMb���@2(!3_�Y�8Z��iۓ���Pam>M9�^���'�B�1� q�hY7�K8�Cj�Fdy�#���[�vh�(T;p�L9-�G�w�_�@dVc4�|�K����8�a���sp�W�dr�V��:2j=��x�̓�a(��ֻ��w�脡��nVEIP��s�L>~��T��#���GX���]�| @�N~̲�;�9@w|�B��F;X���S�%�LIQ8���+ ��c��h��S���cl�S�u{������!��dE��~w�aI�^�\���Hk�tg�T�P<��@Au�����]]$��L᩶=��D��	\�\>����c#������Duu���5�,
��3�IU����������/�ޡ��x~.���]��7��i�>h�n�tܧc�ZGϪ�z}�z���[�(D��@$�Z7�u�\�<�E�!3��i�Զ؉R�C��)��p���ز��!J����c���.ܷ̉�><k�hD6�ص���-�W��aɲL�� �����'�\�?%cZ<��`��w}�y��I�g���'�C4��b�����#���7��֐�Z�Y��\(�I��s#{I�x�kǦwS6���}�����/����0a�쏪�$1��
*-��fD�CC�u�i{�mEeuH=PI�