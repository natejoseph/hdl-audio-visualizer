��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��W��<F�ϒI���3�ާ��$�P��+�L�-�,�86��\5�����݃nB*�I8"�d~��zT��3��ȁ�m݊O"H1���>43d����q�ܽ8Js�ޜ/�1n���c5�{�U�V�Ƹ�s��]����Ͻ�9+�T�[n�i�uv�I	F!Y�XQ�IO�?��^����@�ÙG$�o�֕f"r������p%7�Sk�78�O{�-j���nM�>R�dp��F�W@�!J��[p�(�n����%���w �2^��@�]��1*���� ��ө-ބ�if���qe��&�!J���7y�A��x���P�k�b�s�xW�d��N8��XC)�[�GF�����V�!,�_�lF�3�qd"��s��>H��!�Q�+g���7|FQۭ�P�"xHC^��(�y�\�\�m���(����g}�ڷ�����n�i�qz�1���?���a�0�V[/�W�vU������+�q��bN�����(�+�;�ܒgq9��43��UE+VN��)��p
���g���*1��>$&�����6D�*6�&+���.S�m�d�	�C7^Z�Z�~5i&�����]����c�Y���7s⯠�8z: �/�����h�,�v�o7� .X���b&=!��$�|v&Q"����IԤ�F��,~/�6��(�3.�g�
$�$S7�0�T��\ݞ���
���6߃O d�r}�L@�=�����P ��PP�%}O!&:J����,�-q������8�]�zHݧ�+Pt4��e[A��K}r���0�9]�x/<�aZ����[X�_�Y𻧉
yT���^�����G��\4�dP�nį�F���P�8��}No[�bt�ȩ#�b�s,.C��]zа)� iso�tq�GwMw�����.e��z��ATs���⍧:�^ر�<��t�: /C ���*,T�V���|��k]�a��-t��EU�8��J�bZ�3�Onoy��+��Ċ
��PY��6��]����ăvօ"�p]o˂¦���*�P���D�g1��m"�:d�6[����l�����^�=2� >�����2V��$$�`�؆M}hu1���._��٦�����m�!����e� ��8~�M�:ȗ|�����}�"*��³�M�!�Wd�֦@䶽���-.�P`'�ɠ#�$F��?� ���k'�ra�%@3�Ok�"���5M;I���&r�!��<iǏ�.��
d��PE�#�M� �-6V/-+i�d�c���ռ��6PA�ȶC��p�۽�$�9FX�gm��0V4V}>��cw֡�ʤ�P!�sW��s��l�
Ƽ�u�UC��D���ZbVu��-'�O�"W)ǔ�&Qt��?ۗ޴p����6�f�������h�8�u��`s��Y�c�a)M�l  �E5�����:s;��}��1h{i<K������yPA�{ʁ���m^�_.S�	mKq�յ7̖���s��k��V$/Rb�W�z���#p��P�.�%0���r̻FB`���"Z�XG�O��R��e�K�߈cH�@��m�{˿����?WZ�G��&X�}ݴs䮀D�����7EE�!]8�󹱺sh�[�*��Ά�h�1E �4��4�3ȯ�:˓"T������d��S��Xj�%�.��q3kxv�F��\����7��ڱKc6��"�k�WW�ۮ	h^>c�����<�� .^,)� �;k�&V˗�~&+4��Bdt�=Ǩ���itp�&��2-��+��E}���ڔ���M�9#v�	�{��p{Γ�8���x���C����e{��ר#�pц�mi��+b�Yҗ�/��_�'֮<���塃�:��U�H�{��QC��0f��B��oY�[�J���Fl�����[אַ���{{��i1�ơ��1
�g�_�~5����cU��}���{��������(M��P�E*{��Ͼ(��908�w"X䣐KB�Ÿ
k�?�IU(^����}n1��F�G��^��SB�3��DnOJXG�y��/�G��R�����M����$���%=F����<��&��_P���m�!�B��.P����;X��%�Qi|���O��ڏ;6]�n�>K��k�v��<K��,�}��bI�W
⼦P)?�T���$�&���3 y����=����F�E0�9�T��Xa�G�v�����lZ}H���-N�{��\�Iu�u���J��%���SLM$E�Ԧb+�.�/�Dj���c�:+>���{Ljӣ�f7�B��O�VQ)��]�o�&�tҵ��%_(�SZ���i&�(�O8�(#&Y�����7ʸ��	`O�{Ha	�G@���WS1u0���=���a�x2H
�#>Mܧ��^j�G�0�z/lH6y�����>�O��jT^}F�\&Aƭ��?D�i#����̻#0k�-`1tR�p�P�z�y�
�To����YF�҇����DY�s�-x���9�c�gn�Tv�=a��Y�Hv�[t����#]���w2lW��d��T©ќ_��;�r=�e/8��	$�����d4=��:���O:q��M��	@c��+�w:���(��A&v��VM��\��nz"�VxnK_k�kѫi���%W�q�bǅr.�b.&��{�NHʤ$s9(D�m�T��&?�B�!O`��w璢���Q�O�OzedU�Q-��y�hkg�J�Lx@�&��#��0������g��a�e �p���y�e[r��G)�Pt���!˽2��/Sz��p=��(��+J�����*���X�!Sh�2orڭ�-:Gl�Gl����O#�gV��5�<�b[�E�n�#q�X�� ��(�\(z�t���:��(�R��
���|������}[z�J�0�5$*1��#9>���5�5\��R���?��!tBf��!ŔPh��n��������窥�B���<�H1ۘ��%��Sw=��y�q�7A��!Wg��Aꉑ� �w�:�0��Yv�Ie����R�xΕ ��m�0~�4����r�����'Pb�Dn����R��G���B m����F�(?����/����@���ȵ~7f�=� Q��];�f��I�̋�}�Av�	��+K��r�4p!�\�rז���L >ɮ@]�M��a#7��ˍ�&r�y`�uf����#�W���
��(����ӽ�߇ɘ��2l"Z��h�����eщ�RJFIX��P*	uG�}*�$x������<�U��v��7��-��wG�}[0��� ��˚�q��E=(0��E����%"�=�gEʉ�4�G׺��/�`���7�lk����?�vn�ѳ���=*������`l�?e��/}�
 �g��o�ުiѱ��И�F1�J�+H �{�f���!Kh_�]<���_Y�L���!棄�U	l���2�Iɶ��B2�%8�]�P�O����-9W-6���tКt�lﭹ�G�?kd�*�yg"C�G=��1M��r̽ؾOL ��8Nn!���E+�gwp��~&*yk�/<��:1V�_�
}���t�1��5���j�o�u���]sR�P�`��.z��b�{�;C�C��6dQ���+�^ƚʝ�M-�]�#׌qd�T�\3�HBW��l��g���8O�k���;��a L{��N��2����%��ґ���⻞,���!^�d��!�<���̀(��M���/P��V8�}3��@]Yy/�$��Ȟܝ]�`��Λ�XP��}�S��EE��zf���q�MV�^��fs���#q[{�[B`"��^�t�uL�%9�ۉ����I�1�.� M�4�4o���%ʬ6`�7�"&b�R.�ԍ	�+zax���&�RX@K�H�g���)NsbC�>��h���'����V�
����s�DTU8�Wg�*F$T�#�Vջ�58��cPA�,�������4L9�̕
I]es�2��:MLަmq߄F�;�R��C%�.�ٍ�X�'�8n4��X����K-�jEͻ��~N�c��^?}M���4z"���!o�Ո��Y�B� ����E$�x5��F
P����˾mj�v�5������{:F��W���Gݚ2����_�Z+Y9n����F����92�)^f�Pz�{���g����%�	��,�F�b;F�6C��kD�	�]׃��J�&bu��TBV���@a���F� ��H�9fDmLx}׺7�$*��#.�Ή��u+Xk�?.:I��ᵷ/�1���t�� �PPt|�ŵ�fRw� ~�<!�X��V_.,R�> /l�e"��"����h8ȳ�~gs:n�ǮE$�)Ŷ�P�؆���Y��Ȼ���N''@�>��nЉu�|?�fYf,
E��%uv/Ț��*���<q�����̒����w6B�T\q�S�qߑk�8YC��=��A��ZP�;96�k�e�U��BP��
�?d�s ��V���*';RjSOA}z9���96���� ���[5jTh��h��9�ゴ��:���Qג�{�ic����t�ua�d�l�R�v�)@�oM��8����K��ۦ�����ם��@>�ճ��ڱ*��nۏ�yC���\WQBV�(d{ F�"�9����}���v�ϐ���Dw��C��XI���
��k�S���=t��D��ldsƠ]i��e'�����>���4F��l	̡�ḌMPy�oPP�Ԝ�s� �|K�����Z���M�mT�;��I9=U�����~��A�)�_A�:�0���KpAbD�h����z%�$�^fu'u�[�kL�)B�?��@�s9dQ�s�0�ѵ�v��#ld�M��B4�V����/��`	L����II�~��+�ģ�fD��g�i98�ݖd&���B+�^)�pl+4�F�P_�٠�����U������7F���lx�_�
�ŗȞ�]���rv��ŏ��2�����w��<����6�zʬ�A�^yD�h��{���4T!5ZHi�q?�l�^�l�i�%j��h�i  �ܲF�2��ރǕ��k��Xӽ�Ό
p{ߥ���F$֜!{#�z��.d�cu%��(���:e�[l|$/���=ߵC*�
9t���i"�#��K���6D����5�,g^�%_V����/�֠B6n�1��� M��hxِ-���@:a�8�)�"+~�3B�7�� �`x�����~� ��n�8o���p�Mܷ_��$IJ#���8�B��������y��+����P�X���6�o��.iAf�l��]Y��Rܮ��'�X}�;_����D�������f|E�+l �dכbb�'�w��]ƈg{�WS#��q	��+P_�#�R�4��6�/�N7��P�i�O�aMI��]�y�"�3�,�n�ȵĪ$�Gt	�'���ˮp��N��O�G|�_�}���a7�@�n�w��=Oy�ڱ{k��,W`�j0&QuHm]�{�D��OC`5�'	�0-{5����G&�S���t!�X9Y�BTwňS)�#�?K�KX����ܕ�z�u Z��m�D��v�]z��mwcl�#�
���[�[�ۂ8W}Bhhs`�,t~��θl{F*�����Y+�n��RPpb��#�`M�)*��u��7�6x�Ig�"޳����K���U �p̗6Q[��d/f��tfn�1�V�k"�������̋$��Mn�.t�`����eτ	�p���V"���\�L�G�3�R���y�	RHK ]�]��F��L7�z��j���7���l����ξ��'��=��#�BQ���)���׃�c}��+�{*��� ���VQ[�A|V����%�U�꒥{	~��By�����i�r�af�0 �겞�JP�H8v��p���<Tr��Cp��?�ٔ���+�"�R���(h��	���Κ1�׿x'9vc��5ѯ2"d^��� ��s�;9R�h\y�)#֞H��\���m�'�,;sqt#=�A�]}e2cg�z}� d�/����)w^����6�#g~����K Px�~A�c�U��g2
��icq���	r�EqR+�B��ޔ��}���ey�1k���%�r����a8�7��8�I=���������e�W]����X,R�d���`�D\�gW�r3Ё����Bq�%N[���$ ���c	�Jr��\o�B�<xXԖ1�}囋#vɀŭ�ľ�[�������==����pp�*/Z��hս*���KHt�.�u�|�Ӗ�������iο7�]�}{5h���Jy��-:�sc�@g?�v�����/�	�	#��z�u�����;ZOя�s_A*N��v2G~�3�c��P�#���Qg��t���\#��P�c$�n����7����l�8�j �m��*�驜�YU�}i_'v�y�%�F�]f���������~�
���@�����f�yzBCa������M�A��	��܏q��-=g.���MW��m��<�e��6O���X��rm�M���O轟T�G�^23�cثٯ�RZ�o��Y!�G�uȷ=yB�,!�N���`2r9�.���0[�ĸ��P�)��v����0�(!ܦ
����Ϗ�c�$���g&@�c�z�R���l���z����D�Ns���K�4g#����:d�59/�| żS�!�D�>[e��_����0��=��\@'�,k��	��Q�I
���B��0���]�Z*7���ԯ6{�[>��cU��
%>Z���Ap��?��K���4�����um�GkɯT�i�=nk��/#t�<��l��t>�"C4g�ʬ��JЉ�]u����B1D�BKIOv��~Ǌ�),AD����n����D�Z
�ɷ�"0z�L@���8'�>�S��po����;E$���#��5���Q׃�D��H-7׎�+�CL=�!@a)�F<�Dɋɀ/���[��ʦ��X�zj@���C�/H-���M9F���>��F�0̨���Y|N�����-������	���c��������U�J��k��Ԙ��ڸK8�I�졅^Y1�Kf��bH'L�5d&-
`cNco-��x��p��(�[m}wR8�"���8v�ꊺ\\n�	4���y�jy��x�q=V�Fl��L��7E5�r��"�����d�NX��y��)��̓+�ְ0	��S���3��`��Jϻ���0N��:i�������p��3w2�.!tZ�̪e�5�a_���YG���w_J��Jp͋�K�2�o+닾�����(��)�� ǐ�gD�Hq�R��\��e��CO�|�!�a.�����
w ��v�Бn���<^��M}�os*�*�S\����R�!�T�N���㟈r���+��D+�Gn�v�6Z�Ɋ�l��ݝT��h�@2�9]��R&����3����D�(��8����YS��6:(�^[(]Ajc���َﱅ���²8��^E��J��X�����SUd�$k�c7��T�/�_?/�ř��vf�$���ӒS4���~䣚]�t���W�ٝ2���ጤ#ìOҳK;��!��L��S�@�`�A]'��|2����A�Q�K.�F���Qbz ���z>l�Ƚ�i���B�L�bW4����ϋ�n�;v���PP?��u���V� �)�GHj5��v�K�}DP�"� i���7�!��7ӪlR�c��E��1�$Db��(^���
