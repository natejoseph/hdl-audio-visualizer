��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��=HAW��-F���m�]������6~p���nV�#����@W��]B��̂QH;��W�̥��E�B#H�b�_�0�B�f�c!� bo܏����7(��;�}�.�@�Gȣ`��Д����>ꡋ�+������l���>8������o-Yv�Z3�����{���/�xۭ�Q�!��ٲ����wPc0�<���&�x>+�P��^G��qFtB<u���.�����u9in!������)G8Խ��	�,���E��o�矖���� ��]����%Z��������)���핬`��S�n9 �Z>�(N�u:]���{���ߥ�l���3�G�]���I]zM�j����,�p��*�- �	�(����OY0� �iexm6%��ӬQ]��f�{��h%�Y-���P�3#�[YM�eN4Y��(�[�F4�� �oga<�+Ŀg��z���K�N_��J��	!���������JyW>��*_ ���V����̈�W�07>����߼>����&
%(�M�zbL��Z E���^�Oz�ݯ������C��C�r]=���o��K�K�A�J�G���_F����ea���j��2g��Q�'�W�|��y��α��+˩��3l����5��RI�@01�ŏ�kk���WK��`>�%N!Y��A���K��[e�P�'[��.A �R��oW�D��i��,�C������7p?�ufX]ʌ(\9\�G��K� nf�]���X�Xfh�$�R�� �6�U671.����7�{� �(4�Z�ꁎ��X��d�����k�Fp)��]u�[BݮE�8�E��\�/���1�b��7N�7�.��h��{�2(eQ~oКJ�$����H���4�O�U�֛���Y&Ȇ��$���\����[�m1ޱ?�ð��ڔM42F��	c��h%���ߨ]G+�wGrg֎s5X8i�-������>�"��]�� 	Q��+ٖy����{�.�ڤ��(E:���a�78̥ 4"ϗ��GT�]$���p�U�$���� �%�e���SŠ�c;�@�F5�|���3���A�YՈz�r�G(e]�h�P�fV$ݓ;;P)94��������[ݺ�V�@4�}͈N ύa:�֞��L�qBR1dh��kYTC�w��M3��x�\���_���������T65f��i�l"OK~{�[�cG����¬�ckG�xSfO�>`�;�4}���A�F`s�K}��8qn#I����._q@�F
>��u/q%Nx3��VRu����Z'��� ��I�_I)!]��"���Ð����;��[V��q������p�V<9;��6�Vٰ�z��:�j����u4F���)�.>$���'+�H��IZ�Sڱ ��ӕ��� D�)���q�Qn/ݐ�|�z�.L�Sok?�̈�@2G��H�E����ad�/���t�c��d/BB�3?�Ɖչ83�
P��U�����$>�o�
�1(官�� v�O��`6�/:*o:ʇuڨY ӄ�"=�.���#��'FRʐ�o9&��MF�;s�:��Ց��S�~�~��<\I�3���e�`�B�9 �5W�m����"���R�ۆ�oy�d�����W�X4B�u���t�ew�p��I�������`�y!	[��Ҡ)X���uL�ov��?ib�GY��"�R�l�"X�o&(fDS>#vV/K�j,��k[dV/<����Ǆk�~==5|�θ���[��Ic,�>����R@�@� �Ԅ���{��J��ӺR�l/$�0X6�K��WX]yXQ�5{�d�Ȑh�W��.6w�ۀ�XV���:�lT8tG���v�����/\@�w�]����4N�l]6T���p�X6��vBξ�ќ��3��a�b��N	��*J�$��/Q"��]�ڨ���P�$6r���<O�!��P�'ӽW� ������KH^�_,{k?�x��9�A9��3yǸ6����ݾ����W}B�-_p��M����-��žҪ'B��¶e��;f��
4�r4�.�f�_�Q���7u�G��ģ���B���!.��mߵ��h.�(@e�/�U�;���6�s�x��)i�vqJ�"Z�2����̫
_����`�[�fwjDt��e�R�5qFT��"NNm�a�
Hl�j'㪖@#�a�P��4!�߀:� j�9ׯI��D��M)V����ݼ�o��˂5B{o��C�þ~�b<�!R�\���ٷK�`�Y��	�W-��@+�����ЦNi}U?}$�R-b�D��\�N�xuf���h���C��S��w6�1���Lo�k@�����c}�J���#�n�ٔ�6���>�����&C����M��O$�����TX�g�p��Y�U�>#�zJ��<5gr;�9i����í2���2�P�7��,��Ж��v���LK���y��?»o�w*���X文yw�Z������|bŏ�S_���\x���B�9ހ�?ĉ�ޮ�|78L�q���h��n��+t#�=p��6Q$s{�S����f,��L�m�*/>�C�����,�u�\00����<�R�-�nsIp�X�>��b���)�N?~	��u������F�/�}�Zr��i�qE���T�!󩊳|/7���g<S�󇈝/*��c_k"-~W閭{N{�9�庀����\�Ǭ����3(��R�[=���a@�)!2l^���-���?1�����|��(�d)=⣖{��c�M+dp9��=�d!J����v�8��K	k�4�e�a̜�hi�����Y���c�O$���W�I�e{��`K�!Qp����aS�!�ْ���Oާ����k1o�X��g�Ӑ���� c�QK�:�j=��%#�s�u���Ŧ`:��������V�Ivj���'Iص���q��294��>M h��x�5�V�)%A���U�����k�,dM^�����z�Q��8�A�'W�a�9���(��31q��NS�-QC��?*���)��q(g���,T���9�'^�4�f@����/�a��>���2iƛh�*�/�C�b.�����X�;j�^P�ݴ��Q�ļ\^�PS��L/Gc��Z�D'�t[�o�Z:�\��-5����k�rC�[g��h�*/�m</��?'*�D-EVV�V,��8r��Vp �}� ��P�A����'Ӥ�=�>��v��s���U'���Mc_K3vsf���SKrJ<���S�3{#�7Y�DC���!�n�=��i��L�L��"x��\Q����(����؝�D^ �\'�E�[]m*��iN�M��OW�������9��P�D?dͱx�m7e�?���3y�<����f��΅���Ɠ$c�8޽\%-����5�6{u����3�ӈc�6Abk�mC����c6�����A��o%'�=�1rl��)z0P<����G�=`���˰���پ�i�Ӓ�A2�P/�A�l0 �]*���ߢ��1���Q�R�*~ )�E��d�H�y�� d.�i�G^}h(J`E�3��k�4��K\]��ڙ��zH'T�,�F?BmE��!�)Zk��$W�%߿��j��Y$����(��M�x�N���@`��^W�M@�ۻ(R�L�2F������1>Ցj&b>�e�/�D�v��q� ��]���~vQ?#���)��{4V��<���&'&n���
E�/cǌI�ܚ��cG;Yy���\Ԩ���%�_σ�������Ya6ڲʜ4v�l�3O��#
?{Y��\��}?\��9�M~� :|熨�=nE����k
��ݿS�1; ��.����\ͣͧ� a��~���I�-U�H�č����q���W"7�6���Ǌe�l�C.�r�H�o=2��wu�����h&NKf�as��߈G�8ǽ�W�P�bf���g�?������I��&G�3��������::O7���-��]��U�!�+l|���ѫ�5�u�w���F�=�:��p��T$I뵬Uk�˹Q�#����y�۟�n2���l9׎�����A�D�Z�� x.J�B��T�#����p��c�rI�ɗ�g�q�L��0�^�)�4�3�ܪ��'P\a��P�g�!Ͳ$�W�N�^�\ޗ1� ��Y>/\�������gFj��՝�wKp�H=�4�ՠ=x�Q�������h����f�[�C�#Ɗ�<�n�g��G:;X9Uͧ8��d)5�nX���j�Q{v��PK0��2���\���Z��}���RI�Ax�������.�A��2SCs~6!̚A��K�'��Q����	 ǳ��Bg܁�S�iuB���!Y��t�8Q&?e���T����.7r4�@�%Q(֌� v��(���G�#���N+��Ůn���C��Kض�U��3j,U���x !%=X��&�TÃ�q.�n ����x��OR�dsT�}(��Ih1٪��X)��/�7/���Э2��#徤�w��Lk�}��\߸�#8�"�Zz�e�u�P0KMU�:M1���$>	��e��x�m��u�8*5�io\�����T�?U#͢�j��|���ȫ ��@XKKV�`�`��O�𱔃w�z2��<���φՕ�̯��fM���8g��Pq� ���[o��"�S�$	-�� ��W-��`�,�<�JI� ��d�	᫆��v��eP�hP�d]u��_�'���\�0uK` N��(Z�Z��h��HQrٍ�����<(o��������$v�o�=�=�5n���������[���3-z��dI7���������Q ��]�R����XOO��������F癸���cײ1>h<}m[�����Z�Ѱz9���l����:-�q���գd��
�& EWpO��������@q��K���'���	IR[��0�9A�2 �^S��~���1��P~�s;p�ύu�JĬMGq� a�����m�T#�[�lK�b����&�U�k��!�m��8N�+�_,�48 T4n*�{���LA��:�~C�u�m�Te':4�b�)j`c�LP�#��G)s*A��E�֮���#���Tp����0�ݾx���u�)>�������!�S�����nc��O�ʖ��x���xV���s���W�3Hz��sb������<3�ˋn!