��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�����3ܴ�U����I=\�m�q!vx�w����[o��%`8�p��6���=e�_�5W�뒄Io�SՒ�!`����w�����-B������'M�1�|��DH�]�Z���|��w�����2lQ!hb���L,%�p�r�bF�ΈY
����3(���a�Ѣ��������GF�^ň��(@}W����Xbo���x1�g|W}�r�8k��`�"����J���zn��R�C&}�[����]x#�̍��m6on�{�϶'ʡ�ak����@g� x�}�s���q}w��k��Q,���rb���<������wE�wJÝ.��&���-	% ��-A0�	Qt�r���S|�d��H�l�<��!�'�`s=���Dn�$��a��mu5�?�s�at�
�٨�P�j�\��������3 ��ܛV$	�g��vW�����nnn�)�� �s��:b������R��4N��l��o�u�]����l���PI�m3.�v[P��簗�
E6�ر7ee�9S�aM�L*S��c!l-{���SJ��r��W��fOi�*8s[�����x8`h�l�ҫ��%��-�9���db�ml�yf޵�����Y`�W�l�3�PS������2f�#ת@fض֥�	�DV���r�~�0���`�����m��2D�)*3��4�.ރ���V�>��=rt���Z��De��J$c�ŀ^=}��J�%!������4p�̇4�Z�F� �k��$K.��k��Pove�JѦo���X�龍$���V#�������p�3Bm
@���Y����	t�]� ͢�Y�E�V�[���ƛ�j��>C��n
@S��ue'�m������2T����~���p��t ���J7�<*�R[DRiwY�����ǻh�u*����u+�1��i}R�pr�0�e*����Î�Ub@>�$��9ǋ��E/�p_�� R�N�Ӓ�ȓ����d��j�uhϩ�Y�k�8�<k7L�ް�ph뎕��c�|�:�=O���>_&�(iO�q�p3	���S���+�q�a[I�̢�Ya�,d�3��R�ė��=-y�B����Y���e����R��n�����߇����<��f^�J�2)�G�JV�rDc�Pmc��%k1��6nK��^� �ɹU�+Vx�uH���� 5c���i��7l������F�K�Z�"��T�Q���i�U� ���o�i~`P#ǵ�����#�7�A��[����.������b)
}_Tv}��`;�޻%Q՜c�#��.�I��R�)��<���e1@��d��ɝ�ޖ��ށ�����G1QZU�7�HV�"��
����[����D?ux� ��A��Q_Z�Sp�>����@�X�7�CuX_jy����Ӛ~KҔ�ڇ��{��"뎨�4�x�,M}!�[�-	�b3W��o��$�J�<�t�R�A)��H��9'�k|���D-�N�$�OS�PS��u�Օ]S)��:�2��2��9`�L��Rcy}�9d�n�lG�P�'�6�b�\����8
jY����(�\O��xE�>�'�'���}�fȾ]��TNڛ�J!�9�h}ww��H O�XQj�^8�*��s��-�@��Ƕ҃\-fakM/d�I�E��Ψ#P��я"��N�����!����/�7$�̰��ʕ��)�$�=uC镙�G�.����V:�W��35�$S� 9�}����0���ԢG���պB<W&��+b`���#I)"M��1����/0o������\A'Ѣn�܏s�MS�v�zZ@��d�s^��+Q�&L!����Zz�c�珕p8�Ip!OX�X��F�v�5��G@�W�F����br�^�\	R�-<{U�sg2���Es`�J���r�+���3�PΤ��$�| ��i|�:D&�R��0e�)/�a*~r� CD:���h�ݚ:�AW�κ�Z;�����(.�`y��M�֪M��d[U~΢:o�7�$g�V��V0t�5-	�򰼟m���j,0����=�t��%:�^"̶���N2�hh�Y��W8,�]L3�p�E���a���S���&7���"���yI��$_��s��h��c���<Q����'g_��;��W��=�{�+Θ�3���%3O�8���2�vO ��% OJdS-�7f��O_Kr �UMn8�WY%;�d�*�)�I���
r��xA�Ԧ�ډ<f���Y��tρ7��@��뼿���ؑ?fn�y���+��� Ț�%ڌ3���)����������:r7�=�)y������H�*,e��B��NI�(쉜$�Y8�������
ʜ@����,�I֤V���&����%�x��Cގfm�4��j<&��]�\^6�M���*NW�Rq�5�u_���K�A�k�ʣ|��x\�r�앙����,oB�>��Y9%k���o���	�<>�T:�1��?N=�S��A��d���ɟ�~�\1��0�l�h��?��&�g����wB�C�eM��n@½Vs��Mŉt�#t��f�܀�(�%ݗ���<�$�$�h�9�ٰ؀ߴ6�A��E�"|	vO�,?�&Ѵ1vd���\�~�-\U>��o����7���ѱzi�^3<e�d���	+-�B��p���؋X��լ�2���4)mT�����1����ֻ�(l����nW����)��@M�T�%s?t/�ՂOY2豣HIת!c�B�P��XN?w�m㸎��u���u_r���F/v5��ģ�=�v�%OW��6�
 ��%Q~缪�� &��&>r�� h��h,4R�(w ��.V�y܈z�v�hv�����<�y��u}�PS�B`�R]v������o�<���/U Y?�v.0L�TM*�$'��~X
 �����͡��)���bn/�c��]�}K���Gy�:j`i���T�gq�H�պ�����.��j,�G��@�O��Y��PŚ[r�O���VN�����=�C��Z0�Ռ���ϲ��a���Y���_J4�|��������3E������q�HHB*��B��&�����/"�;� v���{��������v �E���m�,�]���?B���͙�Zzd�!�5�߿��#͑��.Ok��Wٶ����(��#�Ss�[��Uw�I5�#z̔�� Hd芪*չ���Xm^�|I�
LI6��$��l��V��x遲^��^v�eec�|�kTX��R��mST|����(L5�s�x��sr��ʣ32s�XE�t� ��?q�5�3=�5ߑ9
�d^-g���^#�[�*0]��_[;���@�Rl/�Qŷ���̗���V%�T���D�G�@_T���^�i%T�V:��`Y�f|�ڨ��ᨇ1�z������
ܠ��w ���ݑDffǝN�|v�W�xs���.ۡ7�v�	�v9������s$�wè�:82��qo]	��
z'�I���,���D�����&S4���/���������rB�_����rlJӑ��E-0�s���Q����J-�+��<e5ݮ?U���K���U^#x�Ej����E+��C5et�eӍȸ|.�n����R�<��\�GP��,`%�'�#]�@6�@Dv(y��<36��ZZ3��;.�7-��Nj�=(R�11`����� �%G˴ћ*��-��
�d�"��f� V���+8e�;e�˱-s
��#����85I�N˭�#=�f��O�:z��g�/?�~k��b�=j�o�x%���Z�:-���Ҙ9�8g��J������xh�~x Eb��R�?�Mq+2��Y��܊�Kbi�a��JԶ�n�⪔��K��n�*�l|k�,��[uM�T]^sz���/B�O��C�E���4���挧�Ğ���9Y�C ��ȣ�*���%Y��R"�G���>�k�*-�m6[:��x�����&�3��f�d�,�u�)B������r���:a����P_�=�d͸���6� ^[��=D�����|"������k�ޟ�r��#d��}�������#d��9��pZ�}�+kb��\4f�*g�[w�"�R�j�
ʲؘq����5�᳥Y�A6�~�	6{���CS�j<Bgm뾷;��6LQ�'B�Q�7�?�-C�²��q���E<a�:u0�}e���<�����%_�B=+�WG�ښU#{��N�������5���Q�x���6��7�'
$]#A��|�s�OC����1�(KoD�æ<�d�����G�do����`�S�i	GV-!en��/2����Z^KRG+�۶��]̂��NNl�5y����!�1�L@ؔ���{�9m�>R�r��Y]�z�)8�Y[�*`��i�����r�k�N<47���A�Q�S&��y&�»<\�W��C�`����o�[Jϱ�G�6�i��ѽ���o	b�0<�R"�,U�m�]f(�����v�{��~)�����t���l`�` ��nj�œ����opR�{q�x�@O<Z[0�6H�^e�x#�+@�j��5��S��LhP8��@u�l3I��g>�� j0&\<���7�ϫ�V~��f�'^6Tg��%,�Y��$�u�<����,c�T�eN[vH�v�ÿ�d?M��n�mtњ3;	�Zߜ�1�K�������_$6Z�H�c�*�*���8��U\ؼ�nӹ3��;�Q���b%�ٞ����ql������tt�*~kCdkd'�Y>k	#����oW���y�Y�*D�u� ���K��.�����*�_�ʃq���f��:����5 �g���88�f@�.p@o<g_�ں����u�vb�I�x�C]G\�!YNk�&�Βu��%� ���exîq�U=�cU+����S�]�6C.�K���#��6�.rP; H�G�B@��Vw��~�����F�I���R� >�=����I�s��2�5�9��R䝝:��jK������O���C�g̽gPw�ztE�2��8�c wj�f����w 9����Mˋ�	]�!v�*SR����1�y8Gj	�ƜR����ʣ��)3RE�A�F_��w�����3��~Ҁ�{[��!"ܨ�^� ������{b���"љ�ݗ&�= �S$ӽ�i��ѧ��"s[�?x>��[!�%�0��>��z��G�&^�([J]N�"���r���O��dw���z�ͱ(uC�+(S톿?�r)�v`	�`�V��z����<v�gI�*�c�p��v�a��/��
"�?��?�ϭ�������L8�)��M�=�q{կD<
^��h�O���p�W���Z����p�W���Tm��}�H�g������ed���X�ܝ;�$��g�N�m�@*� uꅸ^a.S������f��X��V�8E�q��������a�q�Ե���V��@���q��C�%=Yy�5{,���ma��ϊ�Ρ��9z��#S�KZO�m��	��E��z<�D�����I�-؝]7 繢���u�G!Q��A ٪��W_<ɰ	��;g�H���o�Wtt�)�q�'����.$S�P�U��ˍ3��  �zm'�U����X7Z'H(T�&?�~��îZP�^������$�X�z�6ZsO%#�V4|�P�\>��/�`��g#�O�v��y��ݾ���)^p�B�_u׀��{�Q=�W�P����O�v��ku���CΪB������fb!�y+_[��������;ř��mo�\T0��� Hi㙈 ���E&e "qV�?d�;���>�Q�`�Q��L�#Z*�_B~��*��	��d�o��)�&�	���96[d���<QKH��nS�A��3(5)�"��ye�T�f̺=^~�\�,T���������z�}@��PCJ�#��]�r��Gi�Q�l��Pavg�)d�Cm�7P :�:Y�;'��޴<0��{�YI�#qR���ࢶܫ^��	����ŕ�� ��rwn��m�;A���ǜ��9�z����	G;�D@��gn�*�z�����&�j�� ����m�_����F�/	����&଄vܔ���ŏ�Z'�r˶#AFѿ(��B��ܸȶx��pZ��<Ԃz�7�Lf5	6Kt��;[$ג��/C�5i-��L)��M��6�Y�kQs�o�F����kt!Q����胓?�'X�?�s|_C���xt�����x)cH�s�����'2��Ǒ��މ�4"��Ӆ@�)޾�v�*�QU
�-���9��mF�q*%�~u�!����v������%~���Ģ�HZ٘��"�(C�r�ߠWz�X��FL�e��#�)=�m���v�y��,����'�G�z�� ߞ3x���";�7@!H�Q=~$�N� }{�y�ưCg�/c�'�Nzω���wMpa?�����7����>��n�釪U���Bԡ��UB9~�H!��D�<K=u��h��3N5����-Sp � 4i���,�"o��v6T���1���%���Hro3L�K��Ŕ/{��A����>w���P����P�@��B��8����x�3���,m/�X �hK�"i� f�ěU�NۀqE���A��ڍ-k��S��c��2��+�j�{6���Z��2^�|��T�5��H0��IlД��_^�y��Fk�O�X�.+�gw9fj���"v[k�%���c[�?��f�kd��w�A$~�L���!�(���AJ����a�R~��g���X��HE��L��Q7����I��s$�5��E9Yۍ+@�W�=��1T�C��X}�a��]H]:�W�S��L�>T�U���i�W��}ۖl��	�����7�����T%�V��Z`/|C�A�
d���"��2�؏P	��N�`�)�.�Z+:�O;�����3i�V���G���VH<���'l�KG�inj�dHMK��Mc~A[_�U`UK$�aҁ�۟���V��x��U�O9�=l~����@�U�=��A'��XٵH�R�`���nW۪8ļ�w��t���3y��y��P������n���������l���a��jM�r�9c���[�d����]�Ey�m̦�Ū�]O��W��IH�Z:eeiP3����ҕ�NF����kuBI ԤL��źQư�c���#��o!����|���w��U��O�mUFڢs!|]}�r@���]d*"����1��n�Mw��`~[H-�h2AG��&d���gҫ�T��������]�S0��R���>׼b�H�>���3J}��t������L&��~2����rm�z�������ݿ���Z�S��R��ٴ}Y��	D�Q�J����3��mIS�����@?��CC��-Q��5�>�-[.�Z\C�W�Zn�e�^eW�e��G��@��}��L���1�H�P�ڣk�.)�
��uY\>�M�����<���:�7�џH��D�(K�YZs+%����X"A�V]*��̄�
��Sz[%������˩�)�鋓����ո�+?�k܌|��
2_����̥ZȒ?u�-Or�[8�P��g@��UC���o���$�P�Q
�����s��KK��qG�>UФq]-�3�6����9� ���߂$�K��Y�J��9�C�&|�U���Bgz����!\z#�ʼ����j^���-�3�-��}N9F`Z�����Ѝ�ʊ鰐������9���L%�8��H1!-������X$s��ǶQkw�1�Mc���1`4�s�	�|6���E4݀���ud����/�ڲ�Ε�a��X�h��y�5�S�#��:(�J���W��3�c�/�W�y������o�������\�o�M�:xgq�2�3�M�m1J���?�|�_NhTWj�)���;Ņ1��EJj���䩟_�%
q��wn����@����p�X�7g��?���Ewo�FZFFF�U`D�|�:���i��Ɖ��;瓒8�	�G���{��|�Z;	81���y�-�"�O�yf����Y#��>1sjgS�/��3v1P��Ϗ}Ud���ȎMv>^���N*J?�W�	��#�N�!n�(��[����6���o����H�K	VI�� �b���G�iţ�vy�c�A�76�O���hN'���q*�&��ؿvZ� ��&P'�DE`P{�����(3d�:C48�-�J�,�r;<O඙������nd������⡄��넽E��̗��-�y~�n��>�?m�AB�k_�\:0?�z�yY�D��AjS}����*�~cn�_��^���ލ@�c���.obK-p��@F�m�>����j���,�2A6��$�|��u���}�r"c��z��_^��OD�c.�E�@�5����b��L�����@>����#�r�Sz�I�W��҄į&�4_�� �z>�a̜LW���	�~�W�j%�hp�wXW�Me������1�5 W&hk%f*W<dVUTƅ������̵,v��|B�Ċ"���^oJn]di�n�lU����	�.� �7Y*p��a�ZaB��`�þ��'�"�o.���%H�^aS�q�����y��7m�dٕ�u��Sv[�=�Uz���{Zt@��OÏx�c�R��ͬ�9�D�`׈ےW����O'��OXaP��{dU#l֐S�Jy^W����O� �բ��,x�>hKU��j���bq�L/�F5�e���.9g����[�؞�׿���,����� �>�ua۵�'RS��HtLY��y8~ߑ˧g�%�<���w\Q�+���`�y�#v*A��O���7��X�"<U(���l� ~��)�ع/�%��'��/�Vf��]�(��!�ZF�[J�[f����^^.r���O$U��y�Ɋ&���ɝL}��g�����9YN������%8z�"�����BQ��t��oq*�`{�/�Y=q\D^m6d�T_U��8���I_���51�C��޷=�H�Ԍ�6�&G�=����$�����=?qŝ�$�έy��T�ub�xOE,�k�f�|kE�5U����Z�-��i���0�;��
Eņ��x "��L6&��
�:�_3��4������x��T� ���ecy�q�z�y����� �7���g/��#�(�ZƦjxb����kz?����7J��D�z��I[\�*$��oS�J1�N�/F��#��J0�2R�����w����� 路�Z!^���q!(cĢ��c@'�E�Z]����շ& uti+���� ���G;��
$�f��WJ�;rtv����K��ib�ͬt3��)b�����9��d%3� =���pg�Yk�Wz7T��BOͫP��g����X�ϲ�kXu0�SEM���D̠M��N46���L?׮�7���yP'�X���`4ڪ���ЧV�Ĕ��(����O����+2�|*��J���ރ�+�f��\v=�[N�;Y���K�"���-��W����`ߙ��2Z�L�'�>�个B^���|�$' ���=������EJI�����a���[ lM9������{v���C����wp�Wo�l�������������O�n�\�nF��lB˰�L���	IbT�Ҟ̤؊�f�}0�ey�}q�Y
q8��]ș��Q�������O2��YC8���]\M=���S�D��I.�u��
;4�B/u)N╮���i����:��x��2&צq͝+���g�{�"��ʚ��`��G����x�����y=U�&��`[(�²�i��8m�)�G�J�A�;�꛿�;ƞ�l3�/`�o@T�1�kHf�k��/ʷ'��9s��`evP��60�uA�:�~v��Mո�m�M��I�#v@�����S㸯-��Ga	k���F�P���B8m3,2�J 3���~3����u$o�H���-X0����������ð���?S����
\u�<�(x�Ε5�7�/�T��2��tS)��-qF�cM�B��Y�9o��fSK�?�:�;l�ۑ��d4a�(�r�?G�}k�y|Uض��n�YH�p`��]3\�9 q�ˑ>ex�en}��20;X�+S�Sg`+�R��:	B�ᓁ�!�n�!�dm�WꥥA��FN�FU�=f��!�k�9v��+��Tw}G���׾()v����bg�s�u��O�)�ۡ��@�T,�1����0��F�ĳcX�������ka���&����n��Ll77M�#����[�i)�`��]1�d";0@i	�	7Bg��]�@������cf��O�8+��.�-,&J���`s���C�K*ZG�9)#�aZ�YO�9���&Z2���̗k���QNE@!��`�	�+f4�h��贬CC��%rm�pB\HG�Ŵ���)���s��/b���wX��4{���[�+�����kb>k����#`f��jC����P�<��ˉ�C3��CN��+�;Ӱ|[�0f�6�uT?�� �D�0��|��3e����q�m_�iT��'e�ԧ�R��g�J:�&���걥q��e\:}K�[�y�\Ő��
�!�^38獦]&~{��>dt��A 
��i(({�0�K�|�Ǡ���#L���ґ�h{�d=�E���q>���J���
)�?�5�<�-���]�S	Ā�g�S/��(N���&SХ�F�9�F���?r�~�����.�wCJ���]@f�P!���M� K�l���悔~�*��gDv�a�P~~�\�#`f��ꢼ��mD+ �����[6�Z7��Ĵ��ni��$��H|�#mW���$�]�����/�"��}��L������i�#���,�@�E7�R���b����q��Cψ�l�m�]Swg�>�S�WO�,�d_2�c
��sY�e�o|�k�c