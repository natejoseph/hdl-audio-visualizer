��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��Td��dxC��!k�h,�_�p �]�¤���M��<���BJR~	��FdcB�t�J_�7R�x���F��a��ƪ�~��C9 D���˕VF�H��f��n��(f�Ek���o��"� �&"3=��*��B
y\��3�vC̟>uF��X?JR�����ҍ?	s=E���"k��"L=�����	�,U�vb�F��q�h%썖d7��C�i$s�������u�I^דJ ��+��S�q��
���].'T�h�zw~`��}/�l�B9N�4���Ȑ�?���Rb��$�b���R	�y�P��^�D�3}�=�R���qA�-wMh�#G��,�� ��^�{f���v�x^^�az=�m=���"X�{��E�Ԧw��DPx�޲k�K䄗J�����Uѩ)�LT��N�>��Xpk{��FQ)���DI�a�����)8�/�\����,���$�{�Y3xS�fh���iH�G��A[Hg'UH�}����ȼux<]�-�xU*Q�#^�Q�g��
�L��8�p�/)��w
����;R#�"�kd���'�*����T�0Q�i��Я~�����jTK'���k���5�������,o��Q�!�ֳUzsD��D4�q(��l�Air&H�5�H�w�����&$��?��+A%���Rva	[%q\~�?���������+� ���0c�iu����ﴑ��bR1l-le���[8�N��L�*�|�O��`#�u���8c��:L�TP�ٯ�ܓr�Rn�N�xI�M�D ��e���he�{?}*�I�p��n��9��)��l��v����2��9��>��lH�Z��6rrk5#������e̉vg��L=i��ws��C�-����%�-|9���1�m�Lբ[��,��%B&�k:U��҅�'&x�!��0u�Ug�n�NI ����b
o9[is� ��'�=���
6��b2[�(�*v6�Go=1U������ٻ5���\qAN�c��b8�gqx���SG9��r��9�b�}�o���=+(�PߒU���)���
&�tb&�����Z��/4HXdU�)*��6���g��@n�v�����`d�œu\%���N�QlGZ����*=Jsh$�Ճ��1o��W*��{�(�R*Ty����Դ!�S��*��{�%�۵#������Hq�0¦d0�E�@�8Bѱ8&ϓ0`�SRx��@�R���p 5���q{O����E3�`�C�K�V(��)��^4���9�3H|JN��K��Ny�h���w�y��[���݊o[q��i\��o��-=԰�	XTmq�óFD�E-וuo �Z������E'a0[�������W�Ҽ}Eon2-	V9�<:�tsP�2lv�@ϓzM��v��b�Ҥb~ºcnF���i�`��_�����kp�_�J��(\�<�݂��鴇fA�l`��|���\���6.]?�-|�I���
`Ɍ9{�DYp��xwA)�j��}o \	{����
�o��Kt���
+�L$���ɫ�[jG����V�����$��NB�n�6��t@6��#Uˈ6�P�!�$'g�T�)�d����k�1���rD�QI�+���]��&'��
�X���Uuv"�I�+��6�3GY���Y��0��6��qC98w!G��2ͤ�C��]؜dKz������yh��?w��dV�i%�'�5��j��B��H��x7e`kІ���Z�c��X:Y�1WZ�����%�7���"(9�E�ꋐ\y�s�	Ŵ�=ptګE�r �[~�����R\kHw�`���U��K�����y�5�����#"�7����o֊���Fs��j�Zם��xW��Qo_8����� �նS\�6a�=����R��@Fi.,�j�B-Į?Y�|��!Y/o��1�tk-�N���f;��btB7��l(\aH���g��Dx�����?tj'�Yh��r��{���O�|��&��*x�hn����J���rǡ��G&͗���㋪6{m���=�iOVՐ�3V��!�/�6��k�$�q�U?ݒnw� �sc6i�p��V^A��b�Ws����Z
d��{B :{��"�<v^J�����+�f8���`y`Rp6�1���76|��p�+`�����˪��nR�^����lV)��D�s�5�\�YM�mqޔN$ۗ�m>ȝOԫ����h���K6�8��F�7Oc3��~�@�Md����Gk�݂n���e̩��i �[��̋��a�~u��@&�O����������E��oԣ�גo恣b�3QH<�"�7��tTk�Sdh;f���WQ΋-`Dp^`�&v�������E�	�;hs)e+��y?7�����]N�H�}	9�(%��n謫`�>[Q�FIe D�ʆںƮދ���rS�� �rƛ�ŭ�ʺ-?���d��#�$T��%Sc���i��ӑB:=�nA��d���l���dhM�lWB���Ih�oh�ܼn��9l/<��o�{��4׏�Na|r>T���'�:��}]�� 9�!�j���}A4�K7�(��?�o7z~j�֓�D�x���`��K�5��'k�(Ǉ3�g��wLd�����:U�2����6�'�fp����t�M���N�P��**��km���J�b (�z^�
��;�N�t��{�"�� ��AW�I9����1*>*~F�p�,ȟz�C��]�}�EjK�y@�d����T��a͵`���@㓱��p|��^V`bG���B�w�x��@d6�h���h?� V\��Z�c�B�4�x���1��x'�:�?��I�HA7�;�y�S�"E����dL�5��.D�N�1�7��z�*�H���_�L�I�����`~ >@���NX�����m����L}�4N$�/���6�9{*J�f��ἑ��rtk.���G�[~�bt�5��Rh�U5�e-��Ouo6B1u���h��`�4�b��>�O΋��][9��m��5r�t�qb��°%Ow[���Ն�;ɔy�oˎ��zmgu!�+Ц�8�T@x����	7��~�>�K������aNgY�Qz�o�ɗ������K�F��GF~�y��(���JI�c�g|��($i�ߣ֢���v٫��ޘKRs��s�o���V�Oe��+)�@yr��D�����-�q*�I�Ѱy�6��;��Q:����)���$��em�Y��6Oc�RZ �ؠ��ȏ  _ݮ���t@|h�Ϙ��~���;��5���gMܤ��*eZH� �E��`0'�En5
(hR�e�ɰx��)� N1vQ�7Z�Q��sN'�=5iǬ�<�g���^��?k\3��FUdF3�A!���z�����C8�Y�vN���A��ä��3�M����@�Ӥ�-~�eKZ����8�O�������Ү����ѩ�py�?�@�ű��F�G����ħ-����B(�1]�	v���C�gX���s�WS�T�۴�gw�nl��+{�(����!*�O���'w�sA�na���Vψ9��e0<��vQ�&N� uOQ���M=ъJ�_����1�*?��t�����X�7������`�[���0��R�>1�G�p���HR��Sv|�.gVT앾�m������wcv���z�f�fb:n��,?�T��\�%x�UĻ�+k!k�Fi�Ć���>\��i�pE3[�ü�A-�a�U<�q��9�/�Q?�i�/���?���[���H=�[b1J��+�y�D�9]��.�-�-$����@�z{]F�!&c������픏�T)˻#V�"z_kW�h��Z�#N�2~�k���ګ	�֚^��cq�A�7՝Vd�M#t�-~����2��6F)!�H��F�Q'�P3����d��B����6��gޕ-:`��p!�Z��OY�
�5Vc���-��{{�qmG2(�&�.SQQy�J�����N͗�١��8��H�7]%�3�NA~d�!�٨4��Tap��G��I%1�E$�D��F�	ccn�ڨn�����ɲ�Yx�7�2�yM@yib��R�h^x����WQ#q�5r�7�AϚ�؀���3DCt�$f��ǹsN�1����-�&r�"�f�[m�Q	�όd����5_ W�ߒX�U�o�����Q�(f��<>�P����9u�ڦ�g���Iw��V7��Zf��{�������m8����#���(x��'zi�r5��;[5�M�LþA���8_�6uQ���v��M1����إ���(S;}�Dd�\�'o^��p1�q��
~1:�8��R^���y���7�A��"Ϟ?�Cd־��мA�}mB��H���T�l�63+�h7A:��c�/P�&E:�����A.���T	<��zi���=���>��~���+�2n���"��������¶�k�3�ܽ��|D ���W��5�	3�644�D	خ[��fo�d�:+m����'����ͽ����BJ;{ځ���d�Ō��P)ʳ\j���hA��N'�p疗iR�=�`#~Y1��gv������{��}�NK���Y���P^�l��[���ޭí�8�� F���z^�(����xpҖ�eK�#Hk�l8�Љ�S�(O���Z�A�����lޤuJ6.O{�c�]d.3O?�R�N�u)�{�Qcj4*)]H�=�����x�fB]aV�K�?X�$> 0�����e��x��ݙ��X����B�^F8��ݴ��^zC��g��E��4�.�8����m uo	d���6�r�G��Rg����(�".��&��s�� ��ơ�NaF�J{�r��O5��O3�~��O��\|�#P5E"�x�L���� %�]5)?ʴ/�"R�#G�{m�n$��cRJ�QO.�/Lh���&f��>�b�"+�m�
r���I��"��:v�׿i�����4_���>Hw�m"\ �Fyt��j+�-O��Q�f�Ñ�g#D�yg$�����d�����r!f����$;�n�%:�a�������o�r7����7N$���(We�&K���'�Á"*�����]�9���1���3�E6��|l����Ȫ�`c�V���~�_^ѕ����%Xu	���N3�����T@!��@��7�qW֗O��x�Ų�Pʏ��e�&�{�����Ɨ:�I��̟_��-��fy�w/͡}p�����O��U~�6~8���o��@�