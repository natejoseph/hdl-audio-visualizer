��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C/7B^����y��u�K��w$�M����C�JŧB�� ��Aji@DKuAU����a��U�\�v�g���
R���LTʆ'�ˉ�O��v�4H�C��l�sV�A]�;����!p�{��m?��,��.t�Y࿑�W�I�>���Zꌾ���/�t�t��P��.�(x��vM�r������N ��e�/V�E���_����V���2��.�v�;�;N���rPM����-R���������۞�}��tj̛
�
�񧝜1�Q�?��[O\�&� �m6��8��9�%uA�����5����I�A �?����p��B�/�Ɛ�5x�M!ڭ/x�/d�dG��ʵ��K���}�5��1?�`�#��K���<�B�NZ��_4)J�����<��U.�R��l���ٰ���jīT_�D�@%2#��L�����0N��e��t�}le7�:�g����Im����0�m���S�<��D�#V�ƴ�%����=�Õ�������`��1��F~1�JM�U��鿠$�~Дz���:�`��^̀7?���]���ٖ0L������n����0و�m������_�"f�z��8�]kb�JG��S�tU��"/�$�^������W��T��2�g&�vd ��3�=�p;���.�gC`��������4M&j���L��D@�*{�]��D�T�Cu��A�h^��B��{R��m3�i�KQ���dmN#��Dμ�ظ���8�w3�"�Y��c�@):���̲�KW*jg��J'z�k@���:ۧ^�)K��������阁<�Н_��M:\�	3,}_�����<E�P��GO'�7t���;���4�`��t�稂�[05)��I�O�|&�N�t]_�a��]|%s����EYȧ7�h�����	��B2q4�s��ϯ�!z�ʫ W-I��2�f�X�۹I͑*c�����b�:'�oE�T��	/�j)s0 ~Q�$��^�!z�+'����Ҧ'[�'�P�UPJFJ��bO�Gb�A���Ή�撇Pڱ{��]3�/�95`���há<�D�;�-�'�>�)J�o|KQ-��p�k,%�F�,Mxpd���8�B�z�x�P�P�s���c�c��N?�a����a]�$��1����#����]��10�Q�Α1����t����{��:���I0��j�Y@�Qp*��.}!���v\��)��E�U�<eV��Կ�)�'��5�-n@���_�6��ۙ$���`��Z����Q?L��`�~�]�䌨���1�6G�+{��v����i\}3c�U�7^��.���ٶ�åZ*I���8RqO+����F��BA��a�*��x(Q���Z~�H�v��+��UjR�7)Z�����'���y�O4��є>��RJe�y�����\d��;�kf��S#c���]	��>Ҍ��e��<U�ͱ�.��x� oQ~�9¾��i�/>,�ד�-� �_M��	H&|��M~:���"v+�w�����0c�H��I�H����_��_����o��ip�T/j"�[�����Rm�3�uhI����C(68�aQ���4Z�䨷^��V�</l�4ÆX^���zX��-�o*��ʪ}��� s
�����5&�%�S�$4����'[Y��S���O���5�F�0��uC�F��5T� � ��@���曲����0��-Ïb^2�j��	9�+H;�?����Ĩ���!�N�F#��O{6cd��;MCg?V�ڳ�/���#�����E����g�`���6�`i����$��8��� Y��3�+3q�р3�\���~��>ө�[���)����Q��M�!�Z5i�My[�FY�m�)��q�[�K�e�(��Xf��7�׿.*�k���:^D�\���d�i�ާP�o��d��z��*d�.��b30��<� �I�.?�I���í�E՟���\Fa%��(XË����KrÔ�9��zR�n��y,��yD�\��"����G
qbR���9�m���Ѹ͠f}{I
�[�?���R��˛)e%���W�4A ��õ+���P��%gx
�Z�(�������IG��^�&�,��a�~w?��D�O3%�ό�Q�W���&��g��Ync��ݪ;&���Μ\έK�Ԧ�>�:�<w��)|�� ��B�xm̔���j����*��m��ț�C���~�����
}�����A��f|8D�����[��D͋�S��,f5�m�2�-F��ke&�P9F��c�8]g���$�r�c��с�C�Xo�^�l�f+_����D�y��%V�3�v>o9^�yk3,�?1�v�;dlF�����qM�^��7r������=�Gƛ)au�%�>�$N�F�C�dS�w�@�	x[6������sӌrO�;5�a��n��oZi*AF�]�r3�_�����y��6Y����&�[��s|�1`�x��*�t��U�v�u�nrũ��BE� �p�|\-�|����������1�ڈ��u#:~�Y������8G3mXf�y