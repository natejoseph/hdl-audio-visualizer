��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��2S�W7�&d�c\I ����	[���{Ն���n#�D����������٧�Z�;����3CE�<%�&�Ew��Wh�H֗��Ed=JKj���+��$����:O�g�ps�o�)����������4Z7s�v���{��j���=�	�8�	��U��=���y{�$��1nP����	6r�f|�6���n;!&�07���ȅg��J;�_��"�y�0p��"�u��3�c�~�3ܽu�$�C���y�+|#�?���.w)ݚ�֝�\�~aNs_B!�Ll�_\�(n:HQ��"[Y���5�9!*��x���+B�S�4g�
U�)i
`)�׻W�+YV\PL� RK9M�2���<�X�9,X�ՠ�E���	g7JP�&:D����������/Ĕ��@����2��71�Q��Y�e v�~&]�	��%O+j����+Ov��s�n�^����H}ɗK��B4yS�QU����G�{��� ���Q��fR蕝�qԊ��;ǁw��%�����Z�YЬ�/g"���>e�Qz�J�J�l04�<����<�x\��)p��`��w���F�[�i���75�H��T�JB�6��3���<vI��;QB�;H]�>(�"�v�H0�΄i��/�7�3��d�'�.T�nQ��-�Q�a̗��c���ڒ�DeMV��Y�Wc��j��$�s��(eԿgE))��#����R]G�y�/����2Q�X	�I�!��
���2��5�p�"�.�	�nJ�� �}0d�C*�j�2��і<�	k��,�]����:��:#��UF�X2�Z.(����-˵a���h��BԸ)TT�ތ�_A�/�eAt]�	mN�=�j��P��"n����Ed��ی?��U[���%\r��oݩ3b�.i�of�Ut�{o�Xc��k�"�4ؗ9�7[m��?�6kw1��Tzyn$�1���"�$��9����ow���V9w�w+�>��&,�� �I!Ui�L~c�E��^P�v0��U����{�]:��d�D���o�x�����f����}2L����AP��+��F?Y�u��x����6�/��)<#�V��� ��y��'�n���K$�!��y&݄�a����F�tɬ�̿N��{
����;cB&��!�
ڲ0�q;`<���:�j^�ID�r���w�E\��)�)��W��Vp���V�uk=����M�գA���D��bK��`i](����5$��1���xdpQ)��B���|�wbq���]P^�.���'�Z �s$ϔ(Aԕ��|�����%�����Z��7�dLb�wo˱=LW%,af�WDϬv�'��W3�CR���3|�<=�}#񢈔cS��<��øc�'�_��C��f�L���f��+D-t�$��MG��[����e�����y��������Uzc�����d�o��!�{�6Z�Y
x䨊���T��p%S���+���`�߽.n{�]˹��@��r��V'CW)����UP�^V�W�n8�gW[!4����,���/ц��Р�\���Ǚ�y6�y,�۟u�Q�?�1<H�]'t�azF�	.�������8�
˭tŧ�� ��z��Q���{�U�Z2ȍt+�B�H�͝��	�+?՜�/�h_"��)���Њ]�`i����5�<�l䐀��b��FW�/�TP&>�6��:���G���ٍe�w^�(�.������ި6�G؇��؄/d_(���n���+���$p=b&�x8!?�^��'@/�1g>�)K��`�����p3ζ�������������[��C4���{���4h@�7�eK	�#��[�����;񒃡'�E~�;r���-��i�*Ϯ6�Ip#�G������ƒ���֓i$/���hꏈǨ��; �j��୉�3�m	T��� w#Sݛ�#��E-��T�n�.na��,v0�"���NMV*A}��Ø��D��]7�fG�G�%1�8���Sb��&G��g��N�Rd���ڶyvs�8WE"f����;���(�&Uf8�s#f��q�O<g_o��<�> ���'s�(�(����׵��1K}��
�b��"8Jh�I��b��Щ�-⨔~��r\j�4)_��Y�� gwD��#�	(�v�z>|g���;i�r��8�5E���0d���V�3������P��Ș܅�ݍ�<�;�ݿ����O���Bz���c�^"J�����2��b�@7��!:�E�SAn�c�d�&���~�R�r��8�[c���?�k�&y�m$<������S��Ķ@��E����t��p,����'}<wG�+����M�2�,�8�������U���q"������5�ț���\d�'�ф{�7s|��ΰ!;�-���@?AkpB�#45q1�S����) j���;S�.�^+7�R�^O�X�O~���%����V|^ئ�Mu��͗��;W����婭r�  &@���FNV�wٜ%�$��6DU���\b,L��� �daF)bEg"���84�����Z1?��͕|��dO!�?X[�dah�7x>��<;�,��7�ܮ�`r�/Fb��<԰x�^�{�nUDm3�[\cv�N�����
����S�fǸ��=�v糉��)�BD��a�{�������al�$����ǃ�-Om�>�o���]��H��M ����,|]�Ы���ŋ���h�{'���韽sz��ː�ǌ>�����s{DB�6;V��0T6!nJG�?#�9)x��0׎j��� ����=/\�h]Y�_�	ٚ"c��s	fM�W�����O����E��F<b��F���!��u�t�m��qDV�p���6,��GSo��ꉹd���\��A?,2����,��R	�7|�I*B��, �7�();�<<~)߽�0V��m�^t��I�j:����8Y��PN�>xi�͋����i���&a���ҵL�Z�+dڱ�����(�ƅ�B`�IH�_=����ӡX&���f! g�jJp`����a��]N��W[�����Џ*������R��09Q�@;���Qh�>���5����J�<|��k5lx6ӌ:��_�LW���h���˟��l'u�˧����׹�LH��z-=����K3�j�<��r=��J����������,����pӆ9e�q��VDٕ�\Ѡ���*3
�{�N����F�D^�m��X�dK��EW�Jcg�竹.���%�)�zP�I�L�A����]�Oc0���3`��:ϻ�M������(j(��r?�2��g��m�2ąH*cbG�}��]kڑZ�)������m�AP�z�%礀K9�8,K�u�e�&.D�Y�Jܖ�#آe�ٓW���WG�r��FxɁQ��Y����ri/�m�ZEaw�\��Ú��]�+=C#<
]��/�\T�s�5��/% ��~��]��F�dvݔ���^?����t����s���Uu C��Hg��2��9��:Y�a9W������?� qr�OtK�W,��/���O��N|%#�lMF��~���T���k����6-y8���s��B����J�;ƃ��-'H�]��6k����WV3(�_�$o�x��1�j���J=&��i3i��H8�A�A��L{ky�3sw���&����Z2�#y����k�j�{C��Roa�V�� <L_[ o�# �(�iK�Q�`v�&Wɭ$.
�nV�kĊ�c���n�����|]��1an�m��A���l �����RC{��O��Ŋw����d�,�����~��k*���J�DT���7#���)��%C$=���M`"_���/x*�T��[�"FI\LM���Rⱖm��&%�yUk���{���&�GI:��{"���z�D3
���R][�����MXaӰ>(�ST!qb��½�`��������<��>���X�<��}�u���j�4����A{���$������3F.#ʿ�VA���� ��f�����}��д��m��1e{����%��z/�o��x%�و�楃�������$���cK�Uż-�����bͶ8x�xސ��y;|�6�j�H��NY�Ce�霉;D�:N��M|^���eFk� �b[D������nH%Fk���!%���zn�l�x��p��9맔�弙�HR.�\�ƻ|�C4%�r�Xqڪ�\�6l���Px���4�ě! ���s���	�[1�$���O�-���(nO!Ts|eZ[�(��I��&L�YY��R�u�Ter���?R�-0a��}�h1��Hs�aT^- �JQ� L��m�Q�l�s���1V�hN~��C��`�c%���ީSS��B�m'��������a�Krq�^��TwRh�24k"'��żՋH�� b�j���{�`��/���"���u$��,�L�=� ujz��w�C�5ιQ����q��5*���$r�bn�?_Z��{i���w!.	�*P�������IƵ���XC)a��]�`�� �����s!�N\m��T54�[�c1��	.E������w��EK5Vk �>ዜ]�S:�j�6#g����[z��2�V���^���ӻ�ǉ��]�I�m�<�ұ�Z����s��� ��^�Ѿ�ԣ�5� S�|�b�G.@W�B��k36���[��)6�z�8�!��UV���J�ѵ�P-��Wgƈb~��ʒW� O,N�����Y;������j�{/S^s����4?c�`��)���3���q�o~�6�b9s��6a��X�`�X*��V쀑��%D����Y(�F�7eU>�RQ'oKԴ��-��������R�����d@�{M�)`�A�?m�b���G�9�^��df��_��W���E��P�F��#Ϻ�UN<�+�ہ�Vs�2�P;,��B*�6����xT�m��]Y�W�)�@�T�3��C?��ܝ�gc���*�RT�����}�T�}�jm`H3�3H9�W�����gƢl�sNjt���Y�$Jv���eS�?��B���e�� @D���qw��{���QF�R"[�l`M˃c{}�I�Z����b(�O�9���Ss����:��I°�Z�Ӊ��md"bq��W�[ƅ�dZ �=�I���\^�9wA�5�f�zb]̓�Eff6�n�NW-֔�̀�9��i�CyVi('�5�2s��G�Z:�op��~�@�}N4���A�#|0@�sIQ�2�1I��wL�f3������b"������a��5#H�/�O�{d�B�L��YWF�0=6����ΰ���k�%]�?E6�F�w�NLʚ�w/�.%�I���9���ί�H��{�V��fM!@8Re�0 ��H�)���y!�#�S�	����t�2Z�5���?�#5��yN4�P��=��B�ʺ.s鯒�(n��z+.ս��]�sy&H��O৤��	RIo[~������zQ�3�0���1�|���_�e�P���6�b`'����R�.RJ����)�+�r��N��ww$ć6 �0�Y[)cӳ�W�*���ft�N���+Dڮ�UCw�xb� �xL�S�T����������,o�w�o��՚����I�M~7�'k�[�ztְ�� ?G�W8�
q�Ƃ�޷�FNx�Ʃ�j��ί�v�|�V*e��M`Hn:�/l�F��L�RK�$�xO�iT�&�"ڍ�Y��GЈT%S�R�����ڗ���
t�,l#!��Hx[^�5Fal���'ݨ]>��pv�tT��7�e9�/��كج��^5������Fc��C���x�/F��Io�}�����J�����	y���f��Fq�,�--�-ͽ��\;�82\�"�9��6�AE�r.�1{�%���f��K�Ȕ	3��ҕ&=o����(0�)�ͤ� ~�(.27��D)Ω��w��8N��$��ݴ���7�/�|��0a��&�=cH�ғ����y>N/M���æ���.�)���iح�X�*zO>2�e(P��X�ن�\,���|yAe���#R[����%k8㣥�	1�y�����b��׬V��	�D�P~����ٙuHI����х��@�_��p��m��'��a�&rޛ �'��[�L��c{�S����F~"�i)ǹ��j����6Dgt����G�/�r
M�/�����I3W\#���w!\ ��R$s���b�%02?Y�j��I���U�DT''g���;���+5��q���YF7�������#�Y8N�;�)�l� �	�s}-.�a/��dy�#�݆����j�Y��2^�: �ę��Z�ʈɥ�]|���~m��2��(�v�
�,	�ʷj�4;��7���l�X�� �W���0f�
�p�uQ��8'��,���]�a�M\X��E5�y�~��6�P����&�$�,���*ʔ�!%j��{���^՚W�T��̻�Z�_B7r8�����EN$�1���Nl������7���t;ʅ�`��:\���w�2�K�����f���-F��*^�e΋9h�D�'hp�1yv]��ħ���6H́	��$t0:#����3�mF'4,B��{'��n]�_Ӝ���y���?����Rն�(��"���D+i�̨7�H1�$���Ůi�%W~x)i�P�!Lw�
��J2G�L����r�X�桖�� �9���O���)g��V�L�P��.i�'kYU|���.��G�-��*D~��ح�z���"��͗G��B�4�h�;�r��Ҋ����x�h�/���8,e��h�5�\>��b��H5¼&���j��F����%�:�H���Ì	"��ݻ�n����7��F��|+a;�I����K.�P�ѡ�h�Aу�g��U�^��l�y5-Q�'tB7�Y�!������..U�>]V��܄�-��(L$)��r����o,9]ȹ�E&���^�Dw.a^�ûX�����6_� �'���-�f�M��-�:��kkֹ7��_$Dnq\1�_+>a�jo�-��?T��h����؟7�Wf�u��q� ^8]���E����N�d��8X��[��x���֘i�?�{8؍��֡�e�E5����}|��0�õ�6�M �|�9,5$sѭ0��aJPcm���^ʚ���*��\rٔ~��6{�䀗�q?�����f���d�˸�y�u�a7.,�C�IF����#5:r�	k���A��U.��˭
M���U ��|F
���M�A���(0C�^��0�{�\�06N�Ԡ�d����D��?j��)��2���|%��9�0��~o.��k!nO��z�r���݇����t��p�+�!��OkK��{l*ߺ��e�pyp���/>$h��Z# �%�!:�0��Z@��u!��I�d�#=ǘ����(^�O�j���� c�gI�G�
��j}E{7�r�-�R�
����^ \��N�,,���O^�/�1���|��;M���)S8��
Y�:��V6�=y~�F���11�w��'�fu��ͼ��������=z4Ʌ�$w[�R"ফ����J���)�ז�Qod�+-��'�Z�5��TҒ�-�O��r�X�8'ۺn��RYn��~H-/.� ku��-��S[�n�Cܕ:�ح?u֡��څ2t~�ÙH�Ntx�Z���r�n���G[�\P�{J��ޫ6Rؘ3.YC�]ՙ�ٗG�4��P;{`;�A� WK��n�v�ES�i�1��h�F��z��A��d���Y}4(x�7�`���IC��Z�g���ʁ5TR7�t�Sz�]Ë�Mi;`ڗ��D�4`�����pa���62H���S�}�٤@��v�<���5S�!�67�G2 Ʈ��"c�Rh�P��k�77��6j�?��<av=�qsGA�%_�	T6Z�L���M�(�-��Ai��AK[!�1(P�ȃ�o����A�T���n�u���p��.��`,����b��K���$�f���'UUE�LZ�Ь����W C�	�L<�8��M�/i�A�X��pBM7�V@~T��b)���^L)Ig�\��ɚ�P��iĴ�v�����>�
��1̧�rdC�}��a9�܇&��i��=ìH��7��V߸r��h]la���\�t����E���s՘.����]�h�x��18{ka�uH�� �z��gRz���M�/�Z�K���;��(�`]b��7���7���T��=g��?7;m�n=��9höRl]�����o�^M�ᾠl�I�5��d�>-�ꭀ�R�h������>��:_VY���;ԥ�?��	�T� U�RM�5G��Ό���r��&m���"��;ǈ*�jR�u�|3��s�����F�l0c��b;�_bf��d�������_����V��j���j�P�?\iBzZ�PI�QrC���'��
�}w�Y�D��F����
p��b�o����HK��"��-�"H�l����}�q^�t�dᛎ2��ܾ�G8]$&f8=i�8ol;�eg����=��CszT��	<�M+g��v�~�C�CιN`ğiM�,=ռ-�a:i�nt��̒ee�n��4��v&���"4��ѡiE0S�7w����>�y������d_�w���WΟTJ�[V����t6�p���V���~�1�7a�L�	��x��S���:���;t@���� �������֯��u��욅�=�j9x,��D�d�j��q�Y%�r���SjK9�h=Kf0� ���gD%��I�cL���S#����'x�\	}AFvfO�DQ���T�z�G�Pɦ�@����f5�b���X܁��3m.��*
-o�#1*�m��<��kfNҬ(!�x�}�d��PX!�y���,��e�p\��ޑ{�Y�k���u�p�ܚ�C豶�F#��lC��cg��WZ�VAJ��2YX L���)��y�����G���N�C��7��ςPp���*:�ޥsX�PW�*��x�֌�=*${����<~t�H9לc?6e��7��R���Kg<��B��y��\�����P$����QԼ�6��X]��YZ��
�hZ�:����ϋ2'��"иY3�S,^@�l��,On��U��׻.�|�tn�GD��	S�@����{}I�9a�Q��
�M��u�bL9��U���KX?�'2�B��$�i�BŃUm¾��ʧ�L+`�0T���>1��H�1����go�O�:<&�/#}��C�{周���oIE�nT��	�6@k��켤��ˣ�����s�����6�@o6�:�AO�IO8��*vn�\%n<Đ��\��t�#J21�	�h����1P�Sɸ��6"MSA�����*w�!�:s�����C���T�O����X}V�u!b��Vv���l?ba�:'=�fLQ<k�@r���u��ω)#��~L�����)����/�����L֥��o\����Dj�[����[�B��I�[z8 ��mRD�)�b ?���T�Z�����ǿ����q=z����Mct����X�9G��-�f��s��J)�ђ�N)��h�[�ʃ���?iɲ���S�'����D�+r��4ӏ���U�ߧ�7���1��������F^_���~�9�u���
(|-2��5�Z�`�f�t�4w�ե��*��3Qe:v�I!���*�fI��0����o�B�4?�0��P�
���r���o�)�~ZDg�TTc�y���.&��@�'"s۷xK������ᩑi��'��E��/ک���Z>��E�j.��9e�_�7�8\�7Th5z1�G<9������`�2��66T�5��.�f8l	� �0�m�����h�S�
M��Y��P�{i��C��Gw.F@"�%
�eL�����ѥf�⸰>6E._j������W�[u���3Տ���|��Ϡ�	>�ei����.È��a���	�q�����fl�Կ�خ���7H��Pf��K@��;/� 5�k��@	��oG\c�u�φ�y���� ���!rD��zo���M��H�7a쑉j>��ԁ��e7�,Γdm��M�����@P 3��4����|\�}Tg5Wך���t�R]����Ӑ�烿���o!�5�R�2�4T�j��/קf��)�Yy���I/h�V�L��gs�W�6�H1>���.��]�h���1���݋�tF�1��\E܈`v�3ً���7�`buX
3��bڐ�[��b��*��{}�Į�lL3<����V�-�njz]�iv�&���1�B`���4ɶ�M����!�����dF;�S��T�	�
WCԫ���C«�7af�6ۏ?`�'ƞK՚��&su���8.2�sW�V��%�@�2�Ři�	�U��zT6fܤh�Qk5?e�4�T�j#�>i�΅ tm]�����B�h%�	%I[�ĵ!!�Kk���T��>�G����1�|��12 8��'��]zz�eN/t��D�.-c��:(�?��E�8ž���H�	����>�Z��(ܴ��/��wt۟dQ�R	�g���ͪ*:/��7_���Bc#*!�^C}�j�w�K|
�O�{��۞���Zݣ���P�y����D�Z`̲�j_0JQq�	gջ��^Q�2y�,Od�rr)�	c����g�Y��/�=%���e�fy��.|�t/�����O��*V�O���i���\蹀�J�>��!�Mcrd�i���\���D.7��'X�˾�ԅ;�姡�Þ�٥j�`�l~@:TS�7h��Z(�z��$,c:����mw���G�S�4"`WmN��s��q��I�
�vDw{(x���@��h(<�y�[��U�H��q%{�Β���+=�\��/N_g��
�%%�?��3y���ˀ�(S�-+|��l�d���4l���������c3C9!0��[R�K����;������he}垨�L�L�N�Y�/K0���/⽍}���P����%����?M�2t���<TO+W�\�P-U�����p��� ����^�w�uYi����������Ɍ����ii�I���ǘr>ļ��U�o3x�!<\���RKh e[��?3e������4k[��e�������,����B�$�xҬN$���?�?71!��1�JZc#/��E6;-9J��^K�f"pЋ�=-���e�.�6�}զlX������=�`N�~B�\)�v�Q��Y�
\���^%O�뙮�?�&�u#��ɘ6��Eш�C��[&�$��#w�%�#��¬���%*h�\"��Ԥ���>��^���u��"C)�z�ؚ��J�7����>2��~��e}����N��h�D�0] r%�Ȟ	U���4�����nx�	Nc�h��++ҹ�&�m;�}��x���w���]}��~�"��ȔH�05�ˎb<��ގq�`O0{��:��G=�.�=�q	fJ��{<�mp:�ꂬ3��g{���l��630d�<UN��#���m����^����i�kZ'�R@���1����QǓFx����)ⰆdZM�k�l�z��[M�	���y��ە�Ru_ʤ(JDau�aZO��M�9<����p�h6�̣B_���c=)�OI�o�0%e�5TL�1��ps�1q��M4t�E�W������|�s�<R^ �I3_w����z	�<:D*T	�zp�Qu1hO��*����t���Wڼ%B�`����)�B�fm���4B�w�҆�T�5
E0G�d�>gy��_��JX�����6����C-'���<�n�7.�WϦ�
2) �G��m�̖�鎙|�i��y#�0?�ͩy�e�^�c�iqпg��"+K������&������ւ/;�'�~��N}>Ջ�@��)I�.�WOrp�y�R�8~�5ӕ��l(��(:�
�?� S�CzS7F/�ws�\���KH�Ksh}�U�+>i]�T�|����L"T�Q������hx���P�� ��\<i�s��� dWY��$E=[3��F4�I����#���}��bX�u��^� �șO$��Ϗ6]�m���	�"u!�X����N��xΨs�B�Zf���X8�����H�1И�d�b����&@��L���Ϗ���SA8���"�/z-dR��e]$�'��
����Lg4�H'}F`!�	��^O�uSΉ|$�k �`ڗ�w�P#Kh�7Ȉ�`a�2	�fL�%KBL���*�t�&=���I9�^��o��>9iJ�L�b��P��J9�:�(�0���X�Ұf�'���A�46�B&r����XM���i�����f���H.�J���/\�_�%:�C�6�҉��:%��J*�}˼��Vt_����CY7��w%�����s�N7����Q���=]�9�#��4���Q�c���@da��R�9��� �,�١��U�F�����#%��j�6�xB�<+�2�3�uV*˧w�_��Qp|&���[�y[vRfoF�Ѯ�vS_���c�&���;s��\�p& u$k���v�:M�G�@�?��7-A�pPp�}�u-*��"�MV��!j<1�2�ӝ�>�uD�W���YSf���r�