��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��W��<��9�<��|���#D}e_5GD�[���"ev��W1�+���(ͅ�KxFH�尦>S�h;k� ��oݨ�$�0�,%���'�B �P�>"�h��"3�Kq&!y�~�+G.B6t+�mƱ��6�j،�_���j-K��~����`ʆ��f*B�~����_��y�)�I��'\ւ��~r�O:J��m��"cîX*�[���q�DVo;1���<��92��+�Bww$�y�ܭ��r"����F��l-�+AډFI��)�2.�R�ug�j��?�;���c��®8�H�E�S����K�Xq�V���T�5^J�������^��:��	�����!�=��]D+OhnEJ�x)���Z�q����Y� ��?����k(�v;�(�#k���Q6���"6f��"ì����ʻ}�;����I�#@20^*d��)X�Q�?E>L������)���<�"Z�G�:86�n&{�[FS#���nS�R8��������'�t}{(Z)�r)j����~��k�k���bkQ�n^,n�BoB��w!���rn���ҍ_����.�m-�W+��b�N��r�\:*��; ���3d��Ye8�<�.c���jF�+q�:���L���$=�o �|�+��w�79�G�C�������	�U��@h/��8ߤ�u���A�ߴҬ1�6ӏ�����a,�0��7�>9�m�)��j|g|���ۍ����D ���o��p��I��
u�zI%zJ$��_>�m��6ϐ26,ʲ+�Ҵ��͘،���z�ժ_�8	|�� pz�b�\~/#�B��;@S��.���K1J�`��wqI^"y`�������g+�}��CE���:�~�3��ց�#���	�g��͗%��[�س��������g'�Ϯ�d�</3��{.�k��j��{�d�e�
�������*��'�k��l���@Rб����]Es��7 ����˨*��"��WNz��bk.��۲�"�����F�A��+�M;E84���P�� ���zO���}��&/ix�Tc3�lĲٔ�V�M���#ܕ�:�&�CIa��7;3�A8���Ŀ��㫫�h;��$�R<���E���b7�mb��$Κ�b2]Qcf�ި6H�.��Tf����:QE���Ѝ��g�pQ�H��mb�H�!6�aeU��ͪ	�E���1�C����t��ܗ��4��O��Z!�\�%�9����V�ߧs§�	������w#5x��'���X�yr��tl��}�v���g�Z�4�u�4�e��/H;@к`��L.��w��oQ,��Z7հ����2��1��j�)B��,z�$=E.�H԰:s*����̩\��e��YL�ў�9���
�	R%������Tu0}�+�.�^  �V�A��IiaO|>��6)vabL�8�Lu�/h��{���b��Ǖ���R���(`c��,�27j�x9M����OI�����f��<Z��EB���\*�i��C���F
���v�������l!L���Y����R�[p(�07qߧr��v�~�F�#�>m�Ak��('7{	�E�&-QV�bBy�fct��0�g�7LeK�gǴ�8�7n9CCY��F�Gɞ�����gxNy�$�
7'����Ҩ��)���fe�V ��H�Y��g^8q$�c������-B��4��dS"߰�q%	a>��x8T:(A:\��ٝs���&A��2�D"���݅N�$�خ�m�2E�_�I3-ť�:Fc xD�a�wVR��A�����D�yt��5�7��A�V1P4�K�$9l� �a�F:U;~��:�ܕ��F�	�w����i��Ҷ�X��q�3@��-]&���t/�yHVBnkD��g(���M�]��jȱx�C_P�(�⦠��܎�]���+c�
�C�n�19숁F�r��ܹ�z�c?�Q:o���ݴY,�k�/zō����<#'
�7�q�06:g�0Dc[ �.[����+."��,NCdf�/@��E�ٙ�:���t�;���MU;y-�zi�r�֧|�m��F�Q?��@0��@�2P���i,A��K E�n�������l���+] T�c�U:v�u��us(�A����;�X�
I3bn��p��M��oČ6L8���)�.�N�������#�)����ᘖ!���X-l.o�A����`�l��9����k@]0C_v�u���&\�޾�;�2a_�$u�&Y�Lb4�CǠvV�9"'�-LX�t�6��K��t�?�$�ߖ���D�Q��KG��g3�q�����)��/�n�b��s��$Nqp)*�	#֟�B،[ص}�������t�	h]52f��`ƍ}TꝍR�F��و_�l��۝�qH62]�i��j��E��4cy^N�К�R����M�(�NYO����d?���Ŭ����a�/��6�W��h����
�c�?R�r��E���=Ik7ʎ��,[�'����ʱ����YJ�P��e�j��O�E����c���
)�GF�*f����M���D��x)\����Q��/�F��]�N��Vu@�l������e+��X×T��@K##b8=��+�n���*���e5L�09���J�e7bjK�j�To�S��B:�OSrvX�����&ǝe�k$<�
�]z	dҍ++k���l�ر�=�W,�!�|i!��b���[1]'�gD��e0�g�s-Y�X��U<^�JQC��AY�u@H���]��R?~h` @ӎ��^z~?2����w���,�_nȽE�i���h��̟��3�e	m=��HJUe,�e	u�~�m����!���s0P=a�@�?��Oz�O^=]�t[6��_�I��N�$躩�P�ݑ�@�7l�a+Œ�c#rUqf�Ua�өך�[�;� �	0���̗A���s������`�'��`��Y��	[M�ONCB�JY��`4�i��yt�tmE��+�OYf>�����=|����=�1��Y����֘�����f�x���K��!�Ѵ�����F��Q2k��쓵�.ܶ������8C}�d(A
������J?(�|ML�H�d^ *���XAOѽ��h}�S
m��Iӛ���b@~������u��<6X��M������zP�0�E��rs�$�M�[2�4� �-'��N}�F�6����Q�u��w�7�,[��uh��/�*숫��&�HܛI�z�Ao�qA�F��ר���I�M��0�NTG��YB��$�j���[����W�0��}��b��f}Zi�������mN��4���U�9�p��R�^��K�������A8��d��E�Z�MP����:�V%��B���i(�K>� �AËcemX��������ϋ����5�����44"8�]r!��~�|)x(b�Ntw¹���w��(�kP�y��������:oF�i�ï���7TۼƦ����O����.����h�G�W��̢�d���*��t6s�N�u����4s����a�Q�$s,Ǔ���a�,����j���u��2��'��۶�j�Ҁy�M��O�7���<�;%� �}�O�5JY��X.JLT	CԕwP���`Vk��p�d,@0���(�e��>�_.Z�XY|��N
qXFt��"����,Ե�L�V�t���a3ݻ���7���B69��=7��.ș�w,��:>���~��`�$���	�b͉5X&�/�Wܧ0���	���ڄq/�X3��Ȁ���-�`�|X�6�,�_d��r�?���������7�����}J�G�)qݱ��G%�F��{!�u�"�f�r�(%���Ql�����թ�{t���>�!�8-C- ��x�Oj	=��  I��q>��k�4� {��2��v��2s����G���&lnup�+U��v�}�2����m����d�+� {��:k��qE>k	��;)D/:���2%��qj	�;,j���e������H#�v�� ���!�� D���E�W���X�=��	$SrT�	^�rOjxK�N/AZ�N�	�K�%o�D�G���:�w���l�(�V���9p+9���k溲`�x�-ׇ�{&D
�����e����p�r�Q��}r`�삏c&�q��� �W[4�=ӧȫ���7b��*�񗬕-�⫬����-�u���?;xxej�4�����vzb���Z�nll2�h�Dm2	��/�F�b��B�m:�-*;Q���&�H�9*��X�n6Z=����cu�Anmӡ���HaN����D�4�n�<b�?��p� �׉O����ה���o��z��W�f��x(����7����T?�)�Kr�~���Մ8y�v\�
U�"�z?���A�Y�E����=O�!����46�[�ԞC�879?̭�E_"�
.UE�,�ʵP{x�ޚ���^U�����s��Z�^z��70��!�����W�㬴�� l&��Ϋ�E�,9�yZ%i��i#�/ݻp1{^e6��e�~���+&m.�d_% �7��~3y2lΚ� ��Vc�^8���e�"���qr���rD���
���=�jCh��&s~���ڦVhM�snۊ?����/�� �S7�m�I	d	�>r�[c���c �N�N���૫�i'�<|2OP����tr��2ג�����,�r����u���6M���R>��SS��:@B�A~ٍ��s�(u��b�'�8���;ڹ�����l�ؼԉ7�$�A�M��rj���)Q�3�2��bY��N�%�/���ќx���V�o��`�!�(�9���ZX+�C��`�J�1ſ7,�y�Cʱ;�!",�L��Qþ�lϐ�)��MͶm�Y���G4�$�^\ql��w�����⃵'W�2H[YX�N��:`L����M
��vq>%���<�o�D��mB��z�=K�Ȉ��q�z]�J��l˟9]�n�t9����9�:�P�.�׺���XӰ�����|Dckwӿy�\�"����������s�kb�u~�SbJ��{�'��v��qO��ۘ�פŃ>�a��#=��fM�u�����+t!o�KҦ4���Y�d�l#��m.��f2���1�*�^co�U,����ȆČ-(���|ӳ����qsm�\�����
����v`Y�&h��N[�w���&�)F���=��$�_h>ﱾT
�.�K6��ژ��'�u���)�H	.�,x���ڋ���L�V����.�R?P��7��P�l�y����д@�����RD��y*8H�U�l��fTD��O��U�$տ���,P��:쇢9��I�
E�3^y�eQsrՎb��/6t����a�/U⮫��+Ѕd�/m�W�}V2D���~��2g����DЬ/�'�ɊW���=�y�*��ǯ@Ȭ�C���I���]غwL,0�T����m\��98�ܷu�+,�4�S:�����$�|>lb�]U�U��Ȓu{c��Z�ܴiѥ�@��|�u%��9���âجI���M �^5�t��p���ǰ�.����"~��'Q/�^N���%�h��� Q��b������&������Y�v�7��ئ�0��'py�y'�3m��mc���o� �_�:/T���9aa5cr�:����U�%���c\>k���O/�w��e�wG%���p������6��;�S�j	fX	u������{dx�����QT��lE䚱;�L�AV1��	���߿��-�"cUj�R��G�ӳ蒑���P�%>=�Z$ ���˯v�y�n��쭼��0$9��pAr�_���[eF�0,ү�z��� &�}ȓ-s� i�~�ڟ.53���O�;��"��J�d-2MD�V W�`"/p&�V	[|����]��UP��P9̂�[)^n��	A1Q��$v�g���^xF��`�3C�Cp�Hu��3l�'=�!��'���ӝh��zt������zT�W��d*�[��gQ�m�-{F�L$��~S`�8-]A���eR�4Ly���d��3݌R�`Jɡ��P���3L3���V�PqEN��V9����w���w5���cV�;�),��˔hC2�9��&����P��/DR5�R9;�C72w/��S���g+7 z���f��@�z1Ukc�L�xvsH]������µ��|V���� ��JT�:\s��itE}���Nȟ�-������+_�Hn����S���m~�ϱ(��O�	�����u@�(�@&�ֈ'��P%��]�ߌ��x�%0Lp|۶�	p)�y�W5�8��=�� F詚��F���ڊ`�\�Bb�j�U�I��=�� ��{��ix]s��u`��ײҚ�[���?{�q4R�5u�u��T٦�W�Vk5�7Y�!"�8�A*H(>X�����pZ�zl�ޭ�d|�jJ��٥���mYn�{���BY��d<"��Y�!##([�k�i /�*����S�*Q�2��?/|�@�I�$�2��tM�gM��x�:;n/���ūi�]tF��;����v<.�>Y��40FsO	ɹ�z�%�BR
�m�L��g�&��������E`���sZ 3G���������XK��GB����j>�E����|8|nw��y	!*E�ů�\D�P��ą���T|%@g�
3�A, XQ6\N��=���",��%�X�l����9e�r�N��IȰN��E�B�VI	�Z��B��b�O ��dd�_�z�����D-%����-��/3$�-{̀m����'vWh���n�*(�2CU= �F;�����x��뙽� 1��Ne��H��a�Ӭ:�3�s�����Qh�"wK*��#� �Uaԁ/0ND ��DL)��n���Gi<��c�K��0�Zq}�a�kpІ��a�9�䉌m�z�afA��ffF�Ft��DSE�'@��yg@�(Nb�f~޴���Q��@�)?�y�y�p
K�ܖ[V�e�����̨6R@�+;��oc���	�������h�Y���.8�߬�%�ہ��ST��=D�T��7�X1#�����]"8Zh{i�b�Y�"`���#� Ģr��=�X���t\=�E0b#��T��"P�u�����Q�ŗ:��Λ�;���F�����G.��_Rh}��{-;�����B���r�J��F�t�8N���i�8�-��dnL`,�93`���G�Y��cw+����6���}iT��6�Zܰj��K�qJ1�i��O�u��k��[2��u(���}��ܞ7/P>�oX�^�#?�7��X�B�B��8�Y/�=��j���J�i�YZ��I�����5���9�mи��I�>�ek��:�y~�.8��7��^e��j��:��ֱ����s�U�w�@��.��f�?�����X�X@.@�ZYxH���	&�Z��u��uBsQ*HW��::�M
�f���
\��W����6��OM�G�i�T�ˋ����.u�ҷ�$��I'R'�AS	�~�b�P��#��훑�Þ�f�#U��~��w��Y�워���>G	!�ߙ���3���L_�L�tI7Or�~jm�	��7�ߚZ�s�
��'��? oW@�a�ro�����Z]-��i1�_��r��`�C��n��b��(R�^�s�d�\L�x��\����ѝ�mY^4�:�53�6>��fĪ�	���_m�sa�w)�h'c[���P���D[��-��6����d �r����hHTq�����;Px���>!t��0��Wl0�O?���&Ħ��Jf���G)����9�{��P��E���g���C�O�0��X�[��2��!�:4��s����ܟu�JJvs���ei��{�I2 ldD�RZ�tq�5��m���S��u�G��'�3	�y%td��f���y������bäA��ϑr���Kr���D���3D|��A�{�yZ�A*��Oj��Xԗ�>�qEJ`�'�!VXkk��u�A��b��R�t�LB���I�[&J����9s_r�����撹�{>���
\ɇA�O܋pc�[Zp�!����S�J��I48����}�=$sy�Gh���*���u��%�ӳ��+�?-�	`��f�\�X����=t�W���w���
�ۊ�܃�b�"�B���g� �L�,�����?W'�����D���o�����<�|Xґ�ڻ����P�P
���L��[1��ǥy�cy�� �C��@�[m�ی�3]�f���r�n���	O�s~~{�e���Ǣ:�9�>�p��&X� ��ґ���Ɨ&�V�KE��֋��Z�G���z�(,����!Cy���@w6t�n���pq�B��������R����!��s�.i���k��;Cع�4\����}KB�^\���G�.&����RTu����1=�iE����N߽+�JZ �S�����?a@H�t)p�A�C�P�b�
x[?v�)%���OI�����Ȣ��?�����/S���Ƣ(���n&�^���b*_R�Y�yת����gw�����LЩ���cLUvMF�����#&t��,'���,O�{s�.I�P��t�L��:Cx��#���m�W���fFSkR���d��@�B��V���ǥR�� N&uR<R'�g�C?��vq]�����������-Y�A�'���?֓��!�b�v1�_C��*�g��(-{7M�����L��%�,���=�F����ֻ�p<��U�U�L4$�lX���J���g�<�s
��N(���F]���;yIi�1&?p��[cX%㎭����z�*