��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|Ci.D6�p�ϕ~������jt�9@��]�HjY%e���i�b���gA׽�đ*(4N��<�l@> �,�B��z�ʱ�����pp�6u�����e�`c��Y��}�� �-�F�_��4�68b�F4�o5˺��A-3�Aբ"ԏ�A��Ư�;.J��;̡�)�c��d{����6U	���(�����{�1ƻ[�?
9���و(Wd�>>1�	~��t�,L&>���>��'�'�cvx��� �:K�fF���%~`:��+Τ'[U���	Y#VϨa�b'�S�
��4o��6�x�����&��� H��8��:\� ��#�Z�zV"���c�d�C�B&�F���({� p��m�sq).*Wxl�;��e��;g�<�eʈ ���{i�ޡ�����܄|���g���3��ᗂ���
ΈYo�8[*�۹��r���r�؂7����tU���x�[���8zf ��R�!���*�P�1e��}�7Q�v��b�H���S)>�L�_J��x#ZvTd3z�P���Q7��$dE�뎍��rh�)!w��U��a}n}xc��6�I��"�f�u�6�Ʌ���w�����q�K�~+X��B���ފc�g�Lp��;!tr�y5_ؙ2���O�<�ۙp}(�H�#1A� �'`�x�%j���1����6�$�� �����q�̔ξv�s�ׅ.d�a��O�-"[���/`xTKݥW�"O�;}����N���B<���1N/&Zt��i>-���3��Ut���$�L���=�H��>r��o.�wt"oK�Y��z�ȩG*��}n�EV�x��D5�-�^�D���'O�`�ʬs&�2���n/��F#c$x��_b����D�>n�+�g��r�4���k�7G"X�z�!u2$�O�R�Q*�y�&�|E���Иl%T
�����u��[�#�K�� ƕb��$L*�tu(��@�U�7%�`��(�67���29�ث�G4���s#O�w�s��CO�I3�:P"K�{����M�>�����I��$�l�V�},|<�q\>�K�>�	u|w(qk����D��ZV�b��	�PpOZ'���GAY]�UJV����[B� U��v+N� (M^D7{{b}0Y�7��`�[H�Ys�m�'"�I{�D��܁5�܌�����Y��;RR2��7�W�H�.J	�C��&��ܑ����즶c��]Zq��o�t��2�Dd�Nny�Q�P����GNAO�]a��f�i��Ϊ�:wuX�1��/�8%H���ٲ$L�kUʎ+֑��}#��jg���b�s�#Y��e�P�,`Z%s�R&Ǻ��2(��>~����Qd<99#?hq#8�b������s�5�Z�G�F���W�Ww��M���^��o����R:�f!ѮpS������[Ȗ�3����*I�l�qt��A������_���e�D.[t������L0Z��숂�D-%|ϫ�$eh��P�g�j�3�ʷ� S�	_ ����C�݃�"������ �}��1F=��k�L���5c�1�C����|���ZG2���ļ߁|��9䉧��>'�g��Nt�M����+���qvрO�n�J�XGl�ָ0J�N� �:�̒�C$s�����s��HS�����Q���]?��y[�\;a:1&	�<����;���ز��c���IS��Ҏ���֜y%�Z���z{�)7�B��2W_�=���p������yb6n�$�x�؛�@_g�{�g.�Q���:��x�E昛;�?:���H3D=p�s2���A�i��2����|�аZ�8�QW�4��x��'�tIf�qq䒬�z�d�\���>vx^SUш��N���}ّ��7�~"�+`��Yw��*f����;�^T�|��*���r��Wxh�)�(�<FA9�k�=������"̉��]WW>Dy�[�#��FxZ���I(��R8���)"�J�ea�T����>D�ſgy���xG�hQ����߆yɠ� ?(�hߴ!����|5ک+3�eJ���4Â�Tq����ǖ+�k�+%A����0e2��2o%w�������{��ѥUD�
-%5���3��}��c� ��ۨ�&�� ���?�U버��!+�a��jj�6��c��\���['��>��L/�{0�W j��~�PyF��~-�0T�=1�w.Jg��v�bًG��:�v$��bS���p@0n7ٛ��gx�"�s���Q�Xrp�Mo�U`���@��b���cY�c�k�<6B-#u�(�A�-]X�"2�'�g����haDÌ&�!�?��(�Aˡ�WZ8ρ[T	����o�Cq.<�UYWS�ݥ�럦%0��P_�?^~�=�8��f�t1���������P%^�B�D�5Tz<)'I�I�󻂺/!	A�k�I�D�a'Ψ�BP��u���4n�*�s2^��$'x�M@�ʅ����b�&!�$�ûv�=�G������]��?p�V]�|��yf���Ǖ��F��5E��eq<|���W��G��\�_{��⦦�~;��a�]l���f�Ս�B�r�u����+�2|W::l��[���&�5����A��d�CN�mm���J��Ș��A���\�&_�8�?PӈR�Z���Z���f�rѽ������ߕ�j�˖.X:�eˣ��\�]�ݗ^#��U:=�(����:�mP���T^�+���[:S�% �A?�I��@�����8z�ei��f�%�C��t��xqP���<r��R$2{Ú�Ѡ;�Ey/����kB�z4�
������W�Np{�H�i��9��ô��i��sL����#����²����,�O]��]��^�j���2�;��n#�_�$t�L�G Kh?�`u�y'�lk��H�/V
�W���G����'���F	�����q�����`r�$�cW[�.�ړ����-t�\�XIᘖ��VV������X�D-�=���*Z�F4�����2̤c�-���b�;r�)���%:dr��Z��v�r������	���Zތ��;��҂CՊ��y��PSI�>�Az��U������ujI�\�w�%���p�$o�_yw�($�E�����������e�� ����N�b0�K�c�]N�Z��0�p�>c>��`��0�M���RPy˪���0%�ٖ(TEy^fN��7?���8@�T��0<b����B��� [�#����j��w�!� mW)< �	�}�	�?#�ɼR��Ӧ�p䋘{���ѣ1Bۂ>@�뤔��Z*+8q*^��4�oY���m�e�t�4pf5�����l�o���Dm n�h�0�%��s c���+�!zߵ&�f�m�����b�λw�L�1ln��6	�n�K/h͟�\����ߋ�C���iK�g]9��6��j���c>(A�zx�%2�w�a&P9�n�r���@�wd(�Uu
W�f,�n'U������6B�f5y��<�8Dl��t��	�Po����X)H��V��J]�5� '�h~YGF���	B:L�F�FH[�0!�T����:��8����H��5�Ƿ��6�^��Q���H��N��0�m��
{_��ѧ���3y	+2s(�N|L��ê�\ddv�Ⱦ9L�.�%�Q�J��R@�Z1�CH��M5UU��Ŕ[K�hԫ�=˛#�B�}?`��G�"m��'�ge�<�W���war0�>9�G�	Q�:s�/d�.'��I���<�d��ٷ�s�QQ��e*�u���"�����eSF��n�!�ֺ������T���2ϛ*��K��?S�`
�W �&�L��ڤj�y�����t3of++1>�$���Hpaչ��1s���|DS@���2W� ��0��9mc+��[�a���n#@�P��kG�9��G��31
�'1J����u��w���+�f�hA
W�`���7C�M��2�Y�j�R!t��
�{T�jA������Ƈ��I�a�wbz���]�zq\��Z�@�i�vY9�'v�]TTw#�`Ji�����~Dljdc�'����=��<9�q��~�t�;^t���X�r��G�9��`�0z�r~�Dcc�\��6��ł���,e�+UH+�|���wDIfC�