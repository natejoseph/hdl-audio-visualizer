��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����;* �{pB߆�1h�L�e-�, ���pPt��ºBZg�.�D�хL8��u����k�^�|\;�?H#��%�5���!����esUKd��K"�q�%����#�p���L��z`��kq�	��qY��`QqwY�}/p�N/D���s����^�S�8d\I�R����	���`�J1o��_"�Q ޯ�Yک�A°���b��O	'C�f_��U$�4LQ\w���./�|�Sc$�I�ʈ��A���S}olG�ɠ���l���i�@��N����q8@a�Ү��AS�>|S(����28��;O�Tc�*�w*�����J͕�?�,���=@u��e�^.w@o(��Ep&���\�+��UT�!4�@3�'��N�7�CK�E~[
qB��l3:����&���&������r�n�#�K#a�<��X�������!l��c�b����� OP��a����a�<�*Yr ��i��KӖ{� p./���	���S������z�I讨��&P�vj�Σǘ����pn-`'t��sCf�����T�L���3�Y1����CR��^��>&����b��W�ŋ�>D�u���t�� �0��5Ƽ�ye{"R/*}�ſ�L�;�\���N����y+[�쁸��mxTM�k�x���Ч�m1�dH��?-"�;$�yq]�,���	$��9_(8t��UƊ8̰;��k�$��=:��b�M*=�q3�to���2�#�OQaͫ�=�N�Q	<b��[�� 3���R�.!�X1�uhn�������`j�N ,���O��-�HnҘܞ��&�� Lgv~/�x1��%b4G -V2@�\C�����|��So��JX�o�|s�Y�R���ł��cH�/�!�x��rZ�I����'
�8���u���l=M�8<qO2YtIv�Ӡ�Z[��-���5)��8�<\�҉�wSۇ��Q�z��Y��o��R��`���1��r/w�b�j��5��֧�`+mJ�rdZYXPؙ�ó��{3�g�K��8_��XZ,�Y2R}����L�����Hv�i̎T�s5 �����m��G!)��(T�I���m9���?5�x`��M}� �Ƭ�s�-Gp,E�C���2�'�� ��hDL�,Tކ����8��xhLsBDpƶr�Z>��%MO��6���"�Q��7�{3w�M� F����՜ѪݠG4�큵t������F��0�~�.�ݣ��}8>�z�=�''fD��(��,�r�ܽ���/K$������R�B���j�\�=7��(2�d'�Q���[�H�X��Յ��z�s8�;��fI����{X��x��N��Ϟ��E2�柢'�G�6�*��������P��,?�Z�%6�ʌ!Z��♒}��ƣ�?����+��H�5��nr'��?<]�"��]���pr�������i_U�w�B��y�h4J�1r��F���I	$�Ss�z�#%
ɓ.V��-��s���K�G�O#4��j}Q���5O�c� �	t�l���D�<�Z����L!�YN������7�R+SN�p��&����c����.��{�a��5�`J䥣HQGa�G�2�X�U0e���3LXZ���f;�>F�r�g���D9T�K}�Y»?�3sb� {�#W� t���D�g(e}!��`<Ũ+��5�=�E�?�{��Jlr�}!��9��ݟ�s exǪ�qPY���o��'�.A==)��O��&z[ގ�]�kiݩF����]�+�]P�u[�"?0��������2���z\�9'az�1v��e���d��O]���aob��[�skW>;˲+���j�;eO�����Ho�F�H�8��i�l���2(�ƐBU(#�#����9Qo��UFw�l�dp���KK���,��Mч��\�L���EP�*v+~�ݬ�{����"r��=��ց^�����Rh�U�N�	���cd���ԇ��y��M��$vq���gԅ��}�zS�"UP�㎨�Z&��r��J���@��1"�
���z�qZ}�CM�Hv�|���S̄hH���距���nlР1�sR�!����I�]����ҹ���exm}28����6�V{�IL��G�� �\�;���
���ų��{�נ՗��m|��͙b��(@!>\"��b��}�J�;$��O�%�(@��Y*�ը�j	���7$��E�1ϼ89�s۠4.��c�`s]�E8�`tȄ���R��`�Y�?�����Zc �J[����a8n*�Ԥb3,�W_�D@ S�����V"K�Ϳ�9�8W�[�u����.�CM�)t�ћ�q�]s�A5�O�V�ԟ=���1{D\�2y�i��'�[�����[���jm&�hp�c8pơ�?�(�Q�"�qv�P~�#�s��劜�<� �=u��x�H�9ȉ�_���	L�GV�1��m��r���qfwj�T�K%���IÍ�d�^�˸�Y�n�Z	���0bؼ��W�C�i,�4q�"�:�~���0(��,��)$��N$�j4�Ț)��i�we%��ˢ���\	���>ك��Lq�4��s�':��o�T����&�����~g3|$�0)f2u*B!�~�n<D�vh���d��~�.~R1�i}��om�����7(̒<��3Μ�8$m�������Sܙj��l٣E�	lv~��[�\�~	1Ƀ�5�k���D��Q��NdǏ-{Tq� v�YD�Z!��5tgK�\Ua_��9H�!��!dG8�*e��G���ҍg�,�倰u�j��7�/d�͏>i&tDAzu݉�J0ُ[���Z}�c\䟻 �� 4�{��^U�M��~f�ȑݤ�]&��sF�:⇻���4�oD��Ǩ��E;f��j��
��c2�]I:N���З��n��Q%ba�A��rH>�UT����ƒ�3�� �*��e���� �������S�8�i'67R֎��z1+�cK@e2��}�_9 q7�p��2c�2��n
�S�~0a;�$mN=O0;}C��ãrG�8�e-�y�<�9���! =Ș��X��+o-��fqIH$:[�TIƩ�z�t'ə�ˑ^���4O�$��6�S�E�_-��&�I�6=)�����檋�kJ�s@e�5͋���Wɹ���$�M�P���d|O�Oz|��j}�ᪧ�"F�O�@���"bD���^��[?(��dǶ�I�����#�ʰn��r_��6��j�v�?<���״a�����eEC�v�ˍ�E_N������.��wϴሯb��^�K�f}�Wk��԰]�~b��C��LdI�֓=R��nk��{-�uTߙp���$�dR={�LY���|L#��D}1�@�����g�VL������i�7��5��tv�f�p�Y�<6�C�P��t𡓵p,�z�Σ�;γ0��\�:��m���Y�y�#�G���u�nj�:��e�H��x���
e���-ªg����Vg�u&�,�<�3�m�w?��*�/W���Љ� �n���=&6��q$8�.D/���� �5e^�E����D� �̘��I�q�&��ʲ��5���^�D#�q���m�W��}x��c=p�����u+��M�&ˍ��mm�)�,E?zMF���`@�LC��hvE��<n>{@����P�aQ}�/�]��$���"JL��c�l�uBK�1-]?�|J�RW:Ld�r�i�ɶ��X)_}��[4`���3��ž\P��� �Qjg��\v��>�Z�u��.͹�`�1f�|���U���x��G�˗�o��Pz)��^�$����|]��r'@�U/R���' .����!��g�{��� ��癨)�ŤA#�U��^��f�R�-,-s������,,+�g4���" ���G�����/,"]G�h�&��q���E�߷P��[��	g���"�Pв����V5#3	l��z�DH$g9�O���v��)���A;��I���A@��*�����'w�\�N}D��"��tI��z�lch�缟�?�I��!6�\�n���VD5_�*.�Z���%��:�*a�cRJ9�=ɝ�Twk�i���[g�9U*����h�ӮL��A����4hs1ȃ�@��N$r�$�P�C+=6�?T�ã���6֋w1�?N*]�Ak$�t[0�aq��M�]P���hɋ�;�#�A��i���a�L� 9|'JS�e�q�&O�u��k !�F����h�X�s��IO=�Y��o��ƌ���3��
�s�>�-�7�+Ԭ�>��j��Y���`ǴvL�@t£a�فܹ9L�ij@���Z9q͟�159���Nq]����zNJi�p����u�@��UJhݏB,5��������fM�A^�� HT�e��r�gWt���r<D-�u^��TK�_�Y��W�f�D���4��Ԫ:�\z76��*�-	���@.~������WXdl#0��ШJ� �o��3�%�����yu�7��?+�]�eYf������{��F���>R�7 ���3���]�0�\�G�j�N��1�T��%ҝ�}?�@d�����i��S��z�n�g�q8��Jwע��F����>h���ցh���� 0_� �RË��O�
�1�A�� ��&���E�<�
v �tw�a�g�XQ���DJl�+�Q��>x�F'��zF��ݢ�"B�\����{8#;�WL���J|�
�J�q�B���Q�H��i��H�ߓ��a~�ɩ kІ��\N�!skU/��ꧤ�fv��@k
���)�n��YV����/s�mX�ݑI�c���{rji�uC[~G��N}�Z�n@$�"�J��x���՝�t��9����b;��3��t�D@Q�k�����q�G��'e��-bOU��� ���>�8f�^��8���߁�����fu��&�`q�O���5�8���$��9KM�g�R,ɞ���Io��R�r����LL"Trm0-��6+�=�!^��=��;��"���	��iX�$��"|�ʨ��S��Lw���Y[x��gvɚ
��?mn
�l���:�>E	D���>��>��	��WX����n�l"n�e�Ȉ�ݩ`1ܷ��5��Ww~-N������V�<�����%���+.�/R"�����ئGM�V�(�}���}^A���W��Bu~=qw+S�t-#<MH�qI�h,����/�6�/PTi8�=�-�*��M�DPn�����¨����{�vEZ�Wl7�?��OGZ���8K���O-tMX<
C
�{;�7�R��LJq��Y�V�L�=E��d�iG�� `8&��6�i�Q�����8�����n]G��0��`��z!�@�V�W>j�^i��&���]DwUע�{��h�BaM��Y1��:��� M�R�3�)�W�gFdE13��բ
�)*]<��w��i���g?٦��3�ڇ<kY�{U��������<�]Xm����p�UhƸ]x��L�
|:�]��N�sPPH��E'�uq�É����=2}84ߛ����(����"+j9yF�h���O)7���ʘ({��X�2�6�Y��Iǁ֗����!զO�|�ڐK��pGiw�_���hi��?�*�j��du:�xX$�Ĵ��6.$��*�d?ֵ)�)��K�U��ӊLՠ</�ag���U������9 N��À�� 4��!*�j<x���n?ӋZ?S�|������ 8���'��\����_��p� ��ld���e�/h��ؙ�~�-��)�(Q_M�����fi���bH�?24�\Z���Rm_�o���f�Ͽ����s�9���|���U���=ш�&�?8Ӹ$�o}A���Q%�-�u!�g.���Smǧ��|�����.RA@�P�������\�;l�����WqW��^�l�`�4v^�ЂJ�n��7�D^���b��>�0y��ko������3͸�F�e0%�:i����5y"�4���p �rČa6KY�v� �s��T��۷�D�Q�D���D�T��'kg�!�Ƕ\W�X�Xy� �nア��]d �I������<�K`yS\a����OD��o'����aU��8RJ玆�$��i�*���ޒ��ap�Vۍ��ۦ�����gg`�q\-R/0�
v>B"����=�읟�;d|XQ$@���ؙ��S`N:�
RL�:�u��/���Xbġ^���[����=Bwۯ���v�0��iy� 儦`�S�ۖ���Sz��T�e��X��S�yF�z��d,A1��#�2Q��٠��8Μ$�?r �7��{s�n%�z�1U�q������Z�9+����Qy��n4�9&�ؖ�?��>�5�0������9�ܮ��;��ޭiig��oA۝�{~{_g����KkS��%��4u���{{�v�Z����.�O=�Nћ� t_d��z��l��;c����S���˕]N�����J�²Ѐ_%p�M�-3AJf���a,b:^�{L�s��Α'G��Cg� �\7*m��1����+ޚ����F�C��Y�y�T<�i�(2D>�!��N�2�.`�� �Z&���m�n��?j�:�Z=���9M&QR�;}0G��²�֜x��hO��~q�u�4�Yj�����9wd;�ww�,�RRf;q�o&w|Q����� ���6�Y`7
U���L\7�%�ͱ�f����rCE��8!���b�w�e1�;�ii��l�UC nF@���� �$�c�����-���:�V��9���n,��H�v���A�i��_y�т�O!<C:�uqu:M��Z����ݶ� K��<���:�B=�%x��� 2��B� ��h����@�".�h���a�� �����Ⱦ9= ������[����7�`'� c�T��Q6���ѐ���C��	L5F�T?IT�Ñ�a���U�/��=�?�J�/�*�.��?���' @<p��:��1�vN�`�>��Fh��C[��=�T�a���BS��@~9�]�dȞ:!xDqd�.$�zYq�~y0�V1��(2�[C%g.������C�Ħ���M��(@�m��Ц=��0i)y8��^N��t����K蘩	L��3�����¯H��*cxcJų!{�s!_��:����=UH=�ܛ�*|;=�Y(��/�%Xo�C�ʺy�\>��9�* ��<���ar�Rr4�3ݫ�x�-�=c�6�����z,�V�iTu;�j�sY��,0�h;�o��^���lTU��2�/��l&W�Uy_�%89����1M�Kr���|�ٰ�{�I���**�!�r"'���]O��ߣ�q�0:)�}>�QY��[�_?�/��+�1V���'R�>���Դ���=���%�	u8��V�����á��g)��r+�}\P���<6���c~�4e+vha��VXj�M��4����XĘ�VTڑ�#77�%o�Ej�
(;�	��'�M�æ���Z��$�KXs��8ޖ���?����9q����46�����9)��槄#�:��ՙG��'G����^��C�'Z�C�h�|��h����ףUq�}�~�{{�1�2�W���,�.�{�A`�J�i���5�P��T1��.��.�?��v�ysU�o<�ξ�D����/���o@^�h��oI�?�c���H:1�T
��(t��(y��j���9/��w1�[Y9�Rb$�E���`�"�Y\'y��c�j�%J*eH��!O�"�&@Q弪?��Ʌ7)���^&ܾe=A۸I;���M�Z*���XEm�M�`��O�9w~�ބj� !� �����Gȓs�� ��g��wp�����R(�<O�}�gK��H���9%Gm�W9�ҵ���e�N��IX�6�vo¾?��)>�N�����M�5�3�GF�gS9�D�����Kn��@��qX�M>C�����w���&Z�fGg��y�-��$͢�1�}oR+)	z�z�Лs�&Ci.y%%�9�\?ڏN��pXF�wE��8aP�e��A�O�v�N0x �_ݛQH�ѫ4!�����d����X�[Z��W����Y�@9���G�k�We,S��-�H��LѪ��T�/��0�i`�]A}��N	-��4�E+��	g�m1������j��w�q%T����:�ڤ9��h��_Yg@���.,kJO��͇jT�\r�^R��U%"�0<T������=}�v� >}b��<��Mŝ�e
�7�(��I��r�9]�����R��/���=x���m���'������rl�5f��u�:�8d!o�ef��u����ٚ}�K�SְD���)q�� (�(���x����|��r�� r20�$����U�:���K|uk}}@�����`�?�i!i���j\H��0~ d���P����fo��5�]#^�%@XH� Q��x�b�	�l��97��p�P@Ʈ�ˢ���8�;o�<�耤��_�"�>R�f���"j'��eLw�M� g���*?�\n��J�}p�j��e@<�����JH ٮS1���xG��O�ߕ�+h�k6�}������觺(�'$��w.&�����֓2�w&�tȹ��y�DQ+c���YdIό�;?Q7�@�������b�q�S��7b�r��5�.���E/.`y�NǢO@Hs��"�9!���'�?��]�{����Z�Oi�
@���/��iN_J#�1��I�w��r�6�J�P��5���q���E©�Gj&&f�<K'���:��d
"M�Z�F�N�[Δbde֝�ugV�H��?�-5�;@<��N^R���A��HЌ�Z��T�����{������Y�	����X 9�9�k�.o�%mD0Z�n�C������C���]^b�xQBLʿ��*���|E�䟙I_������MQ+)9�[�d~ŵQ�3����`���ٜ���׺lZ������������WoK��-�1���6�b��Д�3ꧾ�'M{iQ�(O�B/$��{v�����4���G��Y|?�wH�{�/�t��w�=��L<|K6����[�(
1�˵�&���/F�{��of!6����NiP�Ƥ�/���e������+0U��xm��]�.LM�ݕ�u�������� ��C�4Y�1�U�σc!%|�sp��XZ��ټ��P�L��H����Ҹ�r�F#q�d��l���Q���͂(r�'�=��H|������~"!���ܔ��J/}<��jR�U�D�ԁ����3S�k��|���5n��<'�H�PT��v�f�T�*�� ��!��kq-��CY��߾�����m7�� �T>����і�U�����V���=ey�r5C�_R;
��x˶��I�j�Z�Ç�����`�Fs�������$iT��"6'�H*���S�*r����zW{��R�3�nz��h#+e�|>�VW��&k���S2��q&�j>�T8h�_��t�[-�49�Zۚ�w����@���8g'F�5DaW�+K�r\R&w��.��F�9G�S�QdBG��ԇ�j�Ǝ:ҶB�#����|�D;�>qk���<�^���1��B�|����)�'�iI����(��J%�}��;�ȌH�+�J�\o��g�#৐���ҩc�,���Me5x�.uM-��`�i.04~S����{`��_�� p�I�+��bAv5b��B�T	��?����=�2⬊�L0j4/��eKP	������v\k���K�ۡA>�=9�ad�7]PN����
�)Y��@���o��#��dH���sp��$Շ���d풞� >�|"��!�klP9��O�)&ٌ0�V/���"#�� � #3��;�6��F��~�ċ7Yw�R�C}K���3��Α��Fs��2�Z��=�Ee�f����:x�*/����԰q�$�?���
�8�u�ޟu$�Wmq�� $˄X��y�.�+i����ks�9��6D�Y�C�s$�ƴ�4����wF=�|��2�T'��9�_�º�#�����r[�(��K=\�;Jl��_a�+�'��?m�Sג�0�8Rիv�����S�{<�\W<딣ao�lT��:�9y�s�F���ʦ����'��@L��&�h����I�~��#���nU�0��>ʒh{xb�GU��cD믛|�1$�������KJ��u�ͬx�.g@a'9�������eFloJ7�el���V���?7��n}�;oq��w+ܩ�b:���Y_Y������x��A�ٌ��A_�|8��$�"�~�Þ�X���z�]��p������yD}	��]YA�_�&V
�9�q�����e.�����s�f���ܛ9�5�t� �4l���&���m��w�|\�jh�	��VH|�w�}������,.��x��"���k��K��h�/k!^AGZs3Ȃl-P����:3�b9k}���?U^��E�� ^{m�b�q/��o�5m��J��p�%�
~��g"p�h�ǜ�$�rp�:dm��o%.�����c��VS�`�78 �&�h�wӿ�'�(��R<6����tK:�*��T�ܸ�|�\��-��ˈ�-�����
�Oޱ�����)e�IT��`�&�r����&��d��B�Xy)GmH���"�M��藞�YD�L�?�����R�O�ѧ�qkk}�� Kó%Y.�X�z�D/��rv�A�EPJ�1�n�
c����M�A0�27�zor�Ni�\�\̮ߐ,�ju�ͤMH�K^�^]1�p�Һ���W��vQ��Ɍ1Ty)
�r$��l�,�YGG�I
�@���˪T6{�V%l(��l^��D	9�e(��%��oce�Cr�����{6�,O�l���q�یhu���U���v����^y���=�g����g�Z���i�zI.�Q:����Hs�ڛ��zǸf��I�ˏW�e�����%#.���\eי��#��@�<D�^d���T"kmj�X�W�9Qg�Z��[3O�Su��0�chܣ��E{9mLi���8���o7o!I)��=B��/�ҺB��9
��q�\3,x(��^����������6U����"��X��2G�m
T�DΌ�U\0:%S7�id�c��R�k���+[����o#�)=��Q�3�g�C��r��&S��_SѓܦV��� z�������E�9��i����Λ��l Tщ������rPJ�Z��}s�_UmD�M7�����-�i�����i��on�}6Y��7�a�)~GB�n�0΍��x/Ǫ�S��2����F�xGsKy/�?�Z�9���lQ��L�o��q󂿃֞��$V^�7�����\�y��UѾgb��%���
ͮ�[G�ܠ��(����OG±�HN7�]�+�ս�ҢXy�R�C�;�<�rǋ �yZ�W�5ؑ0U�=go�C�M)f�\����&��gf�AZ����Gw������q���c�V�Z��~�Z�$�!8֦7J�����;gOD*cAn���$|90�x�w(�\�������RH�r���A��ײ���*�A�MX������x�B]��qf�L��b������h�1k��ZU�]��s��E/O��
e��-�Eq�)W���m��@_�6����O�^�]�+�p>��k:l(���6��8��M��r,�)��]�u����	e���FM�ݥi]����������gX�LD̞�k]ˀ���2w!���I�=rpLY��8��Dt���w%!�;kBi4�����i�W�Z���q����IC��v*OXS�^�Os� ���q���ه~W+��n����QӃ�?L3͐p�y:RQ����C]���Y&3�5�e�z��XŃK�|Tݶ��S��<O�G��g�R�g��ǖ������@J�7���mw{v�nwĕUb�/��������^V h�]�ci�&,�ڦIT%�6�?ž/!ҷ۪�[��T��rU��3M��I��7u��~eØq�kƢ!��4�Hj�Ȟ=a�-�E��x��,Mꃔ���h�A�C��K[��L����
���4��>�厣� ����
����r{�[8E]π/jL��j~P�N&�94�j9?{R�m6茅`��"S\�	-�������0����,���Sh�(}��1t�Z���%Ԣ��qM[ ]���Y13@eA��U% &w:¤��������Ae.����N��o��W�n��f����L��Q�Xn4��|˕�����̂���?����[!��?��������S��1MaW����I��,;b֕�S�3.|?IG���Ƥ��ߣY�⟤
�c!�-v����c��l&+CA��<��f�"��tZv�b�4�ʵ�ԛ��MܑN�y"vt��N�
����������Jh���=���NkĴ�Q�Ϻ�Œء^�R�b�5;q��ؓ�_��T�\c]��7�k��� ���~�YP&�o�'^�
x㕄��
���^�t�o��/I�`�pz�%�x,��b/���g@�ʘ��C��v�@,��5�h�ĵ�l��<�<L�]�)]q
��ނ�S�6����~�%���Ʉ��r��L�o��;����_'��խآ.�I��`��D��5'+�c���0�+/D�V��\zy99q�A���8�j�*Sݑ�6�*�R98��P�CN�M�����깭�YY�g��F��f;�[��n\~R�$�*[j �aw�Ϣ�R�G���9�M��}�&��;�,����@���~9W�Z5e�@�}n�kc���A���[;KʫW�Os8�����^c��ڜL�AM��ϣ��y�3N�)fK�p[q���ꧻn����������ᎍ�|���	�a��r�u��Q�pԔjs�,�RNXSu=&eߟ�eR����6j���t��
Q,d�AP�]�h�"���|����=qs��Y���-��3bJC"|X��bs�@���HF�:��J�	���G99M�x�։���e�oD3����>O+LL��J��kl�9r����.��8�C`4���.m��;3�y������.ro��8�o�.�?1z��������,,��$+Y�q�� �kVc{ë�9����2�Z�>���B�G���H�+>�/]�Ā���0�;'~��~�I�.ă�t~�~~��_P�M%0�wЪ�U�a�a;��|�ĝ���(aÇ�1(-�-���>����?t����p���pl��һ49�[��Q�b|�i_�G%p���T��̏���pe��y�w�v��z}���#ְ<�.�QPj�l� �=WM{�r���A�ȸ�n	*��>�Υ���y�B���ƚm]\���Y��QA��C���xJ����r���D�ͫcܮ^����k궮��O	�Y�C�G0�]_J�d�V,y��fxC2Tt�u�L�ik���C���{��6�WRtX�ؼ��A�+2~�1�z�%�C=K#�bUj�!��S�X>}dcS��~�ps�ϑv����΂�]�	d��5k�Sv�
��H
�!�\kM���|�+9�E�����g�\��� ODs�&��0���ZI/�yz#?������x|�6��-�}e�p]�龒N#wi%�,�Wi��`)huxQ��,dM!�E���$�;��`B�=i<�t�t����s�	o��Rd)bw�"���I.���e�~]��"����H�P�c��>�<��*�fc'a��p�ծs

��{���{�%�ѓ���Іj;�O�!/�eݵ��G�M9��N�����ڴxXh��:����9ٲn�XZ���(��\�b�*���E+�隞H��o'�6s\��v:rN����h�Z�(9�ZD�a\�=6�cŏ��q�fv����@�	�)�f�GX\E/�������ctk���)jt_��~���x��)5�Y*a�5�?�v��\�n����q� ���\F�D�U���9�CW��iZ	�g���x&�b�K�<���'L�:_� �f7��bPbL����/�F|(ZXL;����Η~H�uX��\1�j�%�i��Z��8�&,��rAZT��il)�i�>	�w��j1�!%��E�lۉ�S���q;"��ļ}��D��qy$}���`ɛ�&�>-��ϩ�&a�0�����P�~�r�n��ݻ�x~�Fyx(�ZHtf���4�v�b��j�q+��H��ީWe�զ<NG29�I-��s�N��8]��~PS��6�B_��qg��!#���Z?m���O'3GpJ@\[��v���+f��=ê�����ݮ`iG�F���� e�+K.O��{M� ���3vs�D�y�3=&���p��.0� !
��T��0g��*_�d_m:t0�4+���G�@�^��2���͓��> sj=�����_]�l3�pR,8a�""M����7�����b�o�a�&薂1��8Y4*�F�R5�hf3�㚌�h����&W��v�2��M��G�^YN D��:2,;����Ϗ��Q����#d�1�Hɠ�+�-�����K�]�p����������Fsh�*���צ���������o�g��*�d��~����TF�
���'C��⑎��1�7��*���|�=4�JE����
�LX=r��(�+!'����.�JY.+������&�žwq�ܴ�����)�5�Óp,��L=ܖO�#]��;��l��#��%��wlz�z3Y�,�ؙ�|�����fL�P�&W�@�Bُ�
�;�N*oY������5��d�1lɖ��^L��kDaǂD��@�#��6J�\����bl8�
,����w9��(oX:�k�"�`����%�I	�M/�hF��Ѣy����%N?d󻃨{�;|�rU[��%�w�mg��L�Չ��g�XRb�y�Aڬl5D$ƷԫW�[o�v��A22�Q�8_4ki�ؿ�.�}�z��^:�8�"���@�\�S�G�᧒���}��d�c�"�n�E��0���Y˞�Q�����>���=>�BD ���5|��D+̀ԤSM;�v��H�3;Y�|?  K[VMz�YQof�Ml�͒*��Gpuh�Gq����VHM��R`7Je�#:nv@rqi�s�����F���'٢^0�f'����6*8��D���I�L-a�i:�-��B=S��`tC�,xq68���K�i� �B�*��Q}��e>��Ξtvi\�pV�bVaء�.�&���ɀ]:�$�k�ޓZ-�#�ש��k�y��l����Ibϸ\���O	ʙ�P�ԛ�0��/|���j-%�Ai��oYa촅�����6 L�9��vžǸ�uϔ�l���w�P5�����Kц�1�����͂���I�:r����OO���!�?��y	P��bVK��B���a���vuN%P�}}��L7�H��@��A�f��s`�C��
A�PKk�f���T! A���ѩ����8q
���R�q�n������F���.��G,@�?z:|���N�4�7�I'A���r���,4��z9�Yc�
6��Ҏ����7�?eZ�WD��ӊ>��u9�eT	��QM�i�d]����4����zg�g� ��"ڭM[�;��
�{ۈ��V`�U�����g��^{:�q[D��-� yV+\h�S~y��Ƨ[�*3v�kZ��Z5�x�}�t����N�y<�r�C�ٜ����f�}ݗ����Q�so&�$H\��f~�����q���ݍ�#����$���W�Ap�R���A��I��������dd{���d4�Ek��f7y��қ~�a��l&k�h&�8���)�^��ߕ�-�	a��Y�*���wT}ν3z�`�`�E�0�\uvy*֎�W�4��^R�����]1�M�2��;��@%f��&�ì���u��������ŞW�xK>���*�}��g_\�úq�`fR<�6I�$�8��Vc��-��v!x��҇�=_aH��˟��
�ȭ)_���в� =:,Q� םb��m��lJ8+�Ũ����
.{W��ԛU#�Ko�d[�A޽��uk���oE�x��
h)���hα�6��>�99�[o���\Z�x�K=$uR�GJ�����k���aƹ�}�
v �=�>;	�!� �t�I9�O�لu+�m��>6q��;��vʹ����qW�z�����J>7��"bg��}�M�@�@]�y&� � ��b�����Ъ(���Mc~��շ�'fY�v��43�$X]���F݇ �5Тת-�uߊ}T�hB�7�w��^P>烧-"Rʯd
�tfi9�+��gF��ǈ�kձot_��	�1v����e��LL�2S�v��ȺI�����r��|���x���v�=����x��?�w ���Z�A�0��{���27]�k(-�Uc'�H��^ ��*R�*/T.�,�#�u4��\�	���=��[f٥ex�a���&u
��@İ�|��SfԊϕ�5#�x�ݏέ�G	 
�ô\80�=����lT�N��[c,Y��(�� �h��x[L�d�>�B��9����](��q���Dm0�C\������e��DhHϮ��
0���H�Fߝ
rh�8�Օ���� |�=2q��f�?\7�Y,����8��2%����ئ
��i��U|>�Պ�n���-�
�h��"Ɖg���>X�A��P��X� ��:�P�FT�6����G�������L��i`,ıO�i9�F������i������:8�w�7�2�u���}��Z���sʏ�Yg.X/�|cP�9����Ӑ���By��O馋TO��lv-��hU��T���(�"H;����� 2�~1�+xg��4���MUYJ��gve'�O�LtR�@����:�=�}��X��>�2姛M���jtn����V!�NŻ+f����ՇO���K���\�
��۴&������;t�L�mw5�d~Ȥ���DE�}9H����h �g��k��:�)��
�5]-�p)H<le��k������8�|,	r��Nmp�s<^�] ��La�<:��,a+$lEb�剸�g!�_�'�\4�n��}B�ۗ��S ,R�/${b)k����2W�{�/�@�}�r?p�;j�3�4Ȍ;�	�EFx�5G�34�,0Q�<p�;k�L���L(�e���a+}5�jQ����i�q�-�[L�]�O�cH�Z%g���3�i/�T��to�57ٞJ�22��p��Ă��r�^�NM'�:�<�	�S��	�1�L��� �8x��)�b� �C��-]��D�S�0�aVK�ɐ��M��'����R��D^����0&x9��;���{ ��>���S�9$CS^���D�f���7R�F]n>�^>N��Z�W#]t��
�O��e^�	y�� �;Sq�Q�Us�w�W��O,ٮ6��,r;E��j����O�M"K2�L;�9����(�T��Z`�J+B�����T����/�W�͡�7���1DĮ�w�"ܓ4F�d�Aڅ0�F/�64�=��+�,�n
%��O?p�bm�����"�7/���V�A !-��ʸ�iY��hK�aͽp�2v'@\���(2��)���)�eI�}$��N�fˌX�3�yO��Q��Q��2�>),p�f�E�A+އ{.N�WL�,��|6o�"�ƚ�4�x�N[�����H� � ���ğ{ �!�O�d�W%1`��v�q�=h_s7e�bL�d���c��Hu0�=�4��0�[���}%=�4�ݞs�ͳ�� ���7�+���lhPTD1%$Se��w����oI��ҰoC0kT/�{߹����+�ۦ����q�+���f�jë��X̦=��N(�u�4�Qv�e�g�v+�V�q�L-�;�7��}��o<B�9]x�;Sl�gV�J���5L&�Jbֳ�`_J���A4�S�UkyJ��Km4�&���t@(�x|�?��X�w�(N/E��N����(���$���H��=�'"�n�Y�K��M�`<b���1���γ��/��C��E ���\nLk$l�4��F�[�j�r�BX�8֭�jo�\�;�vҬ��� ���2&
�A�0m"�Ŀ��֨>=f=����d%ӗRqI3�it������'����Z2��9('�}E�X+U5�0�J�/�;���U`�Ha;^m`��z��Jҝ,r*���Q��x�G书��b%�D�I{.�Z���C�LmR�md|�Zx�q��q�r#�씒;��8s3"������w��+:�'Z�a��U�֔z˔K��bS<5��0*<��~���Fx5)�0��z_y�7��5��7�ք| ��;� �3���;2������VD��,C�f��	9'���z,��F^�˯2�Ў̤82U5jS�![��C�o��K�G��=v��|�;Y��j�"�P��R��?��Å��}NP����@.$�X��oyYk˘����-OmA�Nl�/
��*��(cll)��+#��1�X�^����X����L����.��^x����}���P{�kp�}�"@�$7���U��;�Գ?��&�4�p-�

샐����|;�����!P���=fo��
�E*��/�'��3��4��|,O-�t�e��������VE�����X7�8�/�E�,|����k$M�b�8�"���Ѹq�P�Jr�'e����h���rN� �C���8[s���C��`�.����O=J�p��*)��n�`7A�h	l���J�7Q:*4w�IdL�|&]��`K���d�n����[~_߾�7�C/�	<�)�'�K+��6�c� qt����*a����I0�54�M��di��&z�_�b$���X�E�km�?=�o�zB�G�t��2�����|��ߍ&4�d_�M��֣���મ&:%�_l֣%��||� /D���|��F�Zp������1)�Q�JHk�k�-�W�YJ΀X�V�Xf��d�\��%�'��plp�CPY������E9�wiB�|�3�`�� F�a�5�ِ�xUܠ�r�yA�W�و��fڷ��U��Srx}��B�?K����O=������?��r�P�s�j�f� ��.��Pʔ���E�z��(��4�(E9�p��f�?�J'tdT�Ƹ~���j��,Z9���c�085!�*�q塞�&IL�
f�����$�]^Jw���Uu$��&��k��IW���l��n��R�f/�x��<�F^�Y��kъ)W�Xh�
}��+eMq���W�EK1u�wSDt�9?�*'��Xh��GG��6� ȣ,ŭK�k�g���}v�6�M�C��vD7� ��}����Vգ��3N��Dk�z����1,@ԟ�����xl�WQ&�O ���!\0.�m��	�lH�K��8~>+�ʆȟ�n��B������s�E�lx%�������4>������oP�d��Y��Ɣm���y-��Q�-�$�SYE,#dr`�鐊[�m[-&���^.�:ɎAxT'T犭�dm���/�C`22�O0��Q����Lo7$�-M+���U'�īI�a��͹b��:)����Fgv�q�g��8���}֒r;���K�v�2YM���깕8���u��!6��ko�X����I���B������;-�4�u��s��r>.
�*\����H������c.��=��v�|SF��61��1��M�h��0wľҎ�܎����E�� �˿:0%\4W"�[����L�����@����0�G5�����D�k.��ʎte������%����]���;� ��ٵs�t�9a^C����������C���n�O&C��ڪ���U�I�<��m@2�R��u�l1�W��(CA�n��|i�Ή �Jr����@P�x�p�U}�M��1U�ɸ�d����c^u����N����UJ�탔��lj�S�a9�۩܀�����9������]}	�I����"b���f?�l���0�.�@&ӁӖ_�zm1�$�B� N��xؤ��M�a��9�`����pP�t�KWh���h��<�i�n�
�z��B�0��l�h6��D�����b�$PM�՞����f	��]�����&�yf��1p٨ �Hf���֙-K����C���Y!��s��&������x@'�Ȉ/�����ս��Z��E�G�0d5%�Dނ�\k�z7�Ǖ[;�u�j�Er`I�.hDA��و�wߌ*)�?$����"&2၆�3��Sڱ9�ӂ��qE�p{���T����"�Ӓ���+z߭�N$|��6[)N�~��Ğ�X���!a��K~N���,�a�K�K�E;}'�&�T�d#����I#х��7?�ovP�V��/`v�h�B�nzH�>�Bz��\���'!j�N{жc6T�r J1s�j-)�k�%}k�C
F�v��:��k�ܐ�qEl��~a�+�p:G���N����_�к�왇#X,r��=A����fC���,*�r�^����g��A,B'ju�v�^۔��>�YT�)S��@s��cμ�.� �*�L)4ª�����Y��y�x��.|�l��MQ7W8�����[�Ʃ�G�]U��M��a�$�A�!	D�GW�:�7�k�"�G���`��&g���Q�6�XH�#�Dg�DKm�ت�eW�?iT���X�/Ղ�l�&�5�c�D�F�Ѽ1� '�� �Z%��M�;��'^����&7~�q\�����V����9�+��L�a&��_��̵�\��_�-�ή)Nw�
ƕ�g�e2�hI^>ݕ�ӡV�4��}3�Uҗ;�0(�)�����W9��������Kv^���@0���O,�n�ov�ǐ��c���̬0bc�2R��� &� [)/�#)!���BQ�xgbK��\��
�Jܸ4��u����eVX�cuֺ�Ǧ'�o�rE�B�K��# ��
��Mk%
�LI�{V]�B��<��C����v��	̌tj��6-�o��-j�],+�<V��3W�/1�m����m|#�߼��W��؂ec���,��������@b�%Q��(Y? 8��@�eC����]�&/��`hA��0d���������.����z���LD�sfB�Ě��4�����&�ka�K]�u�J�$�Pf��
�9���q^a� Y�U�}2���5 ����C������1K!��9�ޠ���}՜��Nb�_��F,2�>�x�CMiA5sq>������Z^�"�±F7E��[�mO=Z�(WKXGj�C[���t}i#�[�����z~~���ݞAⳳꦼl����D%�����pb�?W.������'fBk��CFd�s,RC+�Ƞ�(|C�-��A�腅p�R�?�P;L.�����s���lK�N�#���e�w����1�C������|.6����&�X��2?FWR��EhG8�|�}\1�=�WF���~�D̀TB jh�����}����5���tLRjP�ԧj��e����#:ȟ6����7��U�@[Q&sm��0��2`��W��>�v3K-��3&��d�J��錕��	�6w�S��ËA��n�a�� ��rS&}�@}�z%�B��V��@y�g]$��eo����%5+�
=���[��5b�.ʱeP�c�T�5^���`3<R*�����7�0�9�g'�ya��}FLY
P잵�wr�ɻw�����d�)�#��f�R~�T��ԞX4�>��ZS�Z/��H�W{|H̏D%@��<���~eY;W2[����;Ɉ�&-
�XP���W��ܞj*o���I<�K����^���� ������>��o�gYe(J"��wp�
�f�jwSѳ!��f����� H��076�4�"V�kB�l����Ir�I�cĝR�A}`�ZC����4J��&"���C�ڥ�6�l�D�D��U
���H�͙I#��S���E|����מ�`�P|Y�qp_�R���FC03��D�)�\w�_��v�K�a�2k?Z<;��&�+ V�g!c�Y�;��8���w���"(�+v�1�}N֬`�?JLB�(�"C��iN���)\T����2�v"�ݦ��P��L���ؼ�xt-1�n���е��0�����}�`7/1N�V�6J}bs3-�CT][��8l�,i`Oo� �K���Ayv���ѺaI>��i��C�X�	�o�7ؼ3��"S�b�L�2����t�.��gJ�b�<{�[$�/����!�+K,*D��"n^�J�8@v���m*��M����(���C�$n�����gBP�����5��e�4X�wE�����htG�m��V�M����QA�:�f#�p��";ԫ� <�X.g:2@�Sru�xc�}f�Q�u���,g�=]������p$9��؁�{
�� Ya��4��*y<f�>G��G�r���F7ȰB�u+���o��bU{&k��g��V�MO�tr��<O"�%��|=R��H1Hs|��A��N�^��5�9ur����}\�Pqy2��#���_�#c�c�j_˾փg���|�u���
�����P�P��-*�¢Jd�S]��0���F�����ǳE�پ�n�v���{���=�������	�UD'Ռ�F�A�	��p����Y���,��2����JUe��:�~JB�O6b�z�嶔9
[IeF 	D�G�^8D�����Vl�n���iV��",��/���d����Q$�q�����}�-?~Ztc�Û�Ik�/e|�K;��ؿ�.�K�hU�~FQ���~D�E��us�=��������z���sI�`�T �C6V��c�U��1>^�SЂ�<�**��M�̚.����l�-�|�K��d�>$$͟=��p�����/�)9 ���3�Z]ۄ�}̨LA�f�a`9[AvC��d(��װ|ã:���~�����	���8 ���ºeQ���!��/�\��eY����j���9�Ũm����e�[T��k*�*f�o��O?_䝟�;"o���|*�h���$H!/�`@E���c�]c	$����3��e[~Pl(�
M��Qe�6;ǗWJ����_��w�}�B�^
,3?Y1�T���!����oK٣'������[��
$^�$¶�*�_>�s��+��3�8�="�4�����W���$o4+�O1q�og9~�5�e]�gj[����]!é4�*��F��6�PWS���፸��.��'�0���*:�[��؛�W
�����˵GJ�Ʊ��o6l*p_�d��L�=�����ͩ�����J���jZ��]ͯd>%�h��.A�b�}vU5�ba�� bċڌ�5򙞿w�܍:���d���%�Rx6^��?�:r�3�֢��1���w������K]G�"0x�]T�dH�1z��^�aJ�z-�,#q̷�L�)o��G^�ӈ� ��P�"��G?@h,ARc�[^X�8MS�D�Ë�w�!���C����4zh�\���CX��X����dmmo�R����80?� �j0��9CAF�T�`N���'K��;�s�rO��	Ȍ���*���H�����;�����#��M��P���l�{��������ǯ7�� ��`0~�9�2w6�Q�� |S��O�Y���(��زd���Fo'\���K��%
�������oN���W'�����5 goӎ�/MHL�׭�)D���|��S� b�(ȥ��.U� G�C��� K���[��
;��ޟR�����%לJ֙Ć�)d:�[E9xg�j����
{������1�L�X#K�U��+������O�[��8��Z�R*���Y.�@�Ψ��g�P���r��l�^`E��h:!�E�(|��^b���R�q6�$\"�@<�[K�wiᄩ��Tntv�_��p�v����2e��oȐ������M��|)�5�q���=c�r�w�"oG�,Y*3��b���{2p�	3kZG���XS����sKdX��ǟm�N��lvo��^T{ie��ʳ�so�g�|��˿J��=�_�	���[_�G�-��3^b�`�O�PDi~�q+�QĴ�3�}�
����>Y)|k�U���t�0�9�q��]���^#�8�[���fh�7(�)��˳_��^�ٛ-�P=��1�
E��Uώ~����!�g�O�Y9ꎞp��8�A#�����Zk�|��K��B�+0���������zZݧC ���~�9bM�&���&a{4�ŭ��U
�GB�]K7�������\txGD���N;,Re���Gb�\���}�3� C�3I`Ē#���;�6e��u���Q��������`���WP4>���~�{�v�r �����m�0��Ws)K�_��i�q�#�q�Fo�49�H����}�C�Y�ȢA?ǒD�5t��SN���<Y�`J��C��h������:���LQB뾁m
�.`f�0�!~�϶P������C7�����J��b�Fg�*������	������o�f��*p��P9����،��k[��L�>z)�1�
��tC��4��8�������Ku �0 �H�~�����k�S�n�B��L):���%�������
����f~ܠyi��7��cA/Vˤ��c��Ꚋ��i{6rz�"*25;b�k�2�D�B��/KDH+cv@�/C͗H8)&�<�!�!�ۍ�z&��A6����+h��n�e��I��^c��t`B!�.�|^�~��&����:�����p]8l�q�}�B ��@��2:(��8�����i�����4W&�w��Ei�	z��������%��2�6�73_h�=�V70�����]㙧n�5����#�"��)�sb�C=���-pK�Ƃ�����3��F-�͸}����� Т�]�Lʻ�b��)���Ҍ�#ŵ�$�����Ku�廳�B
\v=�0�*����i��9��X2r��,0M�yKkp*��ȏ:�^�
Y!=����A��J�Gs��ג�G���{����Mb�#Cޒ��xj�������2��� �^$�`������H6��['���u�|Z�-�ׅwc���0������UH�8�Nd��e�[\��غ���鑶�YTʿ���6h{��N�圶�OM����ݢ���Pj5]����h����=A�;|v�#Y#�n��h�^�}c��U��3����)�>_{g�a/R�7~Lcu���`w���k�ЌQ~c����>.�<?�v�����Q>yؿb��U�#;`��c' �Z"n�o#��n���3�s4bO����D9��J:�[�M����3�8��uǅ{2��%z��a��/�#	*v�,:^vZ�Օ>���?Gh����'��h>-V���H�v��]|���=��4.�K֭.��qؾLr��g&x1hK��:@��]cJ��]8��s���>�z�����ۡ�U��swO<�*���G�_L���+�[�O����ȳ�5�2�kDXѓ�m)_�4�v+ru��AF1���K ��0%�ik�U���qť3�R0m�u��8}!�7��!�+@κP�q�X�E��\�\�J#3 �ce�)��$h%ľp`�5����;�tL�H�}��j"_i���·$G�Ο�@��	��ˆ��[Rעvʜȏ��d��<pW��.�1&N�N��7z yBeTXc��1�ؚ����"
IgR]��9��*��D��f�N��=��8���!fOc]�BW����H8�%�P�o���AsӲp~#�ʒpg��9+�Y�VQ�ټ��8��[��c1����҄/�}D�i�µ��X ƞ�le���j��U_=J�<�>=E�!3{��xΑ��	J�*#��?/Q&�W�[z���ϦJ���]�EN�K.pBy�rQ,,m�E�ʶ�CX$�����s��ca�c?����� �����S聙8�<O	�Hx���k��0G!�,B��x��7�(��̪����0��.���R6��V��`p!���yK��ڨM���W [� ��v "�r�;�)9p0V��::�2�0�M�k �V��Dz�ڊ�Eї���Rڨ�Ӵٲ[�+W��Rz>Y'��V�Y�@E�hƎ�\n7
Ql�7�2�׺�=q�v�yYlr����X7���Gu������,z>�:$="��2�~��'_�B43�AT}c���4/��}�Tv�хd�\�HqM-̨���b��r�^(�\N.׹�~IXg� �������9�@�	�y7�صvτ�D׆:�����	Zeb5$h� нH���B�h7:w5e+��Po}T��g������~��@���~r2�"k�NAb��˫�ԍ��������3Z�A�V/�H���s0��(T&νU�w�!�N)���_58)��#-���6F�6���A��+����3u�6{6���E�`�d���U��A�Gr��Db�۲�$ݶs��L-���:���[Zxh��i��U>Yc�Pܗ�@��f]�]�^��ɶn��(���pì���L�T=M���d����>Ԙ�Q�|�[���x�A��N��kV"7����!��$���,aT��+�Ι:���akr��Z�ڀ����5WJ�T��_n�	��k�8$;��h9&q�̏u��A+	%w*/�J@��O.X�tࡎ�f���Y�\8U��e&YÔ��A�����VU��<;{$|xB��.&�D�AB�������gf��!#_��\�t���o��� ����;�2	_�RPt���)�Df]�aP~��dJڵ_�)(D�3�u]����h���|P'V/\��q������!t��@�8�/6FqQ���0.� *��i�#:�-å����!��hJ��W��Y	�;����3&C��(�Z�M��QH�|�BO���75�h���C>M�?dN��ŗ9z:��6���!����0�Mοꑲ}ƻړHW���ϒc8��ְ.QO���:�r���F���p��I��Rp��ʽ�XVY�ؑs��M����2,�	���d6e�%0w)�'�D�a?�F���J����Wd
�� ��.��fy�m�<DJ��\i����m�.cP���'��+4����+����F�,u`m	|�TzPd�����5|�uX�u6�w��'�FE�))Ds�@�(Ⱥֿ�Raw�R�r�Z�@����r�����S�f<�lR%����ta���k{t/�iY��M�1<vR�5����_���z�@�I�i|�J��ǫYZ��<�pո0���<G���q�/�ʬ`?A�����8�����m��J�����wU��;D��?���e���<������6��K�,�Q����Wh���d�:��(?!"q��Dv�Ql<A�0�Ēo�K�@O����i�2��9�Z�8lQ(w��Q��(A2ʧ���ũq��,K�?x����牓y��%�C�{_>`�#e�ߣ��q��<G\���ښJ�l��Ǭ�N�nŎg3ۀeS��6��?���]�P�tnw�i��޺����a>�A�h�|���W���v�/P��/�.�X���Lއ�{3��C�l=G�-�Mg�0��4�j
~cDO�i��c�:�V�ޮh��gl]�ebk�_~ȫ?EY&3w�����m��(�gS��SȕאEy�d��ўr���a�
úO�`,��nO��8����caR��m���b,L*Liq�Ќ��am`-�է��e޶$��� �p��0�8�y��C�q~��l9���b�����K�ѐ��b�"��{��s������Z�E[�͌m��+2HW�`_�'l��h���M*�D$��-`�ۣY-S�m}�ő������ϖ�)�uL�������n6�Y9����ɤ�g�KRi��PRj�8�+,�]�?S?P=͎���Sz2�~#��mV6���ك|kD�1�M�ެ�xO�Y�$���5Z�Z�y�
RQߥ@IF��Ӟ�o1���"���R]����6������7�{?��%Ŀn�Xc�$�w�6�Y���w���y�]�=�u����>�z<���
��`�3Pߕp�³}8�'�<jlH�N�������Ū�=̗��G��9��;׼�Y��:����wѺ�Yq����>le�*O�^��ML
��PK䎬��G�����y���(Bg.Sˆ�T�ЖІ>�>83�f�U����Z�Jv�Nޕ�"������Sl)ر�@��������#&�tR�&���m!P�=ͼ�d^�ҍ&~�r���P��o\�5�ex�ϲn+;�3}��E^o�ʇ_DG�D�����
���'' ��U"�����Y95W��ݬ%(a�O�����ٔ�s�m�A�V\r�qiid�l�������j	K [8�;�3��O�����,�X\�3
&ME��
��͊zg]^T��i�%��2����t� 9���b��kW��쾪6T& Wr��L���o�#�RSU�Ȏ�J�c�E(x�ύ��'�\�=��ֆ�@@�hA 0*k.bb`V�q�7;�\yXd˜���ln!Z/x�`$�Rr�����k�e��BWs=+�&^���\���_�a�13���C~k�^��/���O�A�'B�� .r�MO�y#��?�h(�Y"�'��J�h�J�'1��V���kn"v��/G��<&�e	�Zhk"��6�Ĉ=[��>4LG�}�Ŗ�A2�ۜ?PT\�W� �P�8~�������$$o^U:\��0�����Wu��d��=�k=�\>Lu˪N���耈�^q�����`M���:t�{�}�A�Sb6�#�7�ͭ�
��l��U��]�(��yE�9f��@�H�1E���n�J�Z���xF��	D��C=:[�n6�:�4��Q�����I}�W;z���-���"[��5?��j^"�Q�j�*T(wi--#L�;��(����p���u��16
[��KY�l�&����cY$�%#�͔��hjL���gRK
���*�_x��Y�Gގ�z�=J�P�Z:�n�1Zp]B�Z���71���T� CQ��h�D��}������Mr?�Ɍ^���{Vr{��u�4���Q'��aQ:��\�ޗ��@v��C\��vt#�����l��x $�`��Y����%tN���TV��SL��j��߰�t�n�Uxc�N7Hh�����4F�j=nv��Wy�N,M����z��TW���%�YO�*"��3�Ykjl9�b@5Kޢ"r��H���F�uw8�&��3>��.q���hOj�Q��*�<朎�Q�q�.Xa=h/����q{U��Y��l��~��Tp�Є�Y��m�%U�CV�do�+�³.��	,��Nc3"hƻB2=���~-|�/��:����QA�i�K��RG9��>�蚝$%�C�+d�LVr��f���h������F�����{7]*�4F�A������Ѳш�'*МҰEo�wl�-5
�6.o2g�kH���A�)#wQ#j�"S|�?gw)����8斮Թ���˶�wi4��G�Z��N`�q�M� �> ��_$�I�^�`�z}֔ Qj�&�٫B�I���zwl\���a__�ّ��
K�}�W��<�~4"�3�zc�t$O�$޶��L�E%���ږ�3�y��E0��KB�1�����'�I6s������]��}���/ő㯬��m,�=���C�(b�L�����9i��L���XY���U�T��׽�x=P�"��oW3&��ߌ���>�f��͝aV�s	��z�9��mi����?��['�D�'Af�.D�� ����!�X$�>�|��%�kS�ph�wH��Jx�6O'���7~*1V��h�����XJ�@��ΰ.h�'b�to�� {�����?#���x�is�K,"9(���5��"_�a���Rx��
��7�Lo:��tc���O`>Z;�������J`��.�&�_�h*�]�G���w:C��h)�bZ���0�K2���-K�:���� �T=Xɇ��>Pz�?�;:X���s��t̿8m)t�{�q��v <���p�Vi\'ҵR�-��
ܢ���,��z�:o=C�}����H�=�Ͼ�ͯ�����W>��?S{�6����r�~���5�p���v*�l�+��ڠ񗱠����Qh�"�[�EW�9 �Hh$E�X�Yt��2�\�΍��7[����ohtA���xrUWu� �a��n�Pk���5
�T����M�Wp���,�v��k[Vߧڇ@�&�鸓M����Kj��gEp̴������+VpR�'s�s۝.����U��	�>���<���1Jb!�(Y�E׼��f�X�v�4TGH��[:��^�Zˍ-Wj��]/���]
Qg�	v<�≦ɱ�xܾZ���!*6���Bګ�TZ�S��{o��F��C���4h0Agy�"�ɟh����nQ���f�1궓{�l���N�������|�F�-�(�Ze��0?�}i���������_�0[���xv5�ܘ�_z��O�~��@\w<������O�,P�'#�#	�����ob���[�R(�oqٟ̾��<� |����"'�j����Y���js�U�Գ���
�A��N��0�~ZB����0-��()�%Y����4n�/�؏%O��{?Y�W_�x4�F��k6?�U�앍�o��!Fb�.EK��g�p	lD����xX�6�n������fTj�5[�j!�w�8:�ޙ�vV�%�S�5Rs��/N�f_�O��n��W9�G�ƙy�Hp�9n�Mɑ�e��� �2���"ޭy���������<��>a�	�ċa'�_��u]�Mb$���W=*��:�)Y��2��[��u���B��>'�(�@�9	W�Z�+��N�i�a�t�U8ʔ	�UJE����D:�9=�('F��%��X��u���Iѐ[;�Ǯ�Zc);d�������I���J���ʹ*j��!� ��ohN hl<ћ���di�l�pG���.�����DB��|
]A*��}m��m*(
�?���T�dX�"�ПA2�;�-�� S��r2��������ʤ�V��=��O� Xo�H�m��Ț����y'�3��Êў��o��k�$e�%�d���Z�x0� &����2��e�U ?�V�ij>�y�y��Qe�9�@��@��� k�����˜�3�ѣ���������E�sG۬���K�w����PV�;J7ox��P��0�J-�ñ�p�5��H��~{;�;;^E-�֕�w���~��bO8˶�"��+�_��2���Jʃד6e$E��L��,���2U� U�>�g�K��P8��	՜��oQ�W"���R�m�n8[N�?V}�j^�玼d���.Ż����@�B��3͇O��(
;��&4SA�}&�F��}*�Ӑ~i�F�x����ͷ�zU��Ga��,�C�='[V�*&�g���٫��࢑���~BJ�w\Lo��[S;pI�&II��%H��	=	U,���IĺJBڬ�+δ,y����ta/��ӐU�W�0���s��`)��w-+�v�L�l?�Z�~�b}W�}>���R���B���K|����Rf�,3�'t�v�5���xߵd�r�������w��&��d�I(n�߬�����!����κs�C�Bo�u`�Zm-��o�u)6����X>��9������xh
;HzpxGn&�1���T��'��:g�R-K��U�<��a��I�*���;��[f����1y�ũM�B��|� �L-6(���>[��	=zCl�w�=OںJ��ނ�P��p��s�)�GJ���,����ru���<%�9n��/�Q��ǡӻa����?�٬l��t��.��T��\L�֏j��6@>�`�C�i(Y1���i�O� �J6��*w�'pҤ���>*��c���ha"���Nk?Tw'��q8��)\1=���x|B��S�a�"�5}��#��App5T�lK�(����d{�D�4f��E�jr��cۑ��i�!�,˴D�+Tbp�F�0��u��� <��j�&I��2e�VA�R���v(.�fA����J��������:� D��MxT�G���S�	ˉ��l�������I�9��BLԽ)�	 1O��L���v>ń2P��9�����So�|�����v�T���+rN^̞�_JY#懜��D���^Mٮ���S
�KVx�1��S�ث�=�C�9�R�6��v4,��Ό�@ ���H����xG ��^sq�F�� ��T����C����!�CJEb�ݰ�w/��r+=<�W,�[7x������]�Y?+@ޅ#���[��u��T�����-�fMۦNl�>i:#$�<hì�)?Mw��~����tL%���ٲ�X��F0m�j��hp�u�\R}]�|�a:���M+��I�7ҚD�I��NW����?�J�Z��Y�팎"��y�}�1�R��[e�G��S�|h]aM�J����U ��Z����?�����)
Z9ba���&j�G�t3�'�a@�R����"��e֗x�^�7 �<�Ө�����zw���1ȍ���A&�b�́�͹� X�`w^Nm�R	*w���]~H��cp��=���U�=����qdZY��z��۸7F�g�7G��;�~�}��e�������I��p="R�n��	�s=**�?v��I����_	�V�TI��lzeRR��C(�'�1���۲�TM���Ѽ*�?:�C�:��˝d�����p8��j\�En#�Q+�IԊE���+~kj��G�8��c�`g����(E`���:���9+��9�����)�jd(���nt����|�ȡaz�WAPbw�l�[�	C��x@��� �-�L?[h��"*G��`��~�pxVE�5I��WW�V!C��W��n��)�ؠ�9Z;�X(�(��zo��^'�T+��;M���MS1Q �ޤ�Dc��k���$p��GԟmO����V�B������o�Z�H��l�=���(���3~E��!��h����}���\7�n4�И����P�HlʉD��8gCz�S�0�z�5{�K/�#F���@�|�a�F�����n�&m�?�"���g���EH���q-
:�wTI�s�
����'`^��a�:�i{{,y�m`zh�(1�4�H�&�~���w�Jt!(�*[�L��#H8pl4F�K����lv�-�d���kE,a�0*$M�a¢x2�1�oW�fմ�lC����V�/���c_�U����"����og"�.�3�v� n��� �\t�28��o@|S�,�q�Q$�R/}V=� �&��B�����Y%��G�M�*�_����cx��ņxEu�B�QWd��K��Y����GMM�8%��Mo6p�&1�r�-jw^bV:{T�V���\V�vn���ť�7���G �O#.	8�nu ��6 a�QDYs�Pgǜ�8*4\�D\lF��5��h�9A�ǰ� ��r���j����^}�JŦ��z��ʢ��LV����h-4�C��"���A��Mv	��o<�vB>��X{���"����`��X' ����S#���X���gOۢ-a���M�/�#��($ɹc|����,��Qᜱ�Y�sJN�]���z�\�u۰@���ѫ�eo�ʙ��Y��<�~�32��6�0��)�MsX`D 6��X4v�����c�+߳B�U����/�o�s������D:����"��%
ӯ� 	kD���Ah�(��� %�!o�`������L`+��mn"�t"��_"�\$L��90<�����}9�On��� yYBh��_��[��`�#�A2McD �S
���&ZXݸSX��y@����^�8vgӆ H91����5K|�L�x���^m�	�u������u�n��a���+�. u� rЉ�r ����+��e�ל�n z䔡��D�%JyFS˥ۘ�)��?��ov�±9�j�s�t8�1�D��y�)�0�Zib���uQf�'@�_K	�K�6.��.W��2���Dr�On+�y�͸�C�m��=Ki�z�����/��a�VM�xP�"mqŠ+�Dd�|��Vcw��2̶�&yuz���|s'��(�=ڈ���f�^5X!�R�z{C+d��:B���`�U��Q��3�[��?�i�i��D�U?��o�e���*����w_��I<�X�,-�����<{����hk�T����L�5���A<�8���Sq]V|��5���Tm-r���iH��XD��R2��-����	W��N-1Ng+x��k�K�LBa��@�IPdz��d��`�6�s�Fh�]p"9rr�Mr�G�E��d�9�y&Z|�]�`�	p󲗲��\�g�s����:���>(�̅�����ԐY�v��:�C*�=b�}KR��Yً�4B�z�@"->���N�F��W�V��B7���Л�p|UbsʏX#�cDme�)+P�^�C�x*!�i�����l�0Ko��y���~5����e�=�u��;�V��H��^ƅ�?�Hy=v�P����X�N���)��.*�o���R/�=�M֛wF�XÌGlWh�04�;�b)�)�喏�2p!8�YUE|Zd�u Z!�D���g�w��v���w[g{j��G�ȕ�jѫ�9*Xz�0��v�f�Ϋě��ɹ��E%������Ѕ¹ ��fZ
�p�������PT��H#�x݆�ga���-�����r��o|��']��򽓾�(IGF,�n��|��ke�woVoC�9R�	��v&�����_p��Y�v�w��%�ͤ,�Vѣ\q�x;���> �7�'-������R��M�(�� ��e���4_����!�}���X���z�!�ɫ�tn�6�� �~5����?�t*~��-9�a1�*0�Fb��{'��|��*���,ޯ��K;���e:��@��ݧ�5�t�=�?`���Ϊ,6u�r>��Rð�ƣ6���҇�o�X#S~d3u8�=�k����<��p��%�T5=��'��pTU�y(u�ƥL\�X��'��7��m�F(��y.c���$��A��E�!�Y�q�7霨�~�Z
�-�`�����}��l���Tr���bV͖��ͮ����{�)�z�M;m/2��'T��_�-�}�>�r�}��T�Z�f}�C(b@X�ᠯ�����[o;.��hy7nW�j��+�%�}�^xW��T�Į/��sO՜�J�ɺ���-��������z�ֳ�*��,�1���}l�@K��hB��I,qh���g��|l���e��!�`�.����P�
i�0��״��.|
�`����x����*�M��q�Lz�m	�oM "�d;�L�S��X:�b��W{9��m�%R�W�f�����p�~j��ʻ`6��Ma,JHx(Eb��
���J([C�,r��>9�#ll���������q�bDP��%ߕ	ڃi�1�xvc�B>{n����E�j��e\�G0�7��}̑>�����wC_ڷ�͋v,G��]^�kk⾗�<����08��X<�2:&��"w�?��O:��ER��u3�*C2�b{���b����ݍ����'&PX{*��3���}�%A6�}#]b<�鎅~�(��"_�_�lɠ3����/����ލ��G��/h�?�Ͷ9rJ@R�hҳ0��:c{�[�sߥ��h�5BH��c�+Z{��E�mp�r�d4��]�Lk�<.��������{SF��y�0h4����z�[��o�w�|4�x��^�@rjR�	�7�/���hf'��j盤��j�d�-�� �l���þ�|f�����BQ)�K�9�_4
���%Ƅ�Ba��B�~��|6����Uְìv_N�Eѧ��QeyS��(g1�,�[}�a�`��c<B#�+�(�5��)�ȶ������	���<A�d�v�s��HZZ�ܐ��f�oS�=9�s�{��1~q�=@�N[�����Z���[xC&��?G V����y=���q랆O����=H���0;�� hu���r�Q$����3��4�*�л�t?7*�GBL(� �N]�T���Ϗ����&f���q�����_�&�
��w��wrp���y��jҪ|m<����曠o�l��m��VU]��L�>ϸC  �h��~��������܄`^J���e�ܦ�^n����ϿY^|Rd��u�׆A�v�W�=��lBn8����)0�۸����9��i����k�j�yB�G��po�z�;�F�1�)J�q|noh[���uj9��P�,�yvo�R�a&��r�V��Z���/��O������XC0-"Zk��煞���%^�%I��+Rbŝ���O)�����Ml`Tt�㢿>�d<|*j��_1__7�VA�br�3���(NT{
�� ���jrXkW��/����EMs�]
e�Ȥ8;pe��@��(��~�M�|��н�?�G��CO�������v�=lV����y�k���OB��Hz��MZ���Mޜ�>���W3)�2�}o-Vw���	lf���X�F�Կ���N���D�*㧪�}��4�|:��_ʗ�q^nN��Nt{wf
he=2�L�CD�	���?��0�V�H$��t���$өM�ڧ�0�_�[����L|�.b��~�cE���P�E��<Ӣ�[�CT�i���=����9{Lg`&l�� �|gW���M�����g=�ؙ����zu`�Ö�K��Ҿ�4��Mp��L�ɼd{vXp� �h�^ZTH3R�����ˈ9��s@�ND"�sPFn�Y���Z���rte/��q��G����!��Oi4�KְW!�r�

��ð�n��^0cp��#ɓ.w,�]��
��4��Q���x��Bw�+��Dɑ����@��f�@�/K+�z��(Rl	[1]}0:E\�FR�uv@e����M�sJ�l�hg@�>�u�|(�������i�N��|�X�b�x�X�BX�Zƥ��p�8�`��]��h��{W�C�y!7Y�� ��g����쵅�o�dI�n�{Wv\ Vn�!ܮ�l� ��9��xJ7s#�<4}�w\t��=֠D�n ��� e{Z�������?��ǾT�d0A;N��w���I{\��*[?Hˉ�'yR@m��{$�r�Adڙl`A�>�ٶ�(1��^2aE��`ela�c�~̂���*�0��g�JQ=K��iy,r��p�Vp��	���������\�^�fⳜ�J�ͦ�E{~���=;jr�F��c3���q�E��Y�J1"�d���K�i�" �ܺ��X�q�K�s!�y��L��(,Er�W�D��jZO�*�L�~�ȴ�*�1�5�;�u �Ǜh�C���t
\tOn����ڮf��!�kA�G]�}ʆi���L �c�z���U:�T�g�Q��d����!�+Ir�g�/^���E�L�B������{���'��Fo����B�j��Y�
�+�gL�ei����l���	BR�l_iʃtOB_��׺8\�m�h�J#��7�RAbWgŐz��!u��&!�!�F�9[_�����O	���zK�e��O-��!�9���ޱ�M��tKo��^8O� ��;�����0�ZR�+�H7`�R���2�����{,�P�q�S��������B_��׎z'�cZFK��Ͷ�6Ǉ_H������F�i���y�U�H|�&��RHT�r�A���f��suѣ(�2KJ�FP�J���9�s��߇F��9���P���l�M�Q�`������~~���\&,��i2�N{(�11���<��(5�Q$xx9�Ix�u�JU*=55U���,���M� ��/=���kKG���hA����]������D~ hG�̿3�:��XEd�=4Fa+��V���M����1H]+W@t��bD�5�!94��r��5�F޿��s�,���l��o]ر�c����
`{j�������i�ou�hcD]Cr��_C*ƾ_��<�.m��'�b*���[TR4,�`�s�h-�y��v<�ެ*xJ'[j��7RX�C���E$�gLb��4��>��4�@44�A�$m]&�'>7�ޚ�_4&�y��ś��ծ�k�GV�<�kl%'ѿ���7� ʺ��UP�Z�;N��:0�����7�:��Ga�,��� �=Y�1g.�^����8@}�"�G���=�^B&��cv�
`�ь���:ߦ �� wY*��	I����#4��&�u^�Oǵ���-�89�U��덼S�~��:4[�.�`�۴�¡�ɍ� x��4����&�*��@�K�l���]I�
�1��ySP�H�ː�Α"�@��r���~������;����uck�z�<��6��oia��Ǯ_�� ����j<�� é�kF���@1�֢�������,t�z:d�Sj��uʵ��i�Y���@�?��y���1���>�C����t_p�������i$�������*�3��db�)[�X���fI�y�J��|#�'0��19GL��)^|i�^	�K�~�2�kg{�J���%�V���nDC ��<�N���4w ��vH���1lVTvk��V{dY�[� ����CY��x���)���^�mZC�2��I1J���Xq�r�)��A��o���`�#�G��������ҿ���8�#�_o�B�K�&�j���r��f�Y|�%�f��>�p��GQY��֬�Y�h��As�b>
�χ8��@��O}�`@�졙���]�oMk��u����.���!�}D_��4L`�@F-�R�����cѰh��b��}}\p������#K>D��J�J>ѫ�Āh�К�on	T�g���r�&�� � ���6�׆}��^*�푎��3g�=H��0�?낭��*���Bl�p�JY^�/�~�������Ȣ�m�Sg����,���b��U��4�=ɩ��E-������o��̜�g�\���0�u6����L������T��Vd�8���P5��bߤ�N��ٍΈ3���):��@r��B��&5��ϙ���-��|ڃ�S;o;A��,_����H���30T����<�(f��,`A���١�JeU��wW��mA��8Ǜ�����������D5�:��i2:��Y�B[��Ko�oZ���{9��W3R�+��$%��[�W-f�yVQs�#�Yƪ�D3�PƄ�� M���P����g���m��! ��x��X�U�S�]c��;� �b�b����0��p̼��� �2�E�zi����<��@���޿u��+`Iߧ/V�f_� |��^��U�6���ce\���߭�o`��~y�ɂŇ��^��[:��^�W��,�jۗ���*��_�g�i!
g�(�u5�3�u���`ߪPr��~��D�惭v��7��n�@�l�Bz��D�ߤ�5I�G�Kµ)H�I݀+�䗞[��Q& ��@�V�6�7L�F3�l�>�Mx%��{6�7���]VA�C��W_Ċ�ԫ@��K��ʜ�9;Pz���Vr� =�T3V4i��:���ނ��}<��y��R/�5���U<(�D4���i�z}�?�c�d�E[.u��Šg=�^n	俢�pY�Q�1>.�ʦ#t����.������J ��qK�b�g��R	�����n)3���{�x�@_P?h�҈��K ��)�_���1���$#�$�]k̃�*��������:
�0I��k!l�D {�s_�����n�OS�ǘgT��dѧ~s�x7WG:tj(��'-��}���Ru>^	�A�^�%[.�9�zW�`�$}F%W���9�}M=� ��4�������;�ta�>m�,x��6~���dyѫ�G�w��"�����0���V�B��<�CO�����tRJ�ZF��w�c:o\S��Y�v9m�M��� ǎ�'��/Wh%
5a�90��Q�0Ѷ�O�x��]��?.<m��Mm?�,1	U1i{~�N!�>#���n�f|���O���?ɯ�Y�L��`�}���n���dUg.��U@�Mn���o��eS�UEf���!�ߠ�Y�������0|�� �Mӗ��zk絇5��t'�l�-FUk��� b�Ӹ�l�6�g|���^#,ȅ���7R�:��>p7�RJ�g�ҙ�y��1땦=p?Og�L>�|�ڦ6`�=|� �nO?�(Q,��7k��*1���������}��e����՞�,sv��ֿV�}u(2��7��;�ғ���7�T�rQ�Khw��j�O���N�?؁��R��m�N�����W�R7ˆ���n%�:����?4����ťl���Ƹ^U�ӜMl�ڳ�v�Γ����<��މ�1�
x�#�%ĵ�`C��ƊM}�wH6@*3y��Łz o�|_(?��:���|��J�͓��JR�kCko���*.�.F7.`n#��h�4���+�3�ۇ�:���.�-6M���Ep�m�UU51�fA�����^*)��~J����B{Gǜ%d�8���e��q��H�{���M���]��)3GW���US�S�E�o���&�d7�mf�n/k�?�9~Ėߘ��?��W6�ML���X�k�I�{(M�3;�M�Z+W;���Ip�p��� \6.������6Z�9pB(rD�b�ql\0i��j�鴏���RD�x�a=!�Slka�گϔ��ۇ߮Bܵ��(�H�\�tR��b��f_��:��S'�� �?H���s�F��N�x�^����ֶL���-TQ�8��	�Q�:>����uB�����=7}�ۑ�O\��)U�d�wNI.Y�K��\i�ˢ@W��(�)���|W�{#�$��EM?�Y#�B]�ؑ!��P�c���d=	-�ZNm� ����xFx�d�re���a2���X���;\H��Z�x�<�hS�#&*˥R������KV�.�e�lr"�4��Z
�����Wg�"RN�m�����ݨ���;���l�1��0��V�X҃<�c9�H+M�E��F���Z���E�������~���wg�w������� �δ��.���/�] ߼��M3��i�^��AX/cʧ �`��\�B�c%<sw�y��3�OB����N�9������m���	��� 2������w��'�&zx��d��JTD����kQ�4�3w��̓>`��1G��x
�&�]�,�~%/R�u ��w�g`[�4�5�/v6�3���o�_����}6%*�'k�;K�F�H^�%i�|%<;�����C}_����ؕ�ڙ@-ވ���fD8(�;�eO7&Q՞��K�z4����`��k7�^�Hc��h[w�7hC$R�xo�5�J��ld���(�h�8�h��0F��IT���Uu�NX���^��KS��}���!���{X���֚��!�X<�Wr&��֤����V��K�x��:C��M��5���}{�	ldꑞC$<��
�Y^���z&�d،��(��^���`?6y��>Ia��	�@����?eG�k�s��J����նJP�����H����M����;\�Ef2�H� �~���.L��U�![�7��Bo�3(6���k���^�c�����=蓼�L���b1b�6�DpV�X��?a7���H�Q,�[y慵}R��U�=`���)���	F������#��Fn6`�_�رM��㜁�3J�b:�Z괳��>�TM�g(��㳪��bG-�5&-�=j��q���i&	�l�מ�,� �ƌ>/O6�v$GO4@�̸g�#��m~mD��yB�T9�e�:���T3$�m�O�ꯨ�(�u��I2*��:(�G����bm�����:������k��5�w��Ƴ���K����l�o����3�F��h�a���E��(~��u
����ƴ�_�������t_����C8	?���e�����Wu$Dҋ�Қ�m�ѭ^��I�Sx*SYE�	�ڟ�1���V�F�+�S�D�f���#q�����7C��N��i}���� ��;8�������t����&�b�Z@�ǏB#���H���аz��l�� ����;d7��^�VJ5�x'��h9���qk�V���8�BV������2�����:"�>���65.�$�>�aѺ-��S+�^FUD�*�)�H�w�rk���b�y4�!���}=W�����|.3eC�2oZ�L
r-~�7�>��;4=���>[� ������J�='y����;��^���f�j&���WS����<����pY�H��BG�� �l|��t��*����/��~��
���~�x�3� ��~8�r��&FbT�T&�x�Ȓ̵I>$Ȣ@.���Ӏ��#F��F�(��3p=Xc�v��o�� ��I]&u��ko9�������D�l,����}3#�Ahubu,��U�u�s��p}U����A���4`+�dY�`�����U*�ydZjKFg ZOd,���B���F�Z�r��Vô��q�e�����X��!�I7� ���U��-N�������u�
��� ³���} B&�M���~��U�/��1gb����~��_��ڹ>ˑ
��sH���C�q��)m�,���lм�T���K#�I���:���r�Ǝo���Ҵcڢ��!�!�_�� Ǯ4F�q� �:I�]y2��V�=@�FEJXr�4�ı�K|����i�Z�M�ƕ�����b�H��l�g�o�c${�CF�1���<&"Q&ӄ��>�&;3�pA�����k,s9 \<�J�x���	�Kr�{�[#�y�#��q��/ގm��F ���_\qW,㌁�>�I�`s��>	)�!ty�Q���v�V.yJ��yg�须��<"�y�G��@Nzhha2�-B'2�����'��}W��0������ȾX�S�H$.�#x�r�	�J�8i��W�z�����,�����=M%��bg�3K�M��%<� 뛁{E�� C³��c��y9)�4,y��AKl�K���t����.��j~��D��MM�AG҄�#�8�MW��~O�|\�
�I��!҄d��1l�J��ǳUI�/"E�"�)����wK�(.\���}i�i�e�6������IS�N�â�>�c㠮P��Pl���"*���/�o����e�q[f� u_�Q�ʱ��כL�}_�q�O��Q�FO�Nfr����
�G:KP�F��8#=n:;ޜ(5>M�O��;���d������ӷ{s��r�G�Y������w�PPc9z{h���<��"~�=wa�ofɜ�������Sn�rL���ɑ
�i���3�¹٬Z��ۺX������&�d���b�Q�"p�k�Uv+~~P?��u��B�w�ή�[7�L���M���X���F�������=�0pd�$��x�m��Zc��k��Ðj��dde&T<�G<����X-�%��QW-������`�/Vys�[@��LQ(��>�4����3m ��BĞMa�I�[Do@� ����� ���ǁN�H)��;�L���)EY>�.��Q����X@��w��h2�t�ɂ�*^��k�7���\����x��b�`�[v �����z�-��L�?!�������e���"vg�ڡ�)6�i������>l�x��W=%��ۿy���-G�H�ȵ��o-L��%~x��jJ��7D�yɸ�d{'9r��0��zC		ߑt����-5d�8�|��-�_ �S	����s2�⧉ ���I����4��c�Aq�;�:Wu�Bm�n ��G맺�/��bX�ِ%h�f��g����^@|���� �]��gTk
:�t�,��i�0�=0L�iG`�o���E��+��d��ۃ��8cz�l�k<��1������ŉ�\��`���:UG���<��7�y-�"ǊP���qc�D��c��-��K|�5Mf��7O���n�m�O/�?�4�C�J�V�.Ӣ�P�2"H����g�q�q����g��w"�k�Ko�k�y�1�`֬�")ߔ�gE2BhE��{��X�g�ۚ�Uus�����n_b��)���}�Ӟ�����*W=,�#R>_��0�O��y�T�7A�V��Y���΋���~���g�iV`�gZ�3e��e((������Nz��d_�[������BMLm&.�����N2PK�p�'�zEw���mF4��;���#r�S�OՅ����[���;"��\�_{���E ʞ�o��c�z\��W0��ns8L�S.obNŀK�7��{���UJz9~ ��,���g��-�u=�I!�w�j�4��iI�"��i�����ayO��K��i�׃��ĩ�fӃ� �Fa�*�G�<v+8K�1��S�#z ���j/Y�ɹn���:NF����UgLfo��Y�ӲS��E��o���&ϻC��p?��"!��U'G�&�&}�瞩��H���ʗq?�Wf�o��ݝ�=[Rk�N�4:�Y�_�*AV��Z�e��H}��p?ծ"� {�7#AZL�\���0�er���eF���=͗����0���;��5���kf��|���S�e{� �UO��f��=��h�{
7$}�W@�!xgtž�#t>�0���g��d�?x"�@Z���@���`�w/�EH�#�ݺ"�J��F����L��R~h����u���1���*���>O�����̷�1�~��$7hXvw%:
�u�u�,g�!+ld�"4B��D9���Y�����/m��X��v�?6a�!�ǖa�:Oth�0%5V��M��%!Z~�p�uѬ�D\�-�%���K6+ND^��⹁qɱ+�Ͽ��9���x�j�+�t�#L��DIg�L�aG].��=�'r�WY�f�Ԙ/a�<̈��$8%�a�9d�pn���Zt#�D�E��c����5����%wH'���C�&%��v�d�$<9���/����y��8����z̄,o��`�+�-���l�S��L�Ц�<��!^�#�r�A��8*~a�1��ǉ�X���:�'��nw�V��gD�'W��16�&	$��S����<s6yXZ?��@|#�|�:��"'I������Թs��M�d1�4��\!��h��Ja����ty��lnֻs����5;MɊ˚�]��`X��[g�| ��"�e�kq4��&�N�,\Å/r���TN � ��D{����_�3`X�P,޻�S�D:6��i(<M�|�pR&�F�A�����ʴș��r�C~���V��΁�O�v���Mg��rV��դ�.�m5��fb��SB�;�و ��7>�\�������*��h�9�����[E��R�znQ������t+��DK>��)��ԅ�����h��et
�@*��2�Ɓ@��A]�a�[8�E_�
rZ���8Sż�F�~��-V�#�%[D�GYB�AG���*C��8��4�y�>�t��q�M�k��u��M�B��U�Ӧ�-lMuZ����\�f4u�
�U���D|�������s�+"�f�8���HL��x��t�.��{����u�P����&	j���]Ho�4Qnr#=6����[W�h��OkV���a�Z��Ȫ�q�U��?.��b�}������3m�kJ �7-�i�;��+�0�bן�,���G#r{�"���p�ݸ�zڞv�9�Y�����uz*d-�>����#��DM�>��i�6�G��zz;�<FpM�:FX`��\r�
9ˁ���٠��j`y*�2��"To��x�g),�l��b���%����I2��8+ ����_d��۪��3������~�D�1a��S�^����F����e�$5�9;C
*v��V/�kQ��
M-S�NDZ��:B�rH�<L��W�
k)�ܐ�mY�V���>9�n{f��k�[��)C<����F#ct�� �����0Z��|B(B���@�\�aHh�|p �j7$
U5�3�:zvd�
v�e��Ɇ��aaM���US�����N�����=T��I�'��Mڊ�\y����s�� �t��H�ͽ\a���q�|E~v��ki��ƘhG2��F�F�d7i��g�
�M�n���h;�%��W��i�P[�����&\(��K)#Kɏcx�w�K!RQEoL%F���F-D�"���n��E���fSY<sޜ�A�vm�I"��������c}�,2�"�)P5F���F�M�C�`����XTN]���j��&�}�����&���$�Ř=�Ų2�$�J�2ۄ�wh�E�z�H=��
E�5���j*��\Y%k��z�ņ�8m�hT^�ld�����W��_�8�;�`aʜL��J��`���\t��Y����%�߮<�>	�ގ6�?y��k�h�^W��&���Z|+��c�Gu�W
&o�F+]�!%vbc��a#��t!���\8�{�v*U��W�R���xl��	�M��/�F� 7�Hդ�`H�йDc��]Rw�q�-2n#y���Fu2g���B�F�R��W�P
s��
4!���T/)��Pc�&$�X������%���9������{�>G��ϻ�x8"v�zi*�� �"<\h��g�
�A6~g�nu3,�r�s�RBS/V_Y��zo� ��Q��l���2�5�)��+��������=N�'.ߞ�vj.z����|��kgw�5�O���=;�7M�	�����D_V����	��x=���z�e���S��ﱢ�x���q���6x� �׻K۵.q��kj�U�u�E�]q9n������r��°��zb�,o}!�d��YuL�|��(�1W��b�f9�%�:>��d��N��ʃ���G�Ύ�F�1x�r�s��aO᥋B�6r1l6ؙL�����<y,��;��T0�/������Jt�X���CE�QMy�Y]���9t;N+DF�IKX�Wc\&�_F~�F��t�����#���åPIqL;,8Hc�5���y$��2{�*��ٲ���c'�EQ� ��}Gv@��\)8�葢�͔����s����������1��i\����cc2�:<Re8�du.:T�्��3LȢ)�%_ݍ��iT`Yտ8�����E��������G%	z�K�d��)����rpT*f�t�EP��c��t�,�|������A��x�3@ڶì�ht9M�_�>$�HQtT��/*�u�e�-d7���~HZ�yN�x}<�b��+���:�~c�A8����r�a���QĞάL��d')�>���L�b3Sd�щr�+�LC��`�f�s>K.�jR��@��S��l���v� !��Õd�]i�_�N�`��%�ab9J!zv�t�#ѱ�g�� ���3Տ��O�F���գ��GH3�4�%X��n�� xVwc��'��� (�^���-45][�R�ĵF6���H�ǸəfI%?�`{y����}�|�4�,��q~����3�O�Q8;ղ�ĘqH8�.���������Nm����|���
��m�ƇCC�?�X,�v�]�}9jZL�m͗��OZ�W#��UGxz/C}!'|ԅ؜�P���65E�Vx���H��qt?>��f�\=f}M�u�r&�9N60U�%@O�Ye$�.v�sƧ����_,3q �aW_�{���4q��V�s_��(����̴�"݉lB"�}.%B��-�W##��o��#�5����n0,* SlS��N
� �<�����\�4�O�rǔ&�=V����
❙�����U�L/j�x�*W�`F���A��E���#���`�8,��ogG������^�a��!�x�i��X�'��7��������u�4��S4�]�U���
�$��ܺ]���e��R����ݘ�����i
Q࡙���S'��NKv�T�M���}����o;:�y�B�6YO�yܥ�`�}7�z�8��:��I�}衺3ݥ��Rnc�w.��u�����~�G�0;8�$I��0E"�I[���f&��L�c���������N̒E�9��S�
��h��ڐ��_�	#ӥ7���eI��%b�@寫�)kW��ђJ! ��nE��B�O���s<Q)�ƙ�|t��53V?7S�'#u/��-Pe^���Dȣ�\#�_���*�/7Ma��ܷ�s̔�
���r�YU&�
DKx���N�.���Їފ@g�D�x�b܃Լ'b�*5������f;7Y�Yx|g�������|K`<^Ԭ[�+��E�?G0��^��@p����A�wi��5p���l�/N<6�hv�uYf}~�d���f�GS,����Ѽsx�����E��
�9eoV�j[m�ˆ ݍ��^{����2�����Ҩhԏ�iX�=AdM�[r袎�P�*D%灧-��E[<J��[���2��$���őbX�S�f$�L���akc�䁀��cPv�<­��r����bb� s�ӳ��,
���F�2��%�h�1��5e���ܩ���/5�V�ÓzJM?�pKx��\���n�0��!G"�pƑɢ�~��T�?��AgVr�-�0i�������<���{.8*E�r��[�1��P�'=�����~�wh��|-�@c~��,Ů�<49���F}�ɜå��M��K�����r���k�W8.�?�����F�0@^?���I���/�h���s3k��bY�6H?(~/XYK�a�{Z	T!MC�U�Vj�ei���Ђ�)���R@ש̲NGT�	s�s������X�^�(�I�(���)��q�8����k��C$�+<~�Ee��/ x	],�0S'��N.~����Oa\!j����ŧ�tE��Ε}�����1S����`�A�,)]"E%%��s�;p�.�g�S�'�߳�/i��ͧ�����v����n�o,� -(`"�ƌh���=��t�"�1���ho�NuCJК�
�R��.���]�ͰN�s?����ş��Ҹ@��s옂����yU�o��$KJJ���&�T�i�n�x�P�I!<�)���X�e���9�u��h�}j�Q 7��[H�G��TY�~�$+l�|�������� �cH�����Fv����$i�PK���h�$8��.��o�X�k5�=5Sж�܆�W/���%��2�ۙxApJ���&v���j�$��3)�TP$�ϯ ����H*=��A*��}����[si�#����0�o����p��3�}S�@�{}�2���kl8���?~�G8�=�J��Sұu�W�i�[���i3��7��N���.��D6wB:YD蠱�梴�i���i��j��^�vH�|Ӕ�=3�{���y��z�js oժC�ģ��.i��+'�9�Q�)im��AW(��Bv������4��;�� �3��*p���^1��:hk/*�}M�VR J$e�JhzLK�bw�gJK4���O��F�A��_����Aqo��k�5��u�����2'<�s%���
S#;{��8:�����a��|AO�e[�~�0�
a	,��mV1Y��D�݇�u�l���%�/_s�p�u�ґ�	��υȎΩ�.[]:�ԇ%qEQx _��������O�_��cN$��r�mZ�+��x����t�gݪ�.6��O%5�E����wkMgj��a�NS=]� ����� =�ưH��@b�yi˭fo�Ϋ]�p�V�Q ��T}�ׅ�f���zL�dO4�Ha�슴�;��.�BN��k���������1E'�D�e�,����v|�<Ap�5&)�q8/�(�xSv;�A�\]�P��n�� M�U�Xq.�!>{D���+�M��&��~p㿗h^5��A��Ğ�XӚ��_T+딲��� <���\���B�v>�U���2kˤ�d�C%o< k�L�OnwY��r�<�$*a��k�ərFn�/L׼�B�R5T_��[QQ�-fs��==����j��Zgҷ@h1�9{~��$Oȶ��ˊ���&���@T��#?cr�����H���L��S�Ot3'�v�t����������x5��K���R�0�j����W#�T�h��!XgOM��P�b�>����}�9�\z$����׭�*á�<s*mP���u'e���ܧ#�R���?5�y"C��\�x*qD&��mI}�����م�A�y�7&�+�&^�ի������.�A	Ͳ�R��+��Z���ҽ�b��ʙݢԄ�a9$m�����fM%j�M&߂"���C�4_�ҩh�d���4I�R�{{$�4L%Ct�J�:`���ڛ��Z=G}*S��T� 
^����H����p�����D�T7�/Gr�&k����=N�c^��G5kn���U�Kt���7�s�s�%l�R��?#mʾh�����,�gV&�27G$a�~r7�Q�Ks��1g���*�z���7�i��'�.	Uw1�Ny���0K��.m`�]��A^5B��8:�8cڶ8�ag�rLE=�&�-> c�`��x�����������9eQ4��)s%��ZŻ�� �d>��|��ۗ_g�	+*����B�����J�>��N2�3�5B�]1+b�A���U�B�a�ʩ�=���pU�W�i{��пT���l��"��ʧ���4BM�c��;�F!~��^r�Q�Ŭ�Y�TZʥUQ������W�j׻�p�4KB�zԣ� ]u����d���gT��bX��`8��Q�ԙG���\�N��y Hp�z�L�����J�I�2q�d�$9ZX}��9\��O=	I�	򒚗�Q�U/�������[��ϛ����	�BV�6<���$v���ZT�������'�m� ��ώ#wDv��X}[�NAeȡ����I[�P��B؆��=�i���|,F�;dE.��x[,�8�U�Nf娖���8s 0���x*߹d��ô���Ni�q�7bՐ��u}�%)� +�0n�5��G_��)��P�,t���kԁ0��D��0��ݎ��	PB�>��1�OV���|��'9���q��2���47[z1�>�"m�t�ˡ9�M�f�X���g;LN�XI�w�D�(��-Z�f�Y�E�y/�6��,#�۶\u�bO�ni6�}'�Cc}^rt���4��̸Y�̤:�.F:�K����͡�s��Q%��\"~Z%@*ȇ�W���^��\�rD�(J�z£�0�؇��p혣칡ad�2��ë��l^g��i��@���������n�lV�;
8��ܧ��#��,n3�e%9~#n6��ĩL��㶊�M���z���C�1vL.��:��.��nX#B�O~E]orbD�|أޙv�t��8' ��n��#8۷Q�hUN���e�R���ͫ�P�]�6m%���'�]�G'�yc�bS���&��p�忓]�5%�pX|	����N�
�G���J���V�aCW��Ƒ��$�ൾ�U��7�N�� ưj�k�w�e�;�/��֌�sU��WA;�F1�	����٠���)z�O)���Ԧ� ~ؾg�R��P��;'��i;3]�:��4��(�X5���MY:G�r<�//PWc��cF֢������E��t�x���2�k�bf&6K�q��t��Y��0`�Z ��_�^W8�y���N�.}�*�*�٩)�;Y'R�N6R��=�����1H���]�BH���4��"^�"2F�$Mvӆ0��ң	V�e���9WN��6���zwo����%I��z��k�Fup�E�V��+̸����ˤ�_\6�?����י�D�qy�9�,��@�t���◐R/pE��#K��kt��k7$�߿� ��w�\��] ��ڄ�%��r�R���C��9d��Tv>���i@&��4��O���Kc��$��.D���>3M�2��ƍ�Ԯ���7�9�����HD��ղ�H���o<;�����~�Qʦ�bP�zQ�p������l|e����d����aFt<o�L�����>v�z�jQ�4����LJ֝���U�X���
��؆M�/R���K��x
����@{�Ż鹍,�q8T�6Ŵ��.��W(6�F�#�q=��5���TS��K�a���dn��k�[�<Lvf|Q_W��'C��׶�&�#ԭЯ�\;�_��-g�Q���v���8tI��4ma��m��:�dUE`���ӧ1M|x�ߌ��ENpk�,s+|��H6<5��Kn�(ζ�����%�-��&90�=���,o��H�Xu��*tZ��\K��Vߣ�n�+�i
L��Ë���g=��`T�g��pO�����s�axĊg��}�`�9���έ���DcQyf΄u)�w޼�׭.XqC��p����[@�mp �\Eft�"��.��y�^m�>#�(�����wQ[Ă%�%�������E_Ă�%���Ji�hubJ`�C��B#V��֤���L�tHw'�d�ғr��Y���\0�o�������y$�[f̓��'ap�U� �C%$��X����1A�f�V��u�u
�2����%�8��|M�>L�*^���vO���&ܘps$VX�V��]U��+q�y��j����^Ƹ� �q4+P*�/��J0Jl��ӎ��q��d~:)�v� ���g��\X"�s�}��H�W�SZ�4�tޓC�9����� ��ZU*�@!(f
.�F" ixwז�:��=8
|�"G���+|5c����z�{�.zǛfP��^�<�Ǯ3rj��,xD�c��¬K,鷸b6���ΜD1���sD�b�^�+��\���P
ʹi�K��Z�h��\��E+QC �$��sH�"�{E�TC����x18�Wh�����4	���`;m�G��Ҥ�bw5ąd�����H��]8E�]�?5C�S�$K ��O��A:f- ƶ������ u�,�fM�n"B��@�R=PĂ+�%T��]G٠Z[ ��r�r���*	�9����l�JM��	�&��[c�|.�0�����k�� �Q�-}������VD��H�0
�P��s7��f��#u����7�)�jE�c@k��fn�7(dZǳGM�C_��-��Z�x��i	���(?�c��߰��u�t\�ǌo�i�ʐú�o����/���1��@�9C�\�XA$��'�;��p�n���j��Ym��,.���?
�'�k��/�o�L2�P'ْ��ԕ�#�k�	�נk�K��Fi�x�p+��N����b칱Ub��%��C���MS��	��%�� ]N~�U(��`�YK��0�~0+�wg9ɮѢx��d�h\�4[�+�_�on3D�X�
��7��\P=T��sryrm�N�l���R0Ø^�ک���n����j��+}����0�}�#^�� ���/E?��X�-fT�f�e���!��K�L� �|�K���ki,�樯�����Le!EM�y{�y+	��7·lw�s�/{n��Cu�U����U�ޭ-�E��ݚX�M	n<&��NqN-8�z��w��9\I��jPkQ@��S��h�z]����_�%'y�f=Le�}f^�c[�Zu��%�;b`u���7F ���ɜ�پ
ًi,+�Sȝ�%�<	Ce��.�"2w?�R92��2�*S��2Q�������c�9F|���������>���c�l�䄓���%5��Y�=8����(�Y�Fs���'a� Ik�/m˴yF��=:Wᖒ�Cu�s���.a>���=��M�s"ǘ,�JYɒ�GR�xJ�� ��������SY��&�Y�n��o7֨fY18�PX�Q��b��E��]?8A�W�RR�h��}��l�&@�Ѡy�?=4$�/�;�Z�^�����e�U�R���v�
Q�ǣ�vv�Jg��A��,<=I>�2��1B0��4W����3�%^W�5�H��)���CvI�0fA����F�S���Tk�����b�����_�J\��r�0D�$.dijc4�� �nbSs�����A`i�bY�y�Ar�C��\��:1�U���׉����@o��MP>~gqc�n�1)s����8j
��T6V�ѯ�$�;5$fz�D��u1=�z���� �rk^��Y;����q]��1�;y�=�@��@�9^IT�9l4_RF9�1c�ض�\4���}��"�|��!
m�.IӦXD0M(J�䒩0�a� �޿L_z�k7Kjޗ��s� 9��t]���VV/-�ّw�Ԁ;��,�1	^D�)�D��0v��?�GSQ5S{H�4Omf�J�=�h�FP�̵��x�AQ���_Yj2Z�4��y�0e������T����;W�ӌ�O��1kT��؜�ʝeFP̍]�
�����0�`0D�RF�!
_~G�������������w��̙�.��w/�	sI���P�Ӟ~ة�*��؊�sјH��|��R�˱�7=y�Pvڲ
=��#�����\]R��~v���*���Rj"X���Rg���!a��K� ��c+�oAFQ݄?�[�O𢝩sH����ʵܚB����99�Vj~I�����]w ��xu�c��c[�m車��]~��?z��: A�\�:(��\�!�����zj{���Q.�Ľ�(��M�T�N�!�K�wه��0a,GV��0��fY��땳D� ��{,���t���{�q� ����{�,&ʠqdMu.HD��Xke3����A��ʡ*��gXC��*���8˓��0L�Y?wYny��~�9x&h�5�Ȥ~>������c]��\�!��$�&ɽ�!׷a��c2��C/{ͮ��O3v >��n�<��p�v�G��3����
�	 ���
e�8���L���٭j��9W�����ȿ�����Y�;n'�c�����ݴ[���$C1H�O��ykz�9UGt-P#�1ԋ.O��VR�'�:L��r��"��ӓE�����R��@E�`&H�[T�C=�4L@�^;yR��_Ӹ���s-�f�6���o�����
S0@Q�[3�i�o�#{�'?�* �P;��X�灯��M�kͨ;t�pl��T��*�B�!)~��k��Ų*fTm 9��l���J`�`Jn.
�_���4<�6k�k��3Ξ�s/}�a%����N'�~V��$��(0V�y�z���)��|UH��Tt5�f���(�Z�eE��\�5@*z�]�G�%��es!u�VEy��?�5Q��r��#n�vH&+CZܞ?F��q�Py�b ��?��l�#`��DF�,�_�£��X����t�`Ux�wfB�Ռ�1����X!G��~���=.j�(���<	}B
�R�[�K�_�ݰ��.��0�k�-��n� �+q�ݭr���1/{�i��8��\�9�?b�Z����ot�\���j�9�$��T�}�=F�>o�=��W���Mq���{�6��v���ρ�cg����gf��1`��Ɖ�o�.$M�Ƴue�7L�̂y��\ �;�`���\2O�2��(�ƈ��z����!�� [�UJsŷ�3�I0��~�=�=1����88�������S�g��G��l9��;e��]���m���	R��pv���<���.#�S�0{脵iWө���o/�U@�_׃O#��m�)�UL�pg��%�)�oO����B@k�4�d �#�4и��Y��u���o���.#~Kˊ��ʅs����{�^���D'�_���"�xz�ð�D�P%6_��A�)��6_w`�C{����5¥"�l���87�K��ː9�Ҽ��(���<�B�4��]:^��i��
WHj4� �Y�oC�44�@���:��ڭ�Id�]@s��Y�up������>M�Ö�)9V�bʇs�^P���BB�R��M@�f#���צ��'��� 3��2�F�u0GT��r�n|��z�E7����\��<����ì_C�:��̖��}eM�'��&N0),6x)ĢR�׿�<O�����L��A����?�p��B�1��i�5�����Y��oeO�I�I[f/a<��g����>���[�3�Xm���
_o���*�'z���BZI�ٹ��X�|��)�,�X��U���
f>�T�Won`p��|���d�pRό:�9]��{'1;��Мx/�K2��C�:�-PL�6�d���Q�׸}JD��ū��T�a%{��w��Q�3z�{b9��A~��,00^������r���c�5����jr.�P�,�5p*�Ss�.�r������t������,���W�zVD�i���L~r��8fo�wA��f؉q�79%$ ŴRU��C$3.m�w�@�Zm�o�t1}�x!�s>'�T��"ȅ�U�]��(M�Zԙ�a�$΍W��s@p��U�r�K��h -:.gZ��,�e@���ٸps�^
���CH�����1w+��0~��@���`�T_B�L���S4��.`1��D�� Z(���
(�h�G�&���arY�B�0��RkWȰ�Z��Q���V4	�=`�CI��RU�F���,�H�B�5���Z�9����F�s� d�ixH��+A9�K�3�b�d�`̦5��qᢰq��1;b+�H�ǁ@#EY�bB�Q�.3ͪ$uU�|����]�%�V�V�u|qۂ�3�-�4����1ǔ�n�ن)m�k���hX��"�jv/E`��~B�h�n�jY������m�(
HR���]�b�|m^H_9�P��2�1s�K"��*�g��@�_,��rI�D7kS�������^�U�0�����>�I�м���Th(�e���mR��$��T�5[4l98�/�Aٌ�Z����F)i[�~;�Ij]��RU��b���-�#��:��t[����yAO�(/c�7}�RC�Q�J�V�M�M����`����\>�`�����
3>�N�X����L����g�ZP牘`O�����qx.��S�� �d��c�L��C/���Y��<��>��!a�Nr���1 �^7���`R���C�L�4����R�b�HH�mI�Ґ��9�X$�|�jw��e��E ��1x��΍e���
�PJ��!y��V[����DJ�Ei�L�b�`��k��KC�&����l�w��]�$%�|ikjPS-����oE�r��v���S*�.#�O�\���T`Nd�Kiv��w��N���l^�K�y%���WWS�;���B�	n7���p��Bh�Q�/�7kP�|��g0��w���� ���n�I~����ۚ����1���C�c�v��QV��%���H�cŐF��4jϡxX�R,�f��W�LP����EsK:�;�<()�G;E�ù@���@�mz��-K�f�������4�#lއtd�\����=):�1
I�ʳ��z���D�X��n�[�)��4�N� u�0buY�E�4܉?=/�=d��"��l�����)@���|��;���G�F-���胷���G�2�@S�އ���m�C�%����MY��Y��ς�d�ֽ�7��#9����R�lo��gŊsA@�h�ĕ��6k�*�m��~�'&���4zm���F��9\�N)�%iUy�����S�^�
�1>#X�6/�@��Po��G���)J"j��l��сBY6���E�w�=b�&��4qE�S�4�C�>R���@���0���G��g�4����*��
�qf�O/�,�mI�HǂˉA�(^V&6}��َG��d±WR]u�֖���q�ai�9�� P�Ϩ��-Z���Θ *�9�� ���%��K6D�ҭ�m"A�oȏ<�@��$�qअ�xp�h�	Z��@����j`���u�ۖy�N�ə2�al6(W�)�^�ha�t��|�[�ԺyC��^._��*�5�ɶ�XQ�Z�����i�r�:ok�xg�uE{���M�C�*�j�P�"kd�'��(T-aLR�ӑj�/G�n]�\_}%DI���/�sgZ�Z�b����ݺ:ϊ� 	��J�m��,PA+�g����di��Q3kf�W$�]$3�Tұ��.��ϭ��a�������>b��9�����F���EW���\Z�l�I��ޠ�^M��@X�1}��O�<�m��n���jK{��lxҌosU����ĝC�������KVqv��A���z8���**-�v/��ad85Õs�w��Q��<���������0���0[T���9_:#�6%e���u����6b�������M�����/�(��f"�=���:�vɋx۫�}�chZ�)����MD�5(��v^ZuF�9[��~��/sXo�J��{d��RT3����LUO�:k;l����H���':,=��Cm��������ʈa��@�@_U���+�
.��~c�*0�,W�����	�ë��<Ld%N¸{�0��ޘ��9�-�a>���"���Yӧ�z�C��ݫ��N��H~�~���:m7��͢�f��2�ƁK�P�ˬ�:g�& ��[���w|��?��[	h�k*�ڀgÞU𓓗x�^9���lUg:̰؏3#�E#�����pn��|#ף0
�G�Z�?�N��L�6[`P�1<�D�Cf��8,Z|���:|�ݽ��C��+�?�ӹB�@�<:�����V�c�b��k��Ĵ~�A�������D�������`<ȴq�^1֕|��7���1(�Lqt�^p����J�BZ�N�^�C����si6�mM�3:�HҦ���\z�*����:CR�ą���ߺ�.o��$���]��8�(��v�)Lk&m��8B����Y�n���&�mp9��쟄*�T��%�ݏ�b�2�5d:��!�ʘ.#��A&����U�H�8/5���@I���=�Hr��7eD��c��,a�a�fЈuBx�)ܤX"�4�jO4ĸ ��7�#�B�5,o'YF_��!�9{W���J<aUZ��+�8�*5�-ע1����O�g�9���H�QX
2P��r�L�A���ݟ�����p��������2A��
ѸS?�v��55ؑ|�r,׸�KC{`~)�~$��~��@\����#�A�Ҋ�r6@��_3K���::��������Y3����|�qH���T�d��]��98b�
�\L�X`�&s�\c�11�j�a/K��Q'��P[ �v�)�D�����>�V���W��:A3�,����='�a0�=#b"푡<�Θ���*A����y�񘺟�0�3��B�Ta��B��r��
�e��;����k}�<�#�{e�8�|�Nd����)�An(%h��(y��`�Vo�3%(�����q7�,�g���B깓�o����7p�8Nu��/�a��?���Ԭ���V��VC�ێ�õ��Iɴ���0n4�1��~�����=�~O L6�׻�l�v��T��&�]���v���{Op7O�o�Ʊ
�tE:��� _�%�5��SF��Pb_��� �_!�?Nd�r;���t�ʹȒ�!��%bD2c��̄��$��}�A�ߊk����Ʃ&�ۣ��4Η7pm�|��N�W_z��JhO��b�a�i�)ʠ�/w��W���X*��^$+_��
)@��C�驐l��X��@'#����KO�	��I�:mɝRH�g��.�1�I�]�5�t��7�|FB��y������$�w��gӗ��cGԦv�4��t���C������7��A��1��v�y)?8k��:ܻ�@@T�'!Ǔ�,���{8o���\�>둕�O���+HF�B[��\@���V161S.>4��SZAX�C�b�����Q��@��kgn���gO��\m��}S�Ozzn$�M8\�+6V/#ݾ��V�#MA�(3PcI��1hQ\�P����2����̈́�դ�%���=tl11s'��Uw��X���x%���x|x3�9�%90��G�c��n�j�o�h�r��X+f��:ew_�r�ZI�ݓ�ϖ��A�Z)%)�8m�u*��~H���HvnGi�|H��0۲WY��XKò
����$��Y�,�g�BO�w��������� ��ѹ^�䚿Us��!}�{.ST:�xVْ�N��b��@�'H�S�5T���*�Ag�^�0�,��[�%{�!�����	bꍱ��A�Я����k��@w������Y���U�a���kD4l��;���ы3���=+z_x�#U/
�Lm��>X+�Y��ޛT�
nvTj �}���\ٞR�q���k�88 ���<�9��p\����Њ+H�n(���p�fdTT(�X��4(���B��
%����q{�G����t�ǃ��FdA[���?��,bEG��"��IY���%���h��0�]���Q/�x1p
�b�o7�6��s5�6�O𚺃��w��<vp�ߓ��h��NV�Bk�fm��]��'D�ߕ�"@/�����cALt	WQϳ 	�����b�U>�Q���?��%W�@�F��q��p�?�E��s~9u��;���7��hƭ}�bv����m� �'eZiϣ��mD�1b��O��nw/��9cw�2H�$���o�'�!�|�.�%�4��(&-���7�x�����?�(��{�����6��3'����|�]�Uz�!����2a��Ih��E�����X�9����4�,O��]� ������7�}�Q~ʆ[�� ��s@�@@�u�����l��R�v�tk�t|�X\�hab�
�A�]%*K��w�e��C�k��FV�ރ/u���"��k� �����j��#d����i���}Ee[#��(��"Uх���җʗ+�L'.�'7<��aJ���ʳ ʚVv����f�������N
`�<Pp@����=�҃�3�7#��u��K��Dd�:��.�S'+�'D�L,�5�ȵ��qQ��#u��O�y��$vZ�m3��[W3ɶx���/�f��|T��a��6���k��D nP�����ߦ&���)��t�xl��;D'���y*E�E�_��U�]�����t�M��y��
�[2M�P9H�~�Ƶ��@e��x������d�7u���C��e��Jʯ�mŘ�F#D�A��k�d�[�ф�W�6��$�47��n��&,���7�gz/���!���\8���{�?�t��d?qB˄�"��)b�*���j*�ފ�dV%��@�ʹ��si�;��+�"#�����eW�U��Η��m?7b����}�!��k�a\͌A �~IA�A{��%,J39�����w*�kW���r�Ϳ�At{Ɓ�O�e`����� .���p�R�m�,�<�`9�\*��(/�TG�V;�/x��V�LjB � �����*$�����jq����13�ڴR�7��U0o�=7�{a\���$7ԗ
����J�����  'z�������T	�]TG|�"sS�)�����8s��f��+�zkU��8��qG�pc�
����&~\�R`��1~Dz�x6��A,�쐃��y��Yo���SаSl���VE��qj��=�*_f���F���\�X��!�B�W�V�A.zɰ�G@��Ӗԗ9�񺢢Y;di��:�q�(�b�jM��>q\�G�7㖏l����;S�٦���2s$� ��U�T�_�¸���LG�/v�m=�B=	�����C�u��&U>��<.�ۜ��I���lQ\.$zT.g:�\衢��Q�	#P�n�Кƕs�l&�����b;
�΢Y0H�r�ʴ7XY'\H�H󛿋N� |f�����v"�:v��ÀK�_�#� �.�Z7މ����P`���kK��g1�����`���@�GV��J�%��P�Sh�%knEd��������]�зp��:�!�I�oP�mb�����V;���~�aj�zi(�t\'�W���h���.���k��vJ��ͨ����4y�4�����`�ߤ��3��rf=h� E��A�5��/��06;0�_���d	���6�n�?$�����
�-�����\����ʕk�u]���4:�Q�g�f�Dǅ[)�	!�O�����ykf��?70�"�A9Tuz�X�z��&�@\�,�R�ҁښj��B
�:�[�@2�J3 /��D�|�k-u���e��8�f>�K�)��eM�߭���B9 �x# Z��7�fB�k^�"�UX��x�*�b�s[L�O�~H��;��H� ����@��G�(��ի	�5,`13�����|�'�	M��$'�q�n�1����L��8�s3�a��_��-�
�9�J=b��c�jZ��aK��*Ӄ5�`RP�����{�K]#*#��P$�VN����y[���f�K%dSI�M��i�u�DN ���;�!�0��q���*Љ�~���{�h"%��J������<�B\�x�ި�Y��2�����:O��0�;�!�{��$j��eU�b�"����
20ҼI��ӏ^��n׀�e����l�l ��/�J��7�ɗ���Ϡ jM�
^h��;29U��l�>tt�ͻ��aͮ�"
d��+�=��~X�|�b4p���$�
���sf�5�Mb5�$y�t�����9z����J�c��P\�z�fa��C,��o.�s��9�� �M|�%�D��;���iN��:�I���6BZc��V����z�z�� ]��~��#6���2��U�yG>Y8>"�ȣ���
�f%�4��1k���*� �[L<�Ap�l���p̬��f�П=��	%2j�e��_և��!O�,��4���!�ֲ�~���䊣�VN@QN�A�P�jٟ(#���Q&�~�t�ջ�T�@�4�m*~�k�����ĤE溘D���|�;b9]��մ4C�‵q9qY��p���!O���$�J2��@%�he�� {�/�)*�v
�9��j�SV�V0;xG-R�Q%�s�;0����QW������J��6�0,:��
�d��t:�q��'���(�� R�_W�Q�bW�'C�b�"�������N��b`$�}_&9f�|�+X���c0ET�1�sl�N9�g?�(���I��):)��bx>)����# ��J�T�)���$���^�9��;SV6�gq������n|ׁ#o�mS^sj>Qn��W��u�x@�y�^�a%U�����m� :�7@������3������]��	�xbV��a+�x�|^T������4pE��)�hB�{��rV�� "����|D��-��[���҇A��'��ĶK�����)�U+49�]���j>�5pg�׳���GT� �$&e�Yq5�ۛ��)]���U�C	�J9`*�@R�Xg�<J�^Y����2ׅh[*D��<=���EzJ/O-���Or/���$�jD�>c(>[\�����ʂa�pm�����^�"t�q����Ԗ�:���:6k꘱�3�#�J�>�<�CR��^�w�z�+ξ
֢ƨ�&x
D������3Vb�[��@���!����'��M\�d��<*�Yz�6!����YsZ#��Q_˷pi�}y���,�r��@F�$���<R���� ��=g��>S���:x?��_-�R|�Yps�X]������E�?���M��sj{�w��69fq�t%�+}?��R(`,ĻO��4���_��y�g�v�wHy���*���\�τ{=jܯ�V7*5P����!��}���7��6	!�t
�q���AX
Y|9�~Vy�,zm��v���$�񩛙�g�X���1=��\⽎��8ܿ:C�(N�R@��͌!Y2�ꞥ��`_D�{�/��~������"m�O�>��8A`�g�խ���/W&�]U��B3������Y��.
�h�F_5��S���/�ؔvRy�.g8�;mʙ�I���t#qZ�"�I��2��N%��so�/Y�O��Wv>&�a�!u�q������HF��r��Z��,9�a��r���Hl���~�LA�*����I��
�;���~5)d�୒�gs_t���onK־���{!�Z�f8��D�?A߫L>���r���f���[��:-��8IrU��^�����~%ct>�@fyT���v�����w�J�{��"n-��I����Yz�%� -�y�X��xqp�$i�R��a\��J�����(0�N���G�S�K��'�X����:�Cˠ�r�qsL6�E�gpl��|p0Z����V^��כt���!w���#�E$bV�Bv��aԸu���&����Q+�&�ߒ'qn/
�����,��`�ʔ�l~���+��Ę�+c�1��-���y��c�Ю��Q�e��:�/�z��L��>N����z�qyZN���8؏Ks�Wl5���pPc�m"ZΤ��m��u�CE�q>��-�J�9��&�6�O��!�Mg�X���t#���z2��*P���:O��ťrJqNk���}������b���f�`�e�z�GU.鐥w{m�m��4���*Z�\h���g"��T���(b�iZ.3��׮�y���kB]{�6ph�RA�oO����Ƽ&F�=���Nx�	3��`��)�T%)h��5�ޓ���s�Z��k�7{
��*��V#A��Ԭ�=t[C8�^���g/������X��\���85C��I�����	o��kjhJ2ye8G��z7���B��ns������A��g�+&�jg<o'U2����e����圷 a� �)��Բ�ݍ(���1�EB���ɨ��� l���6>�}��7tcN�p)�n�Dt�5M�N� �Y���aёKf��l�%��7�����w�k���B�c�]-0����˘\NR�#�����n��]O�{w��;Bt��h�z�;}�+�M�@]!-�_|��~�
�՝՚L��Rw��t	�Cyi�x-����"'ϰϋ�&۰��q�XLi��/����h2r�t�[�yHE!��f��[a��N,���tؒ�ų�ۿV�KGy���T#�ǵ?_����G��~e�0�8?�����(���f(>_x�z�vZ݊�2l��i�Tٚ���Q���ݛ�IHI{f���oG�Z��o�S�����eU���T�El�=�'��1���)�P�ڐ��|(��c����nՂ���R�_/�U�`L ��"�Kb���,��Y|�o���(�X���X�C �5=�r&�#q���/}V������nx�  �77�$��R����Y:#�9�x���l�U�᠌�Eݵ�TV�kk+Qb�@��!]h�0��	��X�w�~6��|R���M��8�λ�z��H
���𞙻x�p9*�������A�[5�f���`7|����6�e0�#���L��{����#l.D�*GPaHj�ۻ�i��2��3����"�/�.h�3sd��Ǽ�,QϨQ*�ß�
^��5�	lp���%�cj� fj�'ڥ��LX�(�+#Q�p��s��r�q�s���a���!��+,A��޽>l$k�p������9ʝ]X�fa���ƥ�ݼI�f�$b�@R��w�D�~��i�df�Ǩg��v�sL����C`��������_����380�`�����J��^7�����=G"8�t�;k� ]�l4�)��B�S�y��C^�hP�{�d�p{Gu0Ѕb�FY:(z����)���}]}&�~��@�;g�1���14���m�m=����aV��rbM���?V�M��$\�W
����#=�Ψe�Y~�2��=4��G�>C4�ϧ�Q�l�����3l�dN V���;暀~K���?��zCV�+���{=#�(^��B�FH���Amn�i%�*]Hf�2��馾^i˒�Jp$��7(H�맯�E�����e �����Nˤ��ݢ��f[�&Q����é�"�<o`vb��X��K��l{H�O�_C�x�>�Eg�}�ćP�d����d~�$*!(�ݴ�֚&���x������
�l}�{¢��AƑ���o����֡6Q�a�(�Ჷ¯wOޡ8��-2�;�h���!ϕ�t�P�£�<����Z([����n/{�I]"��'��m��|��U�A����g�f��=Ax�J�&6���x~@x���D���f�������wv�)C������#%����.��5��PN-��6�`U� "�(R���D��F0M�=l����FY�.��,�ɗ��8C%ԄO=[��B&���lzrضtO��Jک��Xo��SGC�bf�o� ������dEǁvr����$����5{����T����.ގ����r��ݺ
M�p�Ht�LP.��Ӥ ZZw��g� ����]�R��8zq��Q�O	�uo��8���b����+������BE��*k������+�����H�l�l����+D/��-l�����?y�?Q���1U'�eF%hA�m)��m���������(�E.�K������@�O �	�p��3f/��΁���cK���me`�s�N}��59�+�S����@��h"򆭉wWf���	��'CųXݚ�����3���P,���	(�&:"I�d���`UD�C�_Y�,e��j�5,�'ٹ�h�����'I.�|�>�C�#jh�=p����1K�u"�P�"�%T�=�1�������K���M�=@�ѵj��Xb <��
�/$��Q� :��a[�`����n	�2Vl/��8j��ѽ�9���8|T�,)�^�BVw��s]��0���l�tbv�#
��{ʊ+ӏZ:(?��ʳ�Uȋ8�u�[:n�@���½�f��h�}���5�nMxVdft6�p�K�x��Ⱥg� �8��/�HrԌ���������Ē���h��A٥�Xz�]��.���o�k����h�y�A,�ڋ����K���%��cSΰLY��<|��}�*��n��/�^�N���'^��;|��[�J���f�"��y��ZJ��,y���I`���ܪ1\�?�D��u���!���+&Hgu�ߑ �J�P��t���N�IS�[�i����*�g���c��,~��;�NP�����d%XSU�o��ʐ@Ϛ�Z����	K������-���\h΂��1'[fOX��J�J�����n_�V?#\`�vy���Cмu�}��c����p��އ�J!��uyv	��E��vpFM��Iu@��9��l�P�L��'���Vp2��b'o���#�L\��N�H+눒$�z$�=nHKǺ	���^�c�"n%s��4���N���_�K�bZr����-ny����1`ɡ�q�(af��啃L,%�OQ�rA�x AA1D8ǿ��"-R�� DM�Ю�������D�~�p�f�$�x�a�$�AEP �I��&]�@��
��1bl$��������LQ�2���+�|N?a�B���F�wO�[��7�� ݇}����ȶ���ܽ��N`��k\���Y�B��ٰ���������Ps�̩�)�t�:���d?��E0�W�R/��ő֏�[�W2�D��}�UWL��@���~�Ny��}�`�b���R�Xo)	��Q &gZ�w�Vz<B��^�3��O=i������ōD;������ ��	��q0��v*��B�D��Ub�3V2v����홑���M�b0���k��kL�r�W���Y���c�"P�ÃqO���H]�߀�>P;W"W��Ʃ�OJ�XE�H�����M�~�5�<-�co��u�t��V��z$�����Tw��~뢫� -�5����x�.W
P_/v+��y�ŐmB(�m� �A�N/��t��h]��kv%p���Yq�멂��ɋ����Y�!9��,���c��$��և}C�xGv-N�]�q���5��!O�MY�h�ʹ6_��)c�~�h��Hp^��Og���ɜ����wN^ێc�$mY��'�2�Ȝ�A�>� QB��B�@"��"ߣ?�r٩+�����(,9"BoL��L���e*���WP|K�l#�5U��fǋ�!�����I����9qgZi�j�4��� pКƽSM�%j�)M�K��s5�d������^qc�����̬���D�7}�^��,B��&N� �LiE\;���8S=)�"9��~��W�	!H��s�����'��"�O'�5�<{�nϋ��Y��w��d4MEĶ�Մ�|�I�s݆�Dέ5p��d�F8`\Z�T������Xڋ!A����~ط��`���.�|��}+��N\ȯ&J��0
(�0ҥ-�n%���7�Tˆ�j�w�3�\J�ڸ;[E�e�:߸�P�ԁy�9;�����x��T1\I�"�h_���B8�r�|�>�-��ZaFJ�x"�2О�c`�Z��c�P�(����м���#��$��Ψ��~��j�K�רDa���9�^;���Me5I��R7�}:�h�C�n�<���"�IRsdH;'�"%����x���9��ڥ��%���e�g�6|k���� ��j��|/w�X�+�2JO4�5����ߩ���Y����Nw��Ʌ�����aQE�A��wԙ� ��9p>��8%���u�w��z���.�DC���"|4N4'?`��aIV�Q23T�p׼���®k51?��1��J��j/O5�=r$�y,�9�rb؜)LC��Y��qo�V�Vz�?FN��Ό� ͪ�Kݽ�]sMl������á���)�x#�����-�Wl����RR$�&A2�
�p<��npeР��o����;��w�V�����l�:\9���-.��&���t�}�6��AA�������ǵ~4����,nZ�p��?ز���r�ӑs��P��,�IՎ�B������T���@��Ye���"��Ee��p���at{��ez7<	�}L�d���w��ր�f��"���S
(�i��f(��J��-�
��,�C�b%��ĝ��"�%�l��c� ��ɸ�ŷ�ףoA�5�>�+��gW�p�P�)a:��*_f���3��&ǟm��������o���:J?��1�r����)QVO��O��1m��qlA�������B[��.�Q�46�Z:��O��3����.3J�$<�b�~��U�/�#�� h�l{	ػp��&�9ic�tm��{��U��
�����<u*�Gq0!K�_�j� �A�p�&$]#@�M�x�,�3�uq<ry�i� eݸ$��[��1;b0��Sڢ���\�-�����Mt�qCz)�F
�Į[h��5�zH����ʤq�ǅ?��߫�i���B>᫧�H��R8�ae /*3�̺�����3��c?W�n0��[�|#�6<���}�z�N2��
� ��r��.` Ju}8��-��|yB�9��,�.��Y�"�������O�3t�ߓ�3vg$O�v�7�ǵwB�)�v��#b��Ha�ݦH<3�T��b���\s>�E�0��`�[AS��ۃ�(�ßm4�j�^-J?��C�{���â�B}����R�����۵����3Z�0{�&G�����D���iS�,:��
Ę�:�d��aL�ر�v&"�oc-j��Ukg/���/)���*U<�j�Ag�0!%$届��K���K��̗@��ڝ)�����l'�:�.�˰�g"����b̏�4����#H���v�v,WU��=�o8D��ȳ��c���,nҫ��2~@s��*��q�Xk�sQoݥ�.Y��=�j:�e$�O��1V�΅�[�ݣ������h�Cl��g�&�X�WU-�:2V�g��t?�fH�uЯ���흥����ڠ���}�n�%���0.��Eyr��Ւ��j7��]V���{9%�vdR���w	,VK'��5���gA�w������f���]���f��M	ab���K��u6t���m#E��c4?�]�_v�}�*lrك�%agA�r����,��@����yh0%��3�7,��cLV�f�k0�eh�﫤ㅱ:����T9%�v�؀���Ӌ2e�+�ځ>�����������S���b�x!;p��W�眧sx�q��F����O���M���F��/�ǰ��7/�0���\��KM�/���I��?��}v=���>��/��O?�u~+�dR]P!+�"|�w}��1"�\�1H��ASoQs��[���y.�J���^��E�V���1w��>C��Iwt�E��;z�Fv�j��<�B]�����Ӳ�,g�zJ"֫#�6uy�{	�da�QH* ���.Tz6�C��.q-+y�j���8�������}��~��Bͳ/k���5�}�b^��RS���GE�O6
˸�� ��x��#*�=/�w8[�.A�d1��vs�������c�Qš�L+�`+Rw��91"�?�HdC�汌j.�q��L�z�!{M���z�k�}4lp82km{B⬂:*5�e���0}����d�
���߀q��"9P`;ޝX���fQ,3��H�8�n����"����Ѿ���`��#Z��湭e�V�-n88ٶ��:���F; ĺ<�T�9�pŢ1�v������L31��t��v/ǉ�CvN
f_�Q4Bg����xN��^4�<��~��Yi��ߣ����p��d�q˽Jפ��tb���t�7���_�5A�=d7�(]��P�i�oce�R�1���;n��SQ>6����m���Z|&���}���&b�O4�3w���ٚ�����ͦ����l��<���ZE��XU#��ɛ�'�@o ��z���������>�� T��-�e%��8wc�����%�rG@��~���l�;'���Q^¼<�lH�+G�@�T�JC�=�5w�z.�*��'�}G�|[�۸�6qP3i��v{\����I�琄�$N��\ZL��Jv�K���|�:3�>0UN$7�-��_+�>	���U|����\�^!Sȯ=>��>f������}X���R�[\�X�	���[pO�b RF���,c(>�9�#�͸�j����&d���T��*&���� �g<�X��~����n�i�g���K�m�o������)(�>22�#�?<�8p�x�
����&.����K-:�O���|�{���$��>�G��'ie�|"XO�u�9��33�C�U��#����c�����,sz�}V֙=��Ed*��X��E������2!��!1Qz :L��&��Go�oR�˥
!�8#{�r�^�B)^����n=s���#��@��pT������]��Z�a��=���ޔ����Df��yq�>���	��&zҘ�c�	����U0�ܰ�ExP�ZX�a%�6�����q}�y���<��7>�|�W'A���UGc$S��`i�R��겪�5�MGrߍ	Ϻ/�����[5���q�F�D���=0tf����^��m���J�i�Tɱ�ŀ���͡�Qj9��%���(Ar\M)[�8���=Rt4ͨ�|k��i�a�@ǉ�։�^�Lt��K���*�5�Qs:�w�r��.��)W�����t�����(�(!���,ڑ��$}��o�����'�;j���/趃����M��y[��:n�w�9/���!/ ��.i>6���v�Wq�:�l,*��o֡�%���bj��#;�!3:�����\ 6Q0��l��O�8�Ԕ��ڥ#��$�
[j;]̅���w�75}������m�2�9.;uj�x>��2�t��;�,�2p[�(��C>go�©�i��,�7��.���}R���Ǌ���B䒯fc��DB�c��y��z��jYgw��#���|Ζ�R�v��E��=ih�lB�#�
��mR���2����� ȆT�A�=B�Z?���$Ī`Yo� �O���
@�z.-�ay�T@�*���P�&lm]�F�0��afz-��D��<k��R��3wuS���9�E���5������qL�'|+����{�N��lg�_�J���pu�h�4։ʽFT���̷�W��(-��b��j�7=J��:y��z�gN
��v��8��P�
j-��ٓ2~U�~)"�gX\bL�ǘ��B��pIxŕ
���B�A;��ԂQ�ǓI�ǂ�3O�u�/$����1m��=�t�]<0�oʮ���FYu��I� pAx��6�q~�49������2�Ku:FB�o���_�V��gOeU��O�P`Sn;��c����O�!��~���FMP��2p5n.-����ӊ�����w�uoV�Hr��	�� �R����n������d���IK�ݢ��2dܒ��O�،����U3��odNb^�pn|v��B:NS`.%�^ ��z8�p�<�7��H���7�� �>��`�8�m>���-N3ob�J�H�P�Prao�2��"o���a�8?}���B�
�l)k������5!N�$�k�.jz�u'`���u���OG��T	Wu������<WK���5AL�L�ق2�@5�_Y'w`b��n���3x6���
�������#+�o�L!�� M��9�>1�K"M�����P��fK�E}�\�ɧ�&+v��i1_I�aՆ��FZe~�.:3|u@˵ݍ,�ΪN�����	g>�^	�~��q�i��Zn3E�=���ޞ��(��n���I���R
p���0D/s���:6x;'-�v�Ή3�����eq��~�l<3�u�tʀU���h��H�9���
w/���9��4�K���Sɣ�8}}U�a](~fy�ؔ���&(�9aD�sa���3c���U8Av⚸,���< �aɅ�����!Hq]bkv�W ����*c�t��_�<r%/Hރ��l\�l$Ϋ+���Vp�6k���w>H>/IB\�oޔ�r���;�X�I+��Z���c�ZOamr�d�-O����mRg"�{qr2�m�rd�*�'������+%��zi2�p��_i�_7b&Jxm��$����8ˆ��7D-���3��U�_${|����K��!��sޕ�
Т�+�GCp}�v&8D���/
��:��"Z�@�G��ى$C,�'L�"\��>?�8�jL%u��hT)8,!�4�� <I'<˭��"��@��?8�C.�秩��@R��Y��!A^t����EƚH;JV���f?��3�T_L�}�C(��@���Úm��X8R�Pms[y�I����I��C=�k/�NA��Dј�F���fBÑ3���P�Є=Nl�}oFfdzT�,0G���Q�d�Ҋ�鞶��p���}�8SmE����y��Ȝ8�6v�������:��>�/�ߔXD���/T~�8:�6���]i��?����+��nz��D>��M�Q���H<ښ�h�?����x��[����TP��\��1���v�"�؜�\7QM���a 
�_}ət�	:�lV�;'���!������i�/�܆k�aA%nw=��������?Q4��F�J�N����#,J^z���y3�٪h!�!�U����'Kő3yG?B�C�!RR%J� � ����� ���q�`I߽�(�V�נ���b���~3^P�l\�0��&	<���=�����`�����:V2�6W2���<ð�fX�w�܆p�;��.�4o�{�,Dɹi-k&h��d�c��ԚQ���Vֳ�I�爗�`�]�9�|��9��<�]��[O��QĠ����P`�p'�ԗ�s��=ӥF��/`f��9�=��E���caRe�0	1� s˧����A��� _0�j���_IK*3��9��GC��S�U�0/Z)���!=f�ɿ糈��i	Ve��bUi0Z�i�`�D�ڀw$ ���|�Y����S�\��8���2��$Q4�(h�H&�M�wP�X�]E���O��kU]&[oR��2��>PE����;rL���ظ��a�4E7�b����Qv�x�i�kOi�b��T����|2(%/=N¸�����\9��񑛗��`�^Uq����e���.T�n!5�)�q��D(�����i}��e���.�5��r���D���P>��Q��O%<<+�I6���}3��k�x�V��m�&IJC�~<G�'����
����)跎{%�E�uHM0����l���&S�z�娚�Xq�P���+��0����ʹ����&���s����Lc���m��R��X������HyV��,I[?H�+��qNh���j�� &��ް�{_+GNx݆�3s�NV�z��7�SJ�A�?��Izw�(�]��I=�D���TTL}��f�v��,\�;��n˒�z�N�C|��s�W���mw���Fc��b^z���^N�\d�����@v�=��c�MU�̚�YxZ�}A{�]#��ZUA�dpi��+��ID�dW S}�dh����ԛx�[+��U�������=s՛��ݒW�na�q�?/%��@wR�]. Q��n�Ȣ�6��gV�pKI!DIN����5�`�C��9���HX�Vr9b�Uܶ-�`q����OzS��
	��m����T"�m�J3;	�oT/���܌�=|��A����7e�c'�V�U!�DXY�7+M\�z��h͋�Q�
̀��h����Ϩ�O�?�	m�6��ME\WOw�g���z)g��<tUd�v��3��Ŝ���B�B�+��'8y��v���v�8�X1H�5#�)߽�_��X���������B�Ube������Y���=�t_ٞ�s�1$1U�幦�j�#��fx�*�e�ApL�O����Ϗ���4�Q�]�v~��	��_WW�Ȍ+�?Q�b��zRJ8����^���>��{�6D��|M�gՌ�v�x���#R�U*�J�=�$e��)U�eu,��7�(Yƨt,n.�-���3s����ľ/찆��ͻ�*�,>x��K�m�^|f�_�X��]�|�x��h%wn�R[�����"��BEk�kի�	Ī=���]�k�VH��<�\g��V��\"���೘t�����wZ��^g�6rD���A�Uk����������$?�p�d��$h0��Lu�U@_Hl\eq7���v�YSi�$K��0����,G5��տ�Sf��.d��?�Q��Jg�������ȱ�\��S��6��2�a1�	vs<�h㟯d���V:��0>M���J��EK��k�����4�c�8-�d���h�����	˩���dD�o��㽧g����cY�Ո��B�/��-ݙ��̴��Ha�i��K�,��!�N5C�������*�+U�Y���S�^�t����H�2oML/��u�\K)zB2!g�U��I$P5z�׳�e"Q[�V?�a��:�a�Q�;\Ei��3o,��\�o��q�sS�=q�t�Q��t
����
��Ơ�]��2���0����r�ً�Ģ͘��So�� p�˰i�,�T}$b�p\Ϭ�N��H$	rs�A�J�H��Z���8�l��������M*)�m�<�Y����h Sjimv��S��1W��po>�?߿ �C��JG;���H.G!�6<J�.2.�.hSkw'�#^t��v����􃈑 5}�Wx�M�Ɔs������D�J�O}��L�d�ŝ��I�+y��h][IP4!J��]�+����Ng�K�4x�X����Gd�PeP��9h��J*.��hh���P���<ǟW�m^�!�V ��w�h����-"5�"���X��� �4�r�3=�e^�`*nu�`�a��'��-iVKj�ar#�@��3,�n7e3�͒��p��0I㻠2���F��?0�(����hn���t!���s�lV},-=�	eȒ�Rhn/ژq3C�Xу�B��u�$��?���1T�r�3���g���GV�.�T<* !�E��I?�ѵ�k7p?<dJ:F���@��K�	c 7�♏��)*8���z7��3
�x�}�s7�b	��*�{��7L1���1�E"gɨ&X&ޝ�Zu��ʱx�|��o:ߕřO��V&A96�xM邭�D}|�Ї�y,�8<Td2�?*���%*&�Gx )<���H�\S�,�r��˩�E��lԣ0�T>���kFAAo>m��3�ˈ�m������I���s��&ʵ�],�'a�W��fQ����H�G�獽�m��6��C��ѝ?f�&Si<���1�0:��0��{
�Z�q��fI��ak.��
6��f���֋"����p�[>Ӵ�j�!f5T��ոӼ�As��NG�W?�	O��ƳlW\�����ga�����fz3�rbGB�o��F�f����I̢ZM+u��4�=]�a���ˡ���i�"��d�}F�T�4>��4�S�Fo��:e8��	tM�	-פ?�$���+�����78Z��Xyv6��p���wX%��v��Ű�EZ�wr"��s�P��;��1�UN<Q�k����r�4?�f̾*����tJ��P9���$l��c��rKll����5��zqZ��y!��0����V,S*��=�'������^O`�1�)/�&�wă���7��P�F��j�f��,�_��9� �P3�ޥ�+W�U��L����?��V	��������JH�ސ0�L�O�(d4
l-��˗n��	Z�
-����;�4o@���p��-��v�T�9{ ��X햖�&�$���i�@,���#L��MEX�RN	nQ�u�/c�v+3{Xa�a �O��[3�	[�w��N�	Fr���ocd��_�kV'����H5��H�D��}���hp^���m��nP@�h�;? ��|�aMfc�u�U���H�ۮo[�c�;�+RN�e��
�z�h��lW��ڼz���_����|_єƋ��zI:������Od�БZ�z[\�೿��beB\���k�BIuV�"آ�ψ���Z]4�{�i�3:Ψ8��{�E�5y�噫�e�̆���dʊD�)�S���*�oL��u�5�!��p���q�p��5�bi�7Jj�{o�XlľB<cH�Wr/����h5����x��R �����*�N
̉�}�(��}���RӉ6�(2kWC���N��>0��^$�	EJ_o�Z9@���D�X,����C�h�����ت����Nj��� 3�<5f Mw_��<!Ϊ����w�Z�CZ5�� �a����3+�?�2��T�%�a���Q�Wh�ͼ�ߌR��>���gqفk#{F��I�.P�ڄ�S��z��_9(��4�)\�GB�biR�������0�*�`Cmv֙�`�k��C�ň�UM��� ڌ?�Xd ��L�L�F=2L�C<����myw�L�r���~�\.��]�Qs���kMVM��*y��B�,zΦ�b�T�%i�+9?��<��B�#���ݾ��~@����t�l����+���P��`�ďG���pt��X�)=�#tE���x*ۚ�鲚�C��@s�Ѱ����*�G}�,;��rڃ����C۟WiS���L��P��J���^��K(�H��(���Ur���$FCM��[��Ѳu��\dE�Ci�5�^j|~6J�wҷ	��/%Z��e�*p��؃���9��~�V����]I!� ��;��6���c��g����:�S���n�U�)u�E�A�������]��{�A����2T��?�UO_���0��I�����R�H��-9�hrV����<D:����{cٖ/~�Xd�Y�hjL�b��l��q�i.�0r�z^��Ap�p�g��#����hdG��o$_����2T�T ^��K��!7�ɭ\B���g-���bh���o@uG�L��cW}m���<]�g�Qv�3#�>d���jAƶ`���"B+aL�i�EJ.�����F�z��?�����
T�X�LQ��*���-�#��"��ƚ�ф�h1Z!�6#�J-!�R˔�0�w��r�EG�'h�m�����x���W�5	�t����P�f5ƨ�f�����T��IFP�j�]������9�,H�<#�1�p��x��-2��8V��E~�A��Z6�>���"�1��h���Dyi��ES�Z��[u����6˩*�Fe�
�\u.Ń~�T�ӭ@da<e1�����i���� MK�P�j����Zy@���
�S^�w uԄ͒��}L����tP�"s��B�KC$���8G�Lp�6���=�=��A��a�e�K��:P �M����Q�E@2�6Jr�(��'Õ>CJ�� {����Y��ӕJ6������! j�t[�ۃ�X�p��)�wf��dZTcL]��V߯0�9�6�;�%T�����"M���U�*髙n�Y�E���[:h!�M�l_��#��Q�8�	�s9��+�c�F��߼ ����S4P-,)h���F�#ÿU���p�C��&?��lq�YM��ߍ�6�G Qr��pZC��v��C�͛S��ů*4��-�sǼ�?�+���y����T�,�З�0y6'p�_�͝u�
W~�y�M��X �&L;8/|Ftt�a�_��E���$[�|�0E�֙~r^��ƻ"#!�|N;e?RL�<B��p�rIM��4��XY���NΪ���B�<�*^[<GY��,'����qu������M	]�ü�G� �s��ht\|k4��x;%K���eV�Ja��!�QB �#j�@�w<m/��/̰0QB�q�q�GK��|��/�����l�� ݽq�R0��/������B�ꩣ4zvY�ag���	�o�\G��;�j��0ߧMj��8`����A��؏֡�@��̜��=�������_�X�l,�^s���<�
��E;(�T��c�{-u#��EUa�.���}֌ڇ�����-���MB/+�
RʠW��4zb���"VV����i}��2[�.�hpyT'4Д�����HŢ�,Q�QǤ|q{��]U�7�Il���x�,�@`�;E�$��+�'
�($�C�� �8lW|�*h?�.�ӳ~N-,}���YL�>+翀h/����K?;"�t�eϜ��t(��=!?���a�X���`�;:`�^�^r;g�i��?5�B����a���u��w~,5t��X�rU�I/�+�Mx
&��m�|H/�'W/�b��v����)�ׯq#߁��1����<��?i5:Nq�RR7�#��j#�G�+�q�tu��	�J�6�~Tz���.ɦ�2��i�>�
��,��G�=!q����8]S'��54�e#����-&�|�܇�������B[��^_������9�V��2��z��,sH4y��I�itkN�/�&Q��ף�����3��<����x���PȽ�5� #%+�N����?9����ɞ�h��}��L'),L� ��^6?O��ޣ8;1�2/՗�I���K���%Aثq��^��#~{f�`m��V
w��{I7�'�RoE���<L�4��N]c�%�i�̟�}�	m-lX��'�ʓ:<:G�R#������Kx{��_�j$p���V���9C���ҰN��G ���JY�%k�i:@"��l���b���l�?���a�gkv�G��zc�ОZPN��,a,yZrD�8 ���8nD;Q[,��W	��r689��iR��A�����0��_N�u���?�â'J`m�N�Iy�
S�)v�Wd��"��6����k˕�_,mO�*uTnN#N���]��~�a��:��O��F�df8M��G�K>ZF�I�
��H�; n
e'�N�Fpmf�b��7��oI��
�F⟃v�@�#���ڭH&����0��SK����$z!��W�6WU��P�����]3W&���EE��E	�Hhs�����X!��y��?T�i|k�:OE�.'�PDbgt;] rg��׽��}"ǌ2�������g���Zg�~���,$u���sȉ��[�l�ALەmWxE� H�I���&]�󍂘r����_�OP ���P�1� �joi܋�b:���⡫ E���	[H���Z���UyE�z?�f�4Y���ܠ���Р���@:B�a�%ߧV1��c�z�Z����(:m�u.����'Z���y��H����E�I����\"��Ѝ��X֐���U��<Tv(�3nJ�+I{�M�'s�N�v�_z��7+���������_��������ʾ/�1)�������]3tL�}�������6�!U:�{aMj� bn���C/L�"u�y�N-`n����4~6&at"x���v�rb�F��E�TK�I��_�1%F�oH_Փ�#R�PV��.�W_����D`�e�~K��]+�w��]u�}���s9��������COUE#�x��p!�Q���
@������D}JDф=�ݜyE=z��^�G��m`�<'����˰!�sh�(�Ϯ�c����M�X"鳀��l�l\dB��_g��+��}��΃.!޴���V�<d��b�K��fS`ѽ��0<�pICI�����w�)Feh����q�QS�t(��a��͆�?�UH��~�Zt��>���۸f���& !)#��?�l�a�GD<j%�NcA�V�?^W�I>�d���	����g��E��;4�hN.��Xˣ�T+��p��A�����O�YJ�~8̴�������G8����7�e����f���K���$�ŀ�5�7R9�DH}r���=�b'��&�& �5:�[�i��oS�K�D���z�m���rn�"Hg��"��_���`Hqл���N�� T�X�s�qp�Jjҧ(����v�~m�C�����H�9�?%wu��(��.���/�9
,`�@�Ωg���z��ZI�S����&3cCT+��v��%Q���b��G�?���Oo�N����َ�1��J)�i}����Էv'�~�Ӗ�Q�qOz'FZeV:���5��:�O_��0��Tz�0e	֗9m_��VS��-Ձ w�
��%s�;aŕ.�B_�!� ��[�x��F����8���z ���i���
/�Q���"�C�1�V&Uީ���.�QdH��2╿��iV�bK1¨nߎ^8s
9��0��ݖ���vY��?̳�5ǘ�=��-�+����M����i���);��f<��9'�A��د���+Y�3�����8��
��`��D����R�e� g,ps����6��9��50��b��dR�����_|?�i�.��#��ά�Ų��@��AxH=ᶫ�T �M��\z���V}a'�]���C_����wؤX;ͳ&t`�ڣ�հ�nxk\�p�W�Ճia�S�L!wh`���B� ��W� -��"�Q�ug �*�_��Vi��Jl-�1�a".��eo���_F�Ʃy�)WdB�!��!B�B���Q�H�rJ	G�DŸ>�e�p,��U�S����>��?�0��d��"yj�|y��uG,*�nuR�%\O�ը�ϐ>"�=���_S"������^7��S��{�M��s���.�\8Ϝ"DU>q ]R�F��#�����U;-����B?D�z���qitN�>2� e1������u���5	q���a^l@:�i��r�-5T�b�Fq�F����d�@K�}��)Csn<vݎ�I�Z��3���[�H~�"c?!C���t!܀�M	Z�$���P~|*����F�M2��[}_�e�(����nT0e�Ԍ���ԃ��p���hc4Q�>B��E:�K�PCP`�4T�����$Y�K��n��E�s��6��