��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��TdO��b���F�Ǐ��j�&eR�Bb�ω~]�,��ī ���}�T\�Z��֧��k��v����b����NWP4+z{�G{b��� 
��`⻯��c���s8�)�S����x��|��R}�y�(��H0l��5ؗ{��VŔ1-D���s$�zܒ���� |�3��@�&���9ͳ_� n/��<i�Ϩڴ�PE2���^̓ϑ�I��T6$������Z��wlrTu6T�O�/.���`��6�=�H܅��0&tne��:(�ʳw���K������L1���s�n���A��+��>�fh�����q��}��R�X-��ff�c��K��,ˈ�bU�v�>�@i��F��qf�J�����G�6<�tu�PL��+'*�s���Ps1�@�)��M!k?/<>�RDP��_Y��b#ӋU<0o �.�"b�*T�mԦ��42����(=�pX�c���/�xZ���U.-�̓��\9��K���x�(;>��=��x�|.#��'�u�
��/�������m�Q�|�X���_���s02W�!�IƉ���]C�t\/�2&�B���?��%�IWЛ��"���ӂK&��.����@�UQ6KIZ����h�g�C}�'1u0p���=���ؠ�(�)\��4
_�����6��B�����N.<fO��w����y�c
��d�����C�fn��]!]iN���2�|!u�'�'��m<;���M�!\ i� ����ڽ^��BMI�{�fp���Q>(�wǋ��YƯdL��:REݷ6�Z"B�m�Q�WE��֡��Y�{X��!�͗@��U.��p����"'q�[�t�ey�z���%̶��6�n���W#�m] g[_��҈7n��̄o�n_)J�_�on|Eµ��fW�y�	V�3LԯIy�k��^�[֟,|Ϟtn�<�k���*��Ä;^As�]F1��hv���K�;.5C���G�a�oF� i��xt^�♎нU�hBx����J�m]_�ލ�h��	�j��[*m�*#��֙��5@V���R���#S3�&׋.���j��@� �)�߭�m��럧��6V2�]T��̥T�?MS�eG�_IZ�Y 26�%&�����΂~ТYδ����h2�*_"R�r�t��e�V�p�|�jg,���N��T�\&z^��O�2����c���i�CW8��͍U�W�w�/v��gG��[��ԑA�ՕTz�H�$�i�'��%��4c���3&��]!�&��4���<zF��u�e|;�]6t��FgY���+�����/�OY���R�m��ϕ�cLc�볅���24C���=IQ�Fl�i�f��e?��G�����Up@
=#s���0 asS��PO�_� ZX�υ�ƋHCBa�)�j_$�p��^�s���\L%��2�.�`f�����_����`�j�!���|�G��IBq��X���TX	��t��;�����tf�P�DD���s[��B�s�7 ��GP�f۪�ӓ��}��/�L��4mH�7g�]y�%���3�N��X���E������b�,��������Vn�HmS�5�U����]�$� ��Y���P�+�\M�Y�ѯ2� WK%G����Q�R�no��GGnW�G
� �������]��JҞ	�� �������B�br%6���Zf�y�'�p�]Gs�%��?���d� �v{��t�I��h�RbС2��6�����N�ڜ}�=bUc.'�>�؆`���}��~K��-�x�/X�d���o�1.���h�} �>/	N}3Ŵ����I��4�0&�{�!
�~��46����k����H!�d���:�G�,��"��\s�PH�SŎ>�����bϐ_�u�.�0�JĪ8�ЛÏI��\�f��X1
h�\����߭є����LY�I�H6�����Tsk.�)�O�RXitRF}��9�5��2�	��?<K`ԫu�'��E�潎��`ݐRV��w({,H���]C�Eɚ�%
l4��%u�ךd��F�ġ�x���g�$;�Ï4�3�}Ml���W~�wfE�i�0�����> A�k@��hR�Xx].t����8��-J���E>Fѻc}�Ǧ�q
��4eݙiE�\�*�����{�VSL�(Q�0��fX�XK'�j:�tz��JJ\Ѱ�w
^��{���[80Bh&��]��͕�͜������BV<γ�3���;�s�԰��Nw1�{�!�=�a����2�c��;��j�lʆM��}�j�lv� yB�d���!��������p7(�w��l��'�����rkM�`-�"R�H�̶���|[ ���1��@��X"���_�KPy	��+Gb�q�g�F}>�d�̿N´H�c��	���,�����n{h��������Z��T���'O��6�O���&k��J���
��.>Ѝ�3��$v�^z�DA�N@����nⳀ�Vs�ɛC�:���~	b*�y�P�= �߿������lS�sk]�k�;��pY�����q�K�I�/b#A��,&�
�z�ْ�%�s�U�偰�Є��X-��0Gst���ѡ�\5.:?��A�?dr�_0mb�I^��Q-�wҗ;QFD預I<���Ċ`Ng���U�M��d:1H(i�b������ ƪ��Ƥ��R.1uf10�A�Qt {X�<	T�?�UF��x��inc��'�����+J�O_BlL�Y��f8QJZ��=���y�ʮ\�s����%E�XY��cn�8޿�uF0�]���C�»� ������P�'�ޮF�H���k6��'�n�s��z�vl-�N՛l�ń���%�z�/T�ݾf��DEVÜ#z!F"�k@��(��D\���P9
���J��}����T^���#�P���t�\���d�����z�-�%N�_���o؅�A�Fl�>�[5��k��M��N�`,{>�@X�WIPw������!�K٬��젶�,�0����w3��6��x�Wj��)�'��<l0�\Z��dE�3b?�`�����Q��^��Q_}V������<:��
��>�za��S�CB�*�Vo���&Mp�h2����kC�RVo��|�����s�W�Ί�3�x��1kuՇ�`��$�ڮ�
�s�4��G0{B�)�8��?��v���q�R��O�[Y�i!-a�]|:��#A�֤��
b�]����C�_�^̶��?��ڥ����~V�f��8�e�P���q��x�[O+�	��	�O���F԰���
w)O^[�3�s���0A{)�w��'�O p��C�!~��i.�J���IB����`F5��p���<L���#�L^�<��I�׺�@7O0����%T�*bL��u-͵F-��(�g#�8���7�g�611H?�c>\�0Y��|d_�#(r��G�
>}�C�93i�7&������>J� B[z���K��T\����e�g�m�V���P�r:_��Id�2\i�|�a
�;ȝtx�i&���}�M� ѓ�J7K(T��z�']�-�}����%�1D�JI��3�'+�53q4�0���,�� �8eC��U�R��Hǁ�AnV<�"������B�ȒK�`�������*��ԫ��))�K��U�ќ�3�z��)H����'f���X������`aG��luP>��J����"��5���[{s�6;�^����:+�y5��+}�����S
4=�3U�]��{�Ķ�/����?���r
�V��W{4�Y�iRv�\d�ϒ�oZ�<�Y>V	�\
�B=�C��=�2���z�&���� X�c�	�$��w['����M����mi�q�6��\�ɇ���l����L�֗���sr&B������0Z�£>�M@�����Q�=�@̙�3�d����aPΊ �+w`�D ���5t�vÓ��O�m�

�T�,6bt�x��"�s�G����)�����;|�l��
�����IQ5�ե2�֕��~!7�G,V���.t�fn�x^!iգh
����/SEepao��-:�������p�ζ�x�L����Nj��ͣ�L^
A��!R��,��:�N@�X~J"�|⹎��0z���v��ކ�Lh�	^-��OcMA�.�"W�.��4��N���gC�na��]6�,~<���a�'"��Z�V��t�Z�!�T1<}�J��l�N���B&�1���O�8�ou�JXf9�4�c���W��������w��<�d9�:s�m�{�k\���MʍK#Lce�Đ5ǝ����<�� ��U���Fq�|`1�f+��M��蟠r7A���_r'�x
����5������kb= �s�jl��ԬY��+�1��*3�{�A���s�僧O%'��ce7牢Wֆ�,g��T�����ZaCE`�,o�l2��f�$Y�=����=C[I� ���V>�#^d�Z�ӄ�����8fܩ'jC���"�Mc�^�&U+��8�\�W�A��y�cJ$;\�k��������Z���J�+<$��,Z	���H]��#j��ݪ	���ĥ�-`5�u��+������/�f����㺔8z��Y�1T�ݠ�&�:�������tz�ix��oޑR~�eS�6�߀�9�wF@C^'|���/4?)q�3VPSWː3��<}�\�f�c�،jd0H�h����J���S �Ɠ�ȱ6}��~��i�Q֬�m�[��[
Z���}��v�&���*]���0�U|�4�-0 e�p��UR�a'���:�U3>�|b._#�̾��܄; d��ƠX�t�/a���9<�z0b$^�nhu׬N���*���.�|��m����d�%b���/��%�`�����FB�>NV�)�+nQam�M�H����w�E_6~dHY��]o����h+�
�
F�;�I0%��21����[���[�8��3�X�PH�$	��t��t ����槛j�jO{9�w|�~�E~��OC~���6<�9e)/�$T��5��m4=t`��W����|��B��@a�ĕB�':�i\xC����8�������m��h�Jf�^Ibª�m�:�E+C�Ea�5-��S�a����g�,k�V=���?�&K癆�H���5�3>�IL��6����x�5{���e�7�}t{�-�B#�ٱ�&)��}�p썥VD���$K}2<YU�y�[j�Rd��I}|�5^m���;�y����V6Ҽ�5�߽�N�D�F��z"d9��ۇS��͓���y̧(�P	cKg�j諐!f�p�K0u]k�9�f��"w� uDS��ٗ��@H����2�uˑ��<�1|�.�Oz["���/f�%],Z5��ѐ��3�|��#O1䔗����b���a�R������3ᔄ�,{e�͠�]����͔�O1j̘�?9p�tƈ�!�����ƶ��~h8�DTp�n��g#  N��D��u6WgIe��׉��,ѧj��M�yꅖE%��@n-�E��Y5��xO7q݉���[�|�v������ޞ�wҳ��&�B!����)>kZeSRB9� ����O�4�PD]0����M�?G��(�j�Q+���k��L�&�A��H`!�
���  �#
��d��SQ��>j��P��!������	_ӹ%ג�D~�?��r�(8������lOvcz��"�wlHٮ�h���[�⊼�Ή�j�$����V��$?���^f��{�%p���"���a3м�o��M��2�aE^�����^(c�
��̬���)�>t��[���֜�5q���؛k���5����zZ���j[�Ĺ�͚���Ħm=T��d���E�^��d:�	�j�uwnJ�I�����娶ӂj���v"�(G��9��/C��,���B2h����k�1��,�Ӿ��u�L�gJ�r�.��n�@~)�;��#���T���^�X"��?�\Lا��_%!?�$���^�p>[?'6��WE)@�ʔ�Pǰ��y�K���yk"4U;����h���*	,sZkt���M.�����;x=^ZbF����6�����y�(���\��uh��o�!"�K�Y䏷���a*t���v�kX<��Da�u�6�n-1b�A��L!o�H,�CKIX����6/��������d�y�Z��^�l_�;(|�r�`7u_�C$��3Z
/�9?�Y���h��#q�=e� ��A1Lk�^G7�c50fs3�o���:d����O�5��AܤO�����q�]<��n'�b���]�����3㸛<��|�t�w�o���Ī*��4��`�q�K<A�1���NN+�f�ۂ%ư�I���@�� [+0���@Off]�z�	Q̻�E���5�G�P��xlo�p�q��#�s�C7bP�!���\�6�^���3�F�+� =�v����S�E8���1��d)ڰ/�s.��˙����p|��7�0
��J[M7s����P���$�^'��leC�+����3�	��[b�g���Ӈ���B>x��1�cuUU��l�v�/���R{űQ����2�^tS}i���&	�5{��2]/�Z��
:G'l�_м��O�_N���.�D���`���%�mF����������U��M��/:�\��L��'����@1�n��~�q^]��),�Ct �H�r�K�m�}����(�^,V�.���|S���q�F����yg��Y��wzs寄@��{ek\�Uy�+E�P"��z0�N�N�_v:VZr�y!t 7Ns�6���.�*һ�"��2?��1n����k�WS��Hn�3��͆�:�*Dn�,�K�N^���wv��\��]K�3v���?���,������u�H7K��q8 8��B���Ӽ�(��gX��L�`w+���',��I��ˀ�[Ky9 �DS;gg"vӛ�p�:(��*�L���!��;U���x<1x^ ����z_bvƜ�T +8t^w:�Q:HgJ��h���"6�}��ڎ�f	�F�W�5lZ\��α��'�1�G	?��a���
PL����#�1�~V�!T����c�+ �3��怉�m�^ܿ֍;��:��&�˼�N�Q���a����Bv���q�k�[�zl�j� ����@{2i�"�ֻ�����e�S�x�DF�0�f�;�����K��{g�8���V�n��lF������M/��H�ҫ�G�R(��
�^�Q��JCb;v�J�73|Q@Y�1s��+N�n̞C�=Y��(���UrI���qp}�1�!q5�I")�F�,}p�YT��������Q��V�ľt�ѕe�L]ק�WnT�G\#%�66�}��
�Ȟ���]u6�ָL���2B%,���0I�)P�)�׃�D�-1z��2�V��jKa���Ľ�ʔL�/��q�%�������܁s�_���|�y);����7f��<K�É�tf���3�_�ཥ7��d��H�9p{��7Kf+�٭��u�պ[3���ʧIcx��%��/M)�K�y�2�����e���͞ �1���"B�ɻ;йL��� �m��:��0ͽ'�����$��g��/��S#�m
���Τ�c�t��
o���Qxv�y*�/�0W��h�r��n �y'�)����j|ʐ�_���P���W�)�Kf|���]�z�E�Q���Ψ�v�=���Xr	EC8o�$p<: �p�'��DU���`y��1'��n��HƼ�:�9������<V^��ݶ��A��E�潳E��i�+�F���%^s��U�zJ/&�`_+R�EQ�h�L���O���)�0�RMǐ�>�u
;&��!Ġfbj��,�ow*)ͽ֞>��/ɠ�tF$���.liiT������)k@IF�Q�<��TU���L�
�Jج{W�d�F�m��%�X�w�%���A��P-kן�w&]a�����K�Q�)�%��N�2�9ߨ2��`��CE��4h�bU��Lk�����?���;�\H��\�o�y�U�>��X�:���QM͞FUTu��u��i0n���������=��l�7Qw,�P3*���A�(R)�l��Yt�t�6D'\6��5�nf)�
�_奮�A?B�!�(ѹ��}�1�w.!�H��c���E����f�"�Na*L�6.4>tzb�1)	^q��@I&�ݨ{���7l�f_GA�ޕvXT�#����&�RH�a�w �A)�$Ê/+,�uvӏ�X2�ff�T�*zP����}�����f����Xx��#7�
9���/k����z͒����o����=����z�`�( �_���MM�Y��T��EX��2�f1Ի��]�@���H�_j�_�pJ�.C&αJ�r��^� r����6�.]���@��TRO��uʅȫ_;��\}�,Gz���N T�m^(V��Q���z\��9}6�6��U�ı
���mA��|�nf�0�T��)
t��c�De���x�%) 7(�k��\����P�̂�W�?�]'��+�xOHO$EC��L=F�L��6 )nsF~!���4�˷7c��:s6|�~�m�-���E�B\�4b���"�ޖEW\��v��j,�p�F7-�T�re@�l,�=A��*�QBī�~XC�	\[#��f)U1?��B�ݷ�?s,�i��W㪪��f�]���>O�� ��x�\M�np1%$�U
P7�����҈�eQ;�@.-��v�)���D��y��Ȯ��,S�s�,�_ Su���j��4&��ɥ6�xǭ0>�(:���'&��С��F��#^�
EHO�����*��	��br��@��b�q��G�۞�0љ,��ת^��:�{�̟�=P�C5+�o��`���η(��i0g}�B�_�炣G�0��w��?�	����(�"u�]�z�34K�\��7 �>�_j��[(|��M1�5��$ ˟_��F�(������ƹ\�R�͠�j�l�uĜ�����P>�́f����:#��_k�8^�5��������<�'��,�d|\��9u2ZDY�E�9�7�kȋ�R��a����Ȧe�:�9e��_M���®�w�:�.B��y�w�1��ol	l�xe��,r�`�(�]�Y���o�к��l����"��)^�7z>=nV�t��y��z|?$�����PoNCV�Ĥq�S&�A~��To������`�#e$2V��M�u�L�X^���em�f-��7����ٰJ�h���5��̮����͕F�o��տ��1|����ɻ�]��Czܕb��J�p�J�$U}��~)`���� ބ���V��nofxU�=���o	����b�c�p�X�!V�)�9�W�����)C�U8y�E����J����g�� ��N@�%οW�;/-ߴ���И*���Pc;��e��`YC!o���x��S�8��n0�i����>�֨q�=�C2�ែ� {a�{�� ׳�k�%q:��q�:�{�+��:���w;;�1�q�uȀ��tF��ZA�Q��ݹ� dvSI�O�u���i���Ь��ޡ,�"��l
l߀�@ʸ�v��v�~�_�~�����I(k�H�;�}��'�h2�^i������
`�	
ɦ ��6𞖼|���/�����u��o�x$�`;{ņK?�LL��EX��A ����OK Y�y�X�(��WJ矧�͌j�� ��:}f$����E��,��CzD���q�<��~!'����VZU3�I�L�m�	ւ{;�=l���ŕj�̈́�Y`��㼁5�HXP/R�������yR^���_���aV�7R�B��Muɩ-����ٔ���ٽ��>�-�#�GJ��2j��ŉ��6�G���P"0%�� �]S�M�f���W�L���7��A����j���KO��_��N����@�ˤ�E��\�ޤ�HJU��D�Z�X��P���s�fVA��v�\��K
�Ө�q�^��