��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��.�w�����K�F%�ͨsg�k�A����.�݈N$��_:.?���qi 3��**���p��&��D�.��^��j��!SӲΐ�h>�O����|���6��v�������R� e�<$���,+�*��Gc����L�W�(��^��'�0G�U�� Vj�)�bڅ�Mr�J�.$4qk�R�,��⛟���i��,Y���t�n��D3���k�~d���z�
h#M�{z�f���K9��d;�|τw�'�;��Pf� 瑈5{}�=< ��>]@g LŶ^�::�;vp�		�-[�����ܱ���w���2W���	{.z�gZ�a?����N���k/G~_R�A��j�8H���-Rh�x����5�DuPh�pK�{� :��C|ݡ�Eg�����(	Iű>���P��*h�Ż5�m���	��B����L�XƷ2v=/�u��,vLC�:�
�^��1�C��0י����(�n���GF秊�ꗷ�4�;t�x�� �I�a���-x���g���2�p;�.dG�kᆙv\�`�ܒr Z��8֕�vZO�>���#�^O�_��)�,�(��8���|�D��V�Rm�������Y���*���µ0��k�@�J�p�:V�</�cr���� �!r��.���b�"��A(�IZS>~÷����b��V�#�Eo�G��J�qT��#�!�Ȁ�7�A�2���+c_�[M^K>["��� C܎�=����#:�W����[T`����������=�^{xH��:�|V)Y�QW�&��oo~�/�����VV�����j�"'�����g�	q%4���+C4��FE@2�k�,`�M���$Ee�{}�b8��6#�By��P�w�m��Qܾ�%h��0�-)��R	V+� M���+��&�ؖyA�d���Yڶ�%��W�#�x0�S�J�U��Ы��3�&	V�R��,T���Hic��6,Lt%�w:3[{#j�6bm�1�w�(�J!}E�F� j{����=�1���[����S���&19�Y�p�xD����_�i'P�������3=1�j�LJ\a�T��2�~�)�\}����!/�m=�,��7����z���j�;*��#r���ۙ�� ]>"#����=�&�0��j惩�+��O��W���hj��>e��	F��*�^u��6>H �࠽�"�"o�| �r+�;f�J�l��}8+lZOT�����-B�`�޵��X\P��y�8��:�'m��2�0��p��/o����x�=�R^���~"�h�4�GW%0Ͱ�k�Z_:jI��Da|  ��Ӿ
H^�r��R��A*{��B�����J��֫�5V[*����I��b��k�Ϛ��%�LT���~8�8k?A@�#e��*�*��x�N���m��h�!�H�����Y�X�-X�WB�ZT�_6I�U�c��tVTf���y�p��!¤q	�������6��v������1�*��#�����4.�ү(��-of���n���鶦�}����EB[�	*S�``�� �f�H�@r���_�;y��+ @X��K��>�u����QY�Y8���"U���Py�@h$O5��	�]`�>�|<0Lx�4�ML�-é����ܓP�w�� �Y��uE.�c���}"V�C���L�J�"WJ���em:�զ�$H�]]��+6l���$�/~�~�����X:��W@$� ���&���2
>�T�]��������-bg9����ǔذ,I%H�컇zC)(^�>����ԑ=9X�KG�aY�nY��FW��m��!\���2J/�����K���8��c���<�d��I���NF�Ro7��D��1�6�WF9�u�)��gX�(�/o���8��>��%dB�y\Ĕ'��Ț�_�2�nBs�ۖ�vb�>��X����`��y��#�c�!q�Ϋ���f�1#WX%�[���(��ћS�y��z�.���FeJTKQ{ZcB���η�C]�Q�G�&��k�����5?-3@�����N���T���a��`d�2��Y�e��4�c$��2j��檎�`T��)��A?C2<\<]�u�"��������"���M��v|��9�c��O��x���B(]�C�ν�ʳ���������q��)^tB��m��/�<��1<3_������[M�/���~��a��c7�#��_)�K��y뚰5�3\{��0��]�.��,�ʵB*J�N���s�X7l	�1�P��A�:q7w
�,qzLl�������A���{�97���*�&J�
�s4�[�DQ�n7�Y������K�k�X�M���8ɻٍr��@E�RJzz��3��N솰�\ȫ����d�9�}�����=xQ�A>��*B��$�`�`ƮJ�?�W��*n,�LbD���#Oc��N�����=5�nh�^Eʅ�x�4�N�+�.�)���7$}�Ҏ�	i�%��$p��T�K��2���R�����D�iEn�O��@��2��� 6F�fS��R"�6����<.�Nv5O�6�r�S���a���Ve�N��_m�����
�m��[�3��u���2݈��cTl�u��uf�}�'����7�wǕ�+ ���Ń�q��!;_.n������B�`3E0�fє�˖��W>�9`#�r�e�Pi�"i�$(�~�/�Y{l��O?F��V�I��ۉO��_�!�f>
�R� �"ĳ<U ��0Hk ���T��pK7�5KG��
tSE�I�!PβxI���ߋZ����r�}��+�</C�4Ag��&��O������q b�^�-��ɾw>!�����Y���G(���$0�U���s�Lj@&�������g����!$ήNI��	��	{���[G���#��;qou�%���ׅ�j¥r���R�k�1OoH��7���_�l��q�����9Qx�,���V�[2�_�$$���p㽋�{2N�R7%�	�O����D��!�J����i"�{���_�����:dX� j��z��AU�fLfO_yXx��ޯ�os�m�ds�zF��W�%GF=Dkba7d��I5F�����E"Ĵ����x���z����<��r�a�.���ZR(��}�e�P�s9���N��r�����'�N�5��=;��%��E͗�r\��K2��������:p��0Y:U�$?�Cu��z��l\�BXk�^�1m�S�2ʤ���cؙ�����ĪQ�0Y�޹�9�m��g]W��?pV���=�M�_��W=��u�je��E[4fw��Bx\e��XlC)��ی5�]'��� #���g����M3��J৭�Z�B|�V�� T���*t�?'+_}R��َ����0W@k���OŦT�W�@��=����
+������	1(u�z����Ԛ�m;d�_��Y�܌֚.���Э�<��#��i������uA�U	;0xS����YW,=����ޗ��M��*k��m�[�i���y#Ζ�ņ�f56L}�Ǿ�\�]qɴ�0y�)�٧��x#}��k�Χ@��ص���-`a�݃(�G�s��d�^�|bX^.Pf��Ɠ�aw�z޳\x��k�yϨ#�Gz:$ɿ��;��p�ՉmZh9	���g��݉Xm���� ��\�n)�1Y�$�����i�U�&�0�� wV��%��ַ�2����p������'"'2%�9Yhz�����E-!Eq	�y��[�fR�*?����ݡ���ٝ�����.���Q�t�^�h�j �����(�L$�G��/�jP1�;k8`;��{]ӚB��D䇯�����7�T9�%nC�o$��Uq��%R��a]&"T����9s�N��h�	ܑ�egP���ZV��%۷=>��3qTE:B���AG�G[�$��z��7�~�=���~W�>%�Y\u�ʧ|
ƴ<�	]A�\q��%��ߪF�<���^<�M#��\	�{H��6���(�K��l@����FD��DMN�����j�4��Y��&�Dξd�t��8�Uк�7�Gz�?�bS���T�s
pE�+�ܾ���Z:t����V�������T)!�����}w�$[x�r�����z�،0�^�Կ� B�s�L��[:	�)h�q��j�\:5xz��D[~r��׿~w�f�zW�v �¼W��Pwu�p���D�����C���`�z~+������@��&G��-���~Rp�R)��ͽ�u���]"x�vج���{��۹�!^.�f���m�T!
���V̖3v��o]���´�3R�0���u��</c:�Q���
�	���NN��+�Qw�ۘ�Qw��@%�'�֮r�4�#]U9k�'ܒm����W���a���G�.=)p�.aJ�����f�#6������p�'c8:O��S�u�C�L�j�A�)�^	�v�������dM����e�+
5����'��R"��� ������[^�2�	��!M�۰��j(����O�^�%o	.�h1�\�6@�F�=���#5-V�$��H� ��bg�ץ�F�<���{����2p���:������f*[\�x�������4*��"8���*�&n��RP���M�i�R&����ݔj�O�`�3�?-�T��.�/4sq������h���߰G�D����ם|@;��K�.����n�V^8�g�0������<�9� {K: a)���l�V�7�ڴq���+=/�U��|�����>J3�ϹK�RV��C�0ly��L͉�6���P�1�Y��<�B-���>����ą���{{�U�a�az�I���$���	�fs�t-�S
�<v�L	��(Ax�{C�a��	t	��!<
�����E�%��';�Oِs�x��nξ����0D����nE^i��~�Ȧ���uE�Ve!�%���x�g:W�<�$GE:q�5�`~��ʓ�IL՚j�p��s��0�
�%��;�^����Dk7]��N��@�>Ŋ�h�or^>��i(��Պ�"I�������H]��4�Qa;D��Ң:��(#9:��6[���Dhe��\)lI�C�n/��0B��=|��^����ƽ��& ��9#����p�[Tb�fGX�c-�6�#�bT��aY���8�_Dn� l�3�PQ�f���3��qIl��A(3�$W@o������	�y?��tu*��^/kHU<�ܛ:�-�vP�6�v���!@`H*�+4h7C��Xj��TI����p]Ǘ�mҫ��+��#G㖷T�PsZQ-�Tݜ�PE}&��������>
�T-��ڊ� qJVg�����oTP�N��=+{p�#fv?���g[φ�U25TğQ����pZ���Ӷ�C0��	C�@u��ܳ�:"]��&�_�^���$�I���~~��K﮴�*�%ǀ���r��ڝ6Y�L�� I�.lG�M�	�V��4���\�O���{�m�Y.���F�z{4O�@*��ww0'�5Dw[Jﮌ)V��-���E����L�i8(���#�+81ݡѻ�yk���Β��R��Aq6�q���jٟ���C.�� ��ϩ�8زJI.��6���&�4;=~�ڷջ��
�Q$:�+�aD0�mP!��Ԭ�B#�Y�`2�'��V�0���eY��<'�14�e�.�����r�%Ryū��D��s��ţ�eg���t��O��`����׫�$�\���=5���X��������B?���O6Pkr'ktYΚ���n�����hj�+t�h]�7;R׳���~�?`��$��n�W*=R5l���{V������\��[�j�B�vB�-1r��(!V���x��]�
�+�$
R� ,9
�6�0?���FB�����M'<��Lj��k�n
�[V����V�5%
�fe��#�ѫ�x:�b�u$���:�]4���ZeR��@��ɢ�B��� K���(�QK[�� O���XS�����2��P���W��W��?��b)6òĨ<� <9�~ф������;������@�ɛ~X�0������Zb�M�Q���J,|%o)�g���%D6��ǎ�Y_�?�
td�l�N5ׅ*� �o�S݃h�Qvٻt]�6Z�ڠ�[�/6�m�Cɔo (���c������@�,�Yb6� �~{P_�F6��z)@D>x�����������MO��F!/0� ��7�y�}"zT�*��Ծ���T2�5��_�;j7��g���PRpD�Z���A/X�t�w��B��`�u�5I�
v(��B�����p�$,���31x�K�.ؾ���gIj�\1�������=C\��hw�������W�S���*ְ	��4^�t�������
?ŃM�K�\l����Y�NdQzj5��������"�����qZr�N�>3�?� �n�P�I<���4k�?�c���k9�3�>��I-�g-�ypR7�g��-�,ƴ
o���X���a�Z��P���wZ����bh���<a���	42�
��^z���~\��R���z?��؜���SaJ��c��������:�s#=��?�ٽjH`v���]����a1�	��M�y2գ�����]�$�v]p:�4E=���:\?#�A�.r�/`�Y��LU����yOIط�a��E�-�?��k��yɏ�#d�E�@���<T9�3�P�u���G�h�)�;ٚ>BHβ=���1�c��s���Bn���fhj�9Ac�h���ζ�$=DyEm�R��_t�Qn�;��'��� w��*9�h��LFxt�d�z}p� �1X+�����)�ԇ�Q�B��q�fB*bO�����s^X���I��K̻��ښ�:jH1o�2M.�_��N6,��k9ЩH�[O�/y[�Ց�N~�o�~�z�tfE
,�d�c|��{ �,Ӳa�?%X�ҧ��eW5��J��5}Sq^�ED��ey�u�p�]�$���I���{k�89���;ɕ6��h��8�D[C�>��||ٵ�ƂG|�qEDDG�u}����<P�e�d.1'lbd���S�k��@�;Fľ�3�1<���J)��J�*a�n��F�#����fYb����2MѮ�h�s�Җ@�6�;��sh#�j�a���b4c2AQa����q(A�aݐ�b'[L� �z�i��/�.�����O2ֳ��EUՏe�Ы����ac=��i�S�����X8+���!���z�	���XCN��b����&��Y(.j*Bs��&h"xh@f��5w�"
ú�D���5�V
R��"0=%P��3ʍ�Kݕ��}`���Z�^nǏ��x��MC����?����s�e��\l��o�]V	�H���p�o�H݌��=|�a�1#��ﺼ�,{�֋�]��j9	�1�
�4J�UbC��'����]�_��q��Xr���q��c�Y&�"����Q#2Gxmyl4#~��w�$ !# �s���9&\t�(I_�V�9�"����ȉ��c<Y�+�/l�mj[4Ax|<i���48L�e�q%����,T����#Y��~Oޔ�%�2�^sO�� 	�+����|����@$��_p�T{�������-����З��t-�$ŷ]��.�$���
e�:S_O���ʷބ����m/`���L9<��[*,>�,��?�~�
�U]�*c]ӠrX��j�PΟ�E�p?�s��Z�J�����P�Ify�>5�{<?Z���Զj[61Av^�M�����[:�H.���{m�QB6�v0��t��v�c�6۾I� �UMM�q��J����}�������)�̂H:������%��Y��}|���<��,9�nNO�H��)���/�ak�'LA���;@����׭���|o;]K��8I��iz�Ӷ���#�4e�0�=t��==GÆ�iA�2h�ö�l|5�t%������~�q�jt�UvS���0��e��lH�Ǟ��3:�ZC���<���d��fnn^�%��	���lZ!H��l��x�C�oU�(���z3>`����>S mӪ�~�F�|$�9�@.���I����B;�˧k������&�d�ۏl~KQ!x���Q��ˮ�=L�$�n$-W�7���D�FN=c�[{"�Z�l2��hώr�p���{�K��O'�� �p���;�zI�&�����V�*�<h�l%�~sd~�K�3� ɼŎ��2%V>���R��"��y;��y����{��������jY�Hj�\��8k��l*� ̃=r�D��|e�2d4�~��@~��U�\Ul�F?��6�����Z��@	��ŭ��k��d�9�P�/�|��	@Q�����$�š�ƶ,0������OIE@9KC�\������mɱ���y8��4CIV����8��W<韎oI?,���b m�+<��}�W+�������J�:VU�nc�"�9^�j��u�!0��A2�im�]!��:r�J~"�.���m������0���}d�Et�"���V3�ĥQ>��/�`��ۗ����z@�.��f܆�`d�ӯ2rة���2��;����!�Sv�a�^C^�45&@�����k"���Z�ێMxS�����|�ߕQ���VFe��)f}��;4P�C�"���o;�tkgO?�c-3��rbo�g�d��|?J�g�φ�̩�?�"�J�d�U�F3B�G���[@9���/҃<$��|�p�Y)v.\8��ϔ�o\8��a6�^O�2��:��7i�n�!]���M�;P#��W}���?F0A��7�~�{�8���G�Ķ�����p3xޠ=w���}�����=gK�S�nm1��?h:3��)f���A�i��{�a�����6,ސ	�	Āt�����h0^��bͅk���ya*j̀8�S����!��D�Ϩ/�����#6��:�s�>��!��P2�W�D}���.ô��g7��a	��E��-CCm����.y�S=�M�6w+FB��;�II��mb��-�Ltr�\ʤ~��J1
U޳Ւ
��.�� k)E&T���+��o��w���
�Ҝ�*��c�5�+�����i0�V�24X+�����s��LѼ�Ǌ�;_��Ρп!����k�RΏ鯗K�Oݳ� _,�(�0��
 2�d�Pg��L��=t����å���_%f�VHZ�������9�����d��]���`�����ԉ���	�H��Z��op�4�34�pǩ��fD4^�	
R(qҖzD�N�"����"��Q�,�D�n>R�XI�?�Yl }KB~U�=]M��6͢���F����݁8:���ιԷ��(��m%����;�d�B��A����g/��*i����Ʋ�����}�0	#{ ��]L9LE��jx����k�M1�c���~���w���K����Z��ӿs�����5���'u�c�P����ϰ��]���0�������5�Xu���l�4��n����չ��Q}����G;T�.��t.�ⰲ:�F���室0����`���(��{�ʾ���!���"�v2`�۶oDۏ��cz$�7:a�4>��e��
F���?�kwXZ��O)/".���0��r���ޓ	���X�����	l:��p�g�&YY2�d�:"ě.ɔH���{s!yX.l!�����^|�i�.���<�̝�L�0�<5�	u`�53���Е��R��bV����Ix$���w���N�#�hl�'���o	��{����M����K�-l+�X��u#���:;N[$Vp��ځa�v��=���1�/O:�������ƒ��k��C�j�'=(����f�U�f��;� �l6�W���n�~�j.��.${g�#��ќGb�=�G$��-�����|/��2=ӄ�S�U��x��W�ŉ(=9ǲcᬯ!Ϳj
=|[�i�K/�Bk���_w��J.�J�oc��u�W��u����_D��k���A�u��m�X�}��(9tg�:��nPp|����^�zsO�M1���CݽU�(��x��䥭
�B���8��ȑu}k�z�"���c`�s�A��?�4�r%���d����_w8x%!3Cp�zu���<�O@-��3zc�	$Dizݪ8�����`�i)_5R�|rQ>��$aO^I�0���x��S�V�&��ٴ�=L1����O?��%c)�Gw�^r�]�
NϿm�lq�0�E#r�Wbפ����}w�;�7<D �B���+=ֵ͐p���q��l�I���:+"8Iy�?s�A>���Jam!?����<גw�����OO��?��$#�2"[ �����=��OQ�Z;��NU�c�1��_���<,]��Od	��4By�OY�^�H��|����жJ�
�8�@�|0R�R�� S)n�d�8���A�ę�;D��[]�@hLy9YܩU �ED�k����e��|9�����mY;�ԫ=�6�0����J Hk��=�*e�p�;w-E��߅/O��=�R��	J�h���l��u\���`hZ��9�E
����ģ
��	_��D�k���a�� ������ً�� ��Ni�k�*�>l�iC�?%���ھ��Qq�X��d�܉�?�k��]/SC"�Vj����>�a�o&�j˙߆_�[�j\���o��HNܸ2�c�%y�X	���MR2[�Ŵ_U����g��ߘI߱E4�`j���G�Q+vdަu���}����tF�׋e�MQjZ�"ѫd�q��Jv�$7>�ĵ3�}L�=%���5��?@�3+4�#m)����1��4�l��j$K��r�C��V�c�\��D�ڡ�?	���%S�s�#��>����a���L��0��,}/_o=��[���CJ�)�ǇZ��i����V��i���ҲvFK�����7�:�xG͆�X��
U��]��df�܇vXn�F�R��q�N��ou�vxdf!n0+�g�clq�������Ǒ���IDo�eԅiO�����Iz��	������v�}���iY��%(�Y���"��i�����lt_�{v��r�X�g�Qc����XyK��椫���R#wIW���"�87��N�[��@ʱ�$�`.��Y����3���	��ݠ�.0s~��K #m�
z�mf��Z�Ȗ��F�Z���O�ݥ�P��q�y��~aQjk���<���-�L1�b蠶{o]7ސz|됪Bc�^�2�Ť"����t��@�|�����V��2q>���O��׬6��|��!���tL���U�-D֔�b�T��0֑N��Їc{C��%��ZVã�U[6D��B������4S��_||ȡ&��!���z�2lP��H�ې���_�d)�U�<�����0xuE��6����������@i�7�ؽ�-[��_�I-� �6;c�0%=u	/��~B��B�����Q�i�_�@r�_̹�O����3F�_��V�6ʦ���ErG��1����Y���߄4O���?ǂ��*[bIpT3NSF�僗�-+�m�@ ����|��s@=�zJ�9
^]���J�1vՇ��2Z�:ھ�է��v��}�I�鶩_�I���S<n��ϐ�����H�X9ȫC�P���ע���s:m@�6��9ȟrÚ��B+��������ԕ�%����ؾ2U]3��-�JĮ���~H]c���[T�����7��J�Iz�_����-ޱ�E��M"�P(;��@d���Q���@�j��?��R:�/���P�W�t�H�EG�k�C����<{��|Jg'�$����5%�X���P�p̑>k��D�UZ2����{d��Q��xdp�k�,N%��d�0��ۮ/n���`d���E��v��e� L�1f�W	�P��I:2g����"�fw(�F�%�$�?.��	�� �[r�W�ںbٳ��+y.�'��3��(����4�֙��я%�شt�n�7�G���4P�m ��=���kW�a�E��dU��@$9��z���S^���[��|�M~	���!�Wp���8Y�����=�-�âOw4xP(�o�͸�Tgּ���5�j�|�}q���������y����Z��]�!��)X��dA��,�p|�����xǂG����z�}$
���׳���F�G{{A���l��������.�����Պ�OnK���ֆ�:G^�U���d>Z1��"���ܚ��S��a=X"X��f��d>�t���6�=��,,�I�c���aܦ�j��h��
���E�4|ϋ�Ң�%U�S���E5����+��>�G�j� uj�a3�]�H�m[s���f}��_�,Vs�7r��nCz>	��W�1L���#����v�~���e�(��P�a�_O��-�u�U�	ڗL|�N����A<U�yraM!aə�����J�w�~�A�r�� �O�6
B�f�;,0靇��W�A.��֞�yi�����9���_�!.9-��dva� 4�'3�C[��}p���`N����b[�&�xG�ܙF߂N'54R��ꤧQ��9Լ�1"��7,f]m$N��/��\Q/�WA`S���F�+�z�"�.ʹ{�/Z�v0��~�B�x�	��eR���J����m �.Ht���	��?N��R>lW�JC_@p���.�q�u�I���{�ݖ�Q��Y���M����ZJCǼ��e%1J��Z{!bĭ�A҆�5����MEư�lpI��K�z���Y��D
K8>����5�t�"0J:v>f��x�Q:S�Caa�x�9�9cX�pdTG�\�"�3�X��|���Vӭ2E6olg	���V��g�<���z��@����@q=B�.��j��=����A�i��`l���l��K%�h�~ȺY�����?,��*N￬��A��E�#��u�p-Y��O�U[*�I����̎����Ϲ�ڴ;ĭ��{�Lh�/:;	������@Y�9����� �]#�#H��(��͹"���F���zkG�w�b����}"YZ��j��S��e�|��`_�u���n!��+��/�h
L�o�O����c���;h�:J)_�L�\��,��t_�O8OF-^��q���["�A��֢�̐4D �<���!/.29M���>�N8�2y�\y��_
�]��;�~��ݶ�&�6钪f偞�wX�@tE�Li	ΣD�"�G�,����J���O=�]r��Pj���v����z�!mբ��`e¨d����!�_`�~5ؓ�A;����C�-$�ot�5	�!�A����0�����}�	�-OD_T�C
|�(���]�p�}B�����ju���gj�En���C.�?�r�$�ږK�-�2;�j6{�a�{8�����F�Ȼuѳ>�)�_:u���J�&B�6�F4��5f�w�'O��)��Up���CV6@;Hh�g3��a�;%-���D. 9�S�ޠl��N�����,�6�*V,�fn+S��z�y���A����G��R v}�?%ݦ�0}�h��sTS�������/�S�
��� ���-�{:.P)2���߂M��������5Չ�կ���Iq{�o�K��V�ZGi���1�ޢÎ��J��*�i�B�������^5�T��$=��bd�ț(6��َ/h�p D�O\�? �����n�IRc
��Bc�J������bhH1=ORV�u����=x�LVg%���Fe�_�kq[��)t���Q����X0��=IEnǉQ�[y(�_!�:�Ƣ���vd����{6A��x�����'�����%�̼��Q�6.�I��6��^� �{Y��ޘ�]��㕣��5���v�,\%���;}��ַŉA~���!�{A&��n��l��M9�u�l֓��W�Xn�DZ+����?��_��E��B%�~?��Z�C�U�:��w0%�KÀ1�=�b��8
m����h?ދ���̿=��q��]��8_g��>�����"�n*=���C�)�t4�;�4sqkA��pB���{6KE�fD�p+G��5�^b����2�ɔ�H�t�����ciݚ��I�G�ӖH�S�!m`�4N+Xoe �訔{&X�f� ���J��಻�Z���ZB7P|Ol��i�=Ѫ�)�]D�V��n��J�=cҖ�{�΃Z��+��\ĀoӤ�}����؀���t�<^�rI�pn��`��5)54a��Es�8Q�Jw,@t(���%��	�Pe�eH��� _��Т �$}�܉DGF�$>��&|�}R�.�^UϦ�^���sƈ}��Ά�:
?[��� p��l�ު�%��,=lp��,��5a��iN��в�ԓ�`�6�E��!�{\&��F��C��ғGe���\�G�C�ȥ%��-#ll8��V�͟v�!�ђ��!���VS�q���`F2M���@w{�x:�)^R�>�(��إ>JyНF�[;���1z����:�^����6�	�c~�mU�NF�j�����S�z*@ac� �~�R�ם�$��a�?������Y_v���77�WT�&K��~�6=�3D�QԺ�!L�\Y��m|�*���ȼEQܢ�����4��:��`�0�X�-�4���q��Ɲi�1��+!�9�#��@`�UՔ�D1	V�O\�NJЯ=RJ�ɵ ���ȭb�1��I*����s	��]ҀZi�F�3�0y�V�w�БE�\Q���������(�j�f<��A��u�W�S��6�SA�i�g�������#e<���%!�q�/b~��+w�|���~!�#���#S���>���]u�z"ĸ���[������/Ɲ$s�c�~�Ε�(��u�h��H��2�2�E����)t[
a�������ū����X?Y��ʶ���]fi4i����.����� �wF��3�5��,{'j�5�Զ����E��B�A.��콜�w��Mn��O3��Xp�wG���}�Û�."uI�ʄ�w������V�.'�gRV[op�������HSv1�Ƭ�*ۺ�%-k��
}�B��r�}�C�H�]�ԓ�wh��yG�R�RIR1�{�DDB���U�VK��
�o��log��l���xyZ�w��ѷ٬8����w|&&���O�İW�,�>?# G8�+
y�K�w~�{�p���&A�"��2�����\F;b'�ؚ��������.��:m{���z8E(X|�1�+�P-�r��\�ĥHl�!���Y@� |�r����׫�yX��&dJb�K�	x���!��]ݟ����ai����>�$�R���E��,o��Ŧ
�a�}鍜�Rh{A&��ȣ]�[��:ŕ �fㄨ�E+�w[c���>׀�_XvȂC;~I�ψek���Z������|��_u}g�Wk�<��{d�Ǟ�9���>Q{�Է	m�w����G�A�ռa��C�.%�S=b7h��"ʡ6]�o���n��L鮞�`�E�K"��n3�j�U���m��n8�Ux,���KזK��K�P���.R�:"�%��K��<��������)-�o�ʛZ�vQ\3�� �a�'!w�����m-�����K��ߒ)�\�}l��=���u~n�i���P�����Yg�7ɒ��x��3�)��|A�������mC~S���U�ؕ��.ʙQ�|jzr��� �������T�q��'��fG%�Iy�k,��1��žc6�K!�$W8�wM���n�u,�6'�D/��~J8'{X/l�ofsQ�|(NN9oK��K��_�ӱg�u1��j�����O���������Js����h�G��E�����z#�Z�mG@��x����1�-�.��
��������{~U��w�j�$;er]�%�ۮ�C�c�/&���HbM��թ����B'���v�xz��A	�aC��}�̴�(���0��^NQ�F-9����ֈH,��[D?�dN$��#�a�n��������99�!+_-v�ALyT>{
�s_�S
�_1݊j
Nȟ���>�g��Uإ�ɝ�c���	[~pr�d��2��a���P�t%�c����
�Q��N�i��xNx�Ư�tZ 6��(�f5�Q��⭾���/��,�8m-�T96��V�=��.M�~f]�=�Ͽ�����W)3�3�,2�|�_�H�v�w>�����7h��t����i	���b��b����$��N�e�v��Q��M�"G~���	�����ڛ��B"��:��U��Y��	 s�K�b]�8�hs4ib�?��L��oI���vB3�5��Z��z�%̸�S)�"���i���*)���TJ`�O�k����� 8��"׍r5�8��g�&8N�[���.��X���_�+�L'�"��o/[��/0ҮmJ�ߝLS�kt0Ƥ9C��� M�αU��͝���ޘ~��3��t��}�g>�J�@̂�r3eb	A�[zy�uo/ �b���"+�! ��[Uw?L���(t��TDWvI_a�?�3AK�p�-H��T��G���h��+��
y�2�������Խ�|������9Lju�$k��.]�h�Qe0t����U���n�b����h�e�w�6���i#:V~�X	�~���l����x˼-V�'z�����D�C~RT1�x9�Į�.�*
Wg���d�@9��!�Q���{�U� ߯[Ӊn]����.����$,���ŇQ���s�#�7�%���^����Fy�S\D�r�=U�.r��5��8��G����<,!8��'�3G縄��KX�N�$��i?� lY�����ɖ�=��3[�8{�B�H��u��P���m�ӶRY�j%P������'*lϱu�����/�nU��f�R��]k�\m�־��!'�S�7~�Ź.�ctRB)2d�iUܯ��u����I9|�p����c*��jZ��>�euP/6h{U��	������4���<w��j�&̑"��gpE�q���0Gg�5���b	/����5&��/������)ia4�V	:+�|4��� R���7y$��i��'͆��(�6��#��A�b$נg�=�w�As�F��������+�V$�H����U%�?�^yˊ�N�2��ޗ���5�/�We���b�R�XF��·��ez�}���\�fR*SL(�=�)���@���''�[p>��eGC����f��c]Gȟ���ˈ�� �9c�z�"^0BN�dїF���#�@^����wd�_�IaE^�� �{nS@�z�̣lC���#ံhp��������
H\(|� ]����5�}׶�M���(ż4قu��zȅ�N'��א#�����/�V�#���ڡ�#uwl�-��]-$��W=GC��3m�l�f�jɏAݵ�:&���,��u�o������FGN��>�y�<ۛSGn��۾�vAь�p�e!���O��׊-��U�~-���#R�Ѿ��?4�bu_y�Q>I!$�:�ֱ����ci&������&�{�CR����
�\b>F�L�N'���E�8�s9 b3��Դ��M�'�%E�D'N���@�5�w��7pNL`�,��{���`RQ^&�{�M�g}S����cbOk�
��Fe��2?r"�x���)���ֶm�5��J�//d�)��^hR�X�P^�������g���L��J��/���E�|����0="�:�8��џ0R��7���%1iۂm����1�=�2GF5��5��f�g8Y�ti��x�:����D`���a�r�
�@�w�Bc���4j�+,��$TC^˷ZS�89��ST����ۙ�A���E� �u}�[4�?��0t�zM�}�u/�9�af��!B�����`JЌ���I�������c�JRV�3ִL��xH��o ��Eȫ�gGA^��i��d�7?�O����T��O�/��5
P];��`qq�ƕ?k�l.��rYk���95�nH܎zp��Lmֆ!�c��]�^`�|��� �;��>u1fo٘�׳"�� K�Y���H�T�
����Ԑ��*��~e&�+�E48�:;�2���O*�I {��>�ˢz���dw�䗹G�f�`��N)�Q�>�Th+aR�򚼨��bi;F�����	7|���2DJ�4>w��l�vفJ�qv ����9�$��߸w/��y
!��Tj� �cA��IN��ao��C�r?,vk��:��M0�e���L��	i���w2��iH��](�_{]ۜUW�=���]~��o9��#/a �J�p��r��sw���Q䦣��۳W����7t�; p@��EJ���Ēw�
�?(dRU��K��P3ZȌq��C����v��3��ˁ�pѽ��3���*Κ-����
�O7:dQ]�0ŋq�\��C��
�����
�溑�뺶�8��p���Ye�qZ���g�(䇶��=�f��V�Q Q�~3N���t��Qz�.�VZOPݪ(+Z�DC%������ȷJ��,(-���R5O4� ��u\I_QK)v� �8%!�O#���7(_ĝɅN`�:y)ɛo5�w�%Y]�����Kxyb��s�yiObu�g���d���A��j��a�	����tdr��z����S:�?���� /n�5���h;�<k�־�n-�'�s���Iw���-��[�RWq�Y��o,vtcU��ɶW��Rb�ZO�.�>2z�E0�{�
L��:�c���ܤ35H�r���4�2�|�+���PF��l�OGo	�ɰ���a��|��7H��Y.��q/��u��З(�8�� -�ɟ�{�ڼ�؇�G�0,.j�x���Z8aB9�&�?9-�����(+ͯ�BPv�:67��z�<��bI�U��E��hOy��	{2�V��bUhg`\t��+p��-����.�-,��Ȍ�|���VLX��Fig�)���Ƞ#09)��T�4񯰅^Mld���\���F�������һYnj��(���v��0aY���L�R��W�T�]K�J 2���Qj�$x�|�ȶ��=i\���t�RRbP6�AO��EG7]�=��N߱�qw�K��@�ҝ�XO��V��^��`����"�/�#�o��������1���o���Ǻ���C��X@6�K����=��P�p�U�C����/��N0^�^<f�~+;��$��8�IlH�M�5�!b�*a<0;����"�:.g{�rz���Sy���!d/�q�Kz�M�!'�7��(����=_ԛX �|�Y����n}5���|�y�����tw`B��B���f@
�@����j��|��j�(7�����sU`�}Ae}d�����f�\�?$���czG�P҇��OK�/���p�|c�o,�PD���+���W�����D$�>g��hTu�Wޕg|X��>�9�4<��J�;�j{��~Qh�<A����3ג�c��6���N3��y�e�R[�#1�!��KD/$�UE�F�����Wa�ē�ю)Os��EV,�oQ���- 
㷴�����1���˙:$	(Y�w8����@�C�2�oZ��%���s3G��9C�i�}CȪE�ɼ`h�q�F��ћ4fpSБ����i@(�v���3{3�\@< �zT��6x�f,�Q=�S�Z!�c�=�E�,m -U�Ʊ�  ����-�)�d�/)����*���5��������$��{!i��"��n�O8���z��
���},~�#����9��+`�_:ȕQ�?��izc�������l:�ƥ��2 ���z8w9��a�0�����Ԏ�=J凂�I<���,�e�3���e��8�ˮ��9kY���������O�+;u����v)n
А�P�,�%�#�t�tƮ�D�8vCG�
P +E#^l�,��b�r�UQ}5�z@��#lZ�!�0��M� �Ϧ��k����N�'C;Q���:
&��u�&h����2�\�'��H:~g*,���9�L��^�Y=Ff��M�/Z�]>|}>@VE|�F��F��K�����S	FP��1E��WN�ֱ����T�e=�B	t�0�zӚn�x M]��nr��MV���g�F� ՠ�l6��`: ���u�#��i[*Ӿ n�z��A�(�����"g_�+���G���v��\���Ħ��#���S��>��t����=�6�qIa�w�X�6��q̳~�[j�TGx)��g���/V��E}"����E���0��e ��ݗH��o�f<r��A�Y.��z���w0(Np���yo�;�o�j���8�ۜ �^�a`o��~M4������ߩ�	�2�"^�f<7Զ|I�x���]>%��V��#b��cٷ���
��-Ug���6f˰!
�'NlIȼ���X?�H�hu���A�j^zk��<�4f����t�Q6�He�7^��ҹ<�ڑC�]��8�?�("��p,�����܋JnC-�Y߼�U6��Y�>\�$+Q}>=��m�����H)��ןF�mR��^@s�{�'o}��������})/fP��ũ���Ɨ�q��@E�-��A����S2c�mW��K�F����J�z�0HD�!�G��
,��� ���=�!�c8:�$N�X�K�X���6��%��Yr\J�_����} ��3f�q�*��[�{?��luF-��
o����a�y=���G�Ԉ��n�%�P6}����u�H�uh���H|I/w'�K;b"��yK�˺���u�*(_]J�<�m�)V�Q�6t�<��6hvU�~f�i�HC�,�V�A;�)�#��nҢ\���]�D�nP�R�R0��y=�;V�FdY*z�	^�ISk�ւ�/[��#'c�ܳ��o&�JHz������a��OAy��<zh29xfL��cSY����ʵ�G�D�yH�W��a,�C3��)�+�U|Dpa�tO�=h�ʴ������H�z�C�d~��3��q�x���B��n��L�<��uf��i�x�K^돒���r��1�S�k����f��4 _���}�x�������/|��fv}-�������^7�@z��=Z�jE9=�>��C`���i��7�#���]t�
00�#�ܤ6������G����YΘݹ<�c����:ލgS��^�QJ&�"��z(����[���� �Ǡ�V Jh'�ݒ��i�*e��[\�8���XsI�Z�Rq<����ɯ��ah`"�����GR��A�����gܒ�lQ�*�_�zaȿ����f���PT�{!�j(W��n�J�0���=W�g��8q��|	Ȍ�D���=T�Q���`��J�W���!?8<�o�7����%�o�RV����\��!M���ل����V����T��	���n�����Ȑ_L�AD�j������=���2��웾����4�
������#?���w�����S��nvWn-"{ 60��M�%�Oh[�t>�-A�Q�k(,�N����66s;\h��F��*���1�a�i��y�?�����(Y6;�҃@`��W����p�*ۗ�{�j��7�� �|C���������w*۵�;r�E�b\-�S�H��_!��h�� _0���T>)$��^#^�#�H����.§�{�7�A�Bj�{�ɡ6�A�Bژ�LȬɋ�`EQ����2���?�f>q�|��p����Y�o�̛ZO��$)��nU�Q� D�!P�W���$���b��̐�}A����}�{8�i:�"�����i+�*�m��0��z�M/�y����:�\Jպ|J���E�9�7z&E>��娽���V����OM�X���?s�~��,^^@ kKh�_Aܭ� 6�����X�us� �pG.�TC�׎^�������)]��uO]�A�[� hs��1=A��$L��u��n�~7�b��N�f�q8{�����AdPZS�H�"�d�����Л�tś&u��T�R�����s��Rz`hH��еH�rr�+KL��*���m'����� �W*������<��IvA���]��x�n)Ir��o����t�XM(����ʹٵ�'pO]�8�-���-����E�IK�^��;+���<�rv�]���xY�Mxm������v�?���Dg�㌸m�_f��
�ּ>m{"J�"���g�۟�?X��/ۼ�E2�+ ��Ђ�~B9-���t�~ʸ�P����0�b���+0��a��5N���H��xٝ�M�L���Z~�W6��P�����P�@1N�2����Q3$�į�-B�}6�ЀA�Τ������"���s��dE�O��`O�he'��,����f �����TKtww�1����g��a�}�m~��1���	+���i1J�		l5J�'�6b��� A��B-v@1�r��1���~�kmߞ�%�i/u�,�A��j�"���x�TA����33�7�f�;��q��[��S����6Y����Ҧ�(���H�9(y�О��D�ٷ�9��	Y_�D7���|[:
����tX����~e4X*94+��\B�A;F��2πªژ������&b;�S~ Ɔ���g����喚^�¶`ۚ�b&ʮ����[F;>b��M�]���9B��aD<�7�����๫��?�BL��* �*�f�ڝYb�N��Qr�5RoV�&l�_E�_�فt���<��
��էQ�?�׽�p����q���:2���9�\��8դ�m�����*���W�FR���s���z�D�+t1;�/���C�����o��I��7+�s�����7�D;��f��L�.�P�Ӑ}�+ҩjs6h)�۽~uZ-l	OeD}/*^�) l�9�/����r�\���*?�7;+�OlI�L��:'�l�i����vpY��ϸO��`��+���yb"A85='&N+إV�KKG.��d��0����V�mqp�)�H�A3}���yھF f�J:SB��/� �%��l6^{"�<�w��ZDmE���ҧT~tQ��nO`ԃ�1�"Q&I��iH����u"D2Lp�N �\D�=��w>����8�|��t'�J$�c��s��
�'��\���l_]C�͛�4��{���ӄ����8T�MuW�خ׿��A\�m�U��^�ܥ�qM�7�������f4�/��=���wYjD���Y�B����'
�w8�WT�n��Z�V��3�l��%G��ObF�,�.VT���ˠX��X��<.����k��
�Fe��o�]5w\��d��7�/@pK J]��:�$�6��/k���P��{�D�[��&�g yP�}�P����(�v����I��[�
����l�Ȉ˽�_��V8�sF#�S����	ײ���x�z�JJB���N�3��m�g��H38v��7]�/�#@5����mD���r�b�����+�pt����P`o�����j&S>�1��E=}�QA��g����6�z�r��c���w ��dȸsl6	=�w�е�Mxi�s��eo P��㈈,�{0>���I�5�L�����q��6���m0V�x|�BE�C��3��a�_6�r�.;!%�^IJ_-�/�������!~WI5�O���W����	|q�ug@7ƣ���Y󝃜l-�F�#����m���Z3���ļ��g��M��?��<��W������W@9R��UF0y��B�#W�������t��^(��Pq[5�	��<�}z�ޑ^�) ,?���-�м��.9��3���J�Q��B�l ��NX�r1��?4�'TN��R� ҈��0m����O �I�s+�0����Eb+D>��/����,97Q�Y7�W�JA�#!Z�-�5�AA�/vsͅI^5NT$�Iߺ�I�g�~�,N\�'.�$ `��kXs)�S&F�{�F��GcU��H�A���/����H/�ѳr�^A����Ϙ�2�w�r���o�γ��¢i���lc��UfH��~��Y���.i����F��Jh.4X�#�����AT��cF_�9Y�ο���:��3{ID_̸D[�aI�k�專6<����i���b
.�D��l�i�!=���n�:<�P�ѧ�c���V�:���G�����	jepg`0ש��`�(�ҌZ��ꂶ����8��|���="�����?U0m��j�k#�r���$k�K3�]o�T��dF�W�����Su<���Մ{�'�>=�\�������
Eb��N��s�;�sO �@ ��� #�h6���[t�}��n�/�y�+UWڪyx��2��h�9L�P�Wo֦K�00�"����&�4��h�v��5L�䧵�~w�l�m�rL�|��.��"�I!�`������l�]m���,޾]�>Ĵy�F)�k;׊urV��J��4L�1��?�5�4N?U.Ωd�����Rn�Xu	�L�"��I}�}�����p��u����[���tq�^�� ���Cv�bU�pS�8�r����OM|��oj�@[�ֺǹ*�03�u�ک�ę鍬^� K���o/_Q�x��Q�g�R�s����`��+T;���K���fD��q 	�r��|��9ǁ��ܯE'8�i�%�j3I	,/,�pMc��Ђ��V�Μa��\m`��@�ʳ��9�
o4�C�����1���ޫ]�y�I�eخ,��D�vuv���-��߹	�[o ��!6ȧ*�(�o� �:?��z|堚���Z�O������:��2�R.�	�Yj0���w������ s�<��"�b�@�[+ˣ�w�o;FW�.5c�@$de�ۮ.�W!�����λ��"!���z�/Gz*��/����|h�Y�EM
�Gl4��m�^���?��F������&����u0�_}z`�=<b�ٵ@eO��-�*��ý*a�dU�f
f���x������Q��ԯ*r�P�l+ֿ�
w�*9�[�E.\�e
$�O-�Q�vC(�;��Wj�B�S�0:8+UFl/q�FQ�5�|���N�A�K�4y����s��_� ��R��D�؈��{E��h$�=�W��^=�)o��+��s����:�S4����i���8}֜�&Z� 	f!\̈U�PX�pm�t���߼ux�M��d�<�9_R��M>�,����S]'+�96���>#�E������:U��~�\�>e�xw��I�����?���tSŶ�m�wZ�?�������ZM�f4=D�GT9/���>�lf<BW�8��W�p�V��>w��f
i+@/_>�p�%s\S� �U���*@r^���a�`H�ȰL�n�ܲ?C�X3i^�'ggH���|�G�4P&��x��^�P ��OV4q�_$m��3��3�g5�MغGRwʧU�W�Z��E.a{jU�F�ֱ���EQvj��ظ�W�ſ�ı�K64UM��}����������k4�g,�ev�%���_!��%�6�{�)�V���8^��4_-m�{b�*������P�:�$K(��HJC�d�"��*��Ԟ)z�8���?�$������w���ݱ�@��1������C�ph/��龧_�}e�<̆��1����P}q�V�O#"�*N)��$8�F9ID�ƻ@��Aq�t���]3�ZH8��$k�`�RO�t�{����;�����IC�:@��=GFs�o_�Ŋ���+��s S�z�\��3��I��~���T����{�LݧN1��OtS8!����C���O���.l�P�����+A1�q�\9�&�bI!���M�	�+���F�e����vd�NL���Ȥj���jɟ�D�Xu���`�`�W(p@����"�q�Kl�x1<���3�S?*h�7�����w5��ymh�#�����̮X�q�#�`����ҾN��,	7���aM�P�Ҷ���1σ�R4hxU���45q��M���>@�>�dwwYy��7�6S����+*st=�m0��LA�w��GON�N��s�׼�f�O
��6-�mɇU�੯,Z�Ŋ(��t��ďf����#���.�����JUt�-H;�f@a?�q�����w����љ�A������f��D��M)��|�k���n�q8U��[��؂�\J��y)����������B��q��5�p���ʧs��p�O�k�o$̯v�;DC檄��s<#:�xS㌺ ��6��6�vSS�=��	�mJ�ԟB�q
�G�F��F�`��j#'��آ_�k3u>��0/C�Șuh6/l����14���حd4��qޣ����9����qL��/�@��Q������p�J̠�O��Z�M%�����#���A]۴���F>�+L��sH��`&��>,k$����=��*�^YG�Ԩ6�@X]�K�'��A�5�{�5������hV����/L"7�k�Hw�ȡ�����_��w��7�x甋k|g��I06���',���Y�<zﲨ�MS̒��8D	�I��K��_ "�ӗ������˶��%���ޣ�.����ͅxjs�~/��(r+!0�n���](c&�^x�}JUg�)@��ƂC���vۜ�@�=�F�u%�9u��O̘̽����*:�~�`�7O�����S�I���?�e#oS�_�W"�I)�5h�7��w��P��s	�SgbV�uH
*)A\�Wk$~�R;��Y�����R������0^+��B��4�5OGC �y�5C�*�$�����(]y`�mϚ��;��uU�mGM�ሸ|l��O
z�	_������H��4�4-��F A��G�����V�!@��s�/c3U	�!) O�|,�D�z�M�~4Hm{�?�TK��q���w*�pb5�A �F�#\���6pՎ+5iK� ����$�iP��?LE��"he="?
�
T�,��-�{�j��ι�_�&��R����T�!��5�J�h`����mDjYe4��s5�sT;I�\�jcf0���
�9��:"I���Ωt�I�z>^H��Fͻ���Jp=6p3�o?�<��$U��[q��u��l{`���j
XSTۣ���@}IZ�b���e����xR'`.���#����^lSc����Ļ���5�m���U4�X��!�}5n���͞=��X�/�T'�[q��~(�U���=�B������#t����a�;�J�8K�J2��B��E
�k�w��o\6��S��9K��ap\����j������Q��	�_��7�i��)��]�1!�3����S���-7b9U@�G�}f�x������̸�6�Z�ov-f����i���a��tv&*��H��c��@��l�x�ud��r�x�W�1�;�B��QV��~$������Vʓ��0��'�CɇAؖ�c���g�,/�
�~f���:N�N/�1�8?�Y�	{%;����{oi_�]}�uT����.��W�rur-�tm?Пl3��3;����\�ɹ;�������O�c
 	�S�sA4��Ӑ�1��=���8?̛�u��.>g��?!���a����N���EV�F�i��{����Y��ouB@0�(��;��]���x�A�9=�X�`�]��,*��u^5��6Į��+��ib](�m�fP3ְ�S_��a]н�z[�I�﵅���qj��>N#�($��*�=���2�X�}v{�hmp�}�៲g汑g�iX_D A-�����r�$���gt�M����~����v-�<ό�Z�אP�|����3�����f�\�u�~}�كH��_*�bΝ�f�̭CDA��'�Č,��Go��d��c;́�R���G�s��u���w؈l_2��K�U����O�}���]
��F��5�z#�9g�x~sɋ�X�54,1�s��t�	Ym�ɵ|�����p.�l�ͯ!�Gu"��ä�1�cb�����Ǆ����7���3��N\�[+e$�\Q]�p'���XE�q]�^���I���|q�?�A!�E��#I���ח�X{О��e�����>牔��(^i�J�������C�T�峼JgxE�8H[- �$�F{�3(�oԋ��C�03��p$���W������ƹ���H��͢�4�b>+���^��9���5:�����}�����-�&*[���a�w ;�Q�ҩ^8�`���I'AuO�����ŝ����l�dOB�Egc���=����ҩ�z�F� Q������h��W��\*�'=�����y�.SWv7y�l>gD�˫�b��g	����㑍ڧ�����	xb�~w�t(��A�L��