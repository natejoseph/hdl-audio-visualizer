��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O���=e�h	��f4O��x�jrs\���ô���)7��jꢤ��b�h忿��Q��Q�s]��Øpءms��u$��{�pS����� ��J�|էS�1�M�n��r�ZD��ˑ�U�_��J��jg���Nl�G�OqV�5��(n�����5�U��:X�)aZ�|����R(��n��n��i}I� ��R-~�lE�0y@������<��a���ycS��vr��j8�$���b#�Y4k2����Ch�/@���Arn鳂`#�n{���ed���Z�e��}�Jؤ���+6A �T�>o�g t���a"\��0�@��@��!�<Ӣ������^-k�JL�Aܟ���������!�i۬�>�܆Vf��Jx2��Xp��2����<YaƠ3��D�[������^j�Q��`	V�)`ٶ0��ԸѲ�
�t�I
� (D��\���W�4���1إJ\f��Ȓ��[����?b��@Zp;i�� � ��/p���4W���&�3jK��lꖩ��n�iv���Ɲ�;�� �����΍b��{�=\ʘn���e�VKIP={D�-?\n�����Pʇ��ө��c,�2�7���8 ��O���
o6�˖�LW����m�*
Ґ��DL�"Mf�N���|��4��v�Ɯ����-Z
�-Ҳ��
�(��`�oR��PGI^�~F��}f<Y6�o�`~Bo�U��C�S�W��F���{^$,ӗ��o�T������j$A�wDZ��;��@��:�x'|yh�Ä�m��Nd�·����)mR�U.x�[2�R�{���sm� 2�p#S�Rrܶ(�Y�Ғ�N�ZgY�o�oE#��?���� ��9������+�}�F������}�i'm��[Z����d~�"��[���
ǫ*�:Q�����)��;s�ȹ�'b1t�b3�-ܱD'�+�Hm�LV'b�֢��z�hU���������t!:	�i������$ɨn�;������D�mB\�o�%Շ���Q*p-B6G���Ձ����b5^+��}x�b�Y��Pi��h��%�m~�:�¾%D8�͸�k�q�x"8$�j.w�	�̇�sw��O�����ZL)f�w,�����m�:�F咢�s�,?m�����f�t�Aa�qB� D�����/X�l�ݖ�8!��{��ch?�"Ԭ�Q���U�!T�Q �F�7+/cFc���F:
�ݹ�:v���`���e�YYT\pT^۪ֆ￸��(��{���ɴ���"eZ,tcMC�pd|9��#.X��I�C[���+��E����a\����X�J�X偨yD;]B^��r~��B��7Qm���"��\mL�����g�5Ku��&�]\<�{�n��C�Zy�;���}�1�,ؠM0���0w��t��cDG�<T�{8
�%�����P�YJ��E{���;���~��bbsÚ~
�����V�cI��(}��P]H�J��L��	Ckұ�f��*�aQ��8��@6Gs�b�ѱ���#_�U�9Qs�j���v�EW�%o"6��f6�J;�I��n�G�3�^����gZp��
�\�q.@ٓ��Y[��U�U�T��Q�O5�[�MH`�N��"���`8�!�d����GE� �ܪ��p�ϟ��Z�4��)�'�;6��}�fY�S)p`�r���ft5�/�t���� |�b���vOԃ�ڝ�Ԓ
��f�x@Ŝ��ȤC�9�w�o�y]P��u��Εcͣ���7�ƀ�h�������	� q	������²w��%��������>��i�g%}��\V�J8*���i�2��!�� ��|zBUC\߻DT�"�N���@��c ��6���H��y�2�������V�QPF<ؕ�p�\�2x�)*7��s�?ޜ�%}f:�){=~8�����.��AV&��/\%hDI�7��!#���G�J\+�\b�ڲ'/-�jy��m��=�����g��Q��g�}w���o���C0ttQ�1� �Z_���WY+̼gJ�:ML�^1b�#n��l��v���g>A��)U�����rS�<_�}��ܖ�Y��i9�yg҄�ʂ��{��j�v���Wbq	���W^��ҋ�ᕾ$�5���qNt�l���	��e0���l��"!0!r�WqX�Z��S�?SN�J)r�e;K���lȢ���)�]2��I���R�kF����'�`B���� Z�T�c��K���Y��ʋa_ÎK�_{y&��z�t{�I�'� �:��f��7Q�C@�]1B�'�Z 3�4��⋁r+K�`FZz�{nJv��X�n]�]Z��q�{��@ޙ���V�R������8���9R|��Hז��i���-����Xe�8��WP��Nt_���Tl����{\[�.��a#����pw�A�gd�BYB溠���َ�]���c$½0�|e��<��^z��^�ʀ4��� �>�~�gn�I�'�i;����(�.3�s�~�f�콛���2�ߓ�;K��#���Hȏ5�U铁\cj'a�\je���2�U�^=jY pgG�k $��#AW�l��O�
���`d��J�쇇�Tn�xщ�?�Q~�y�3byFT��0*��˞!�4��T��tfc2<�e��(�7"?��A�q�_�]�?EU��+�{$�k�Ud;6��<�UO���?�X��w�i�(�I����Ü��q�(�a��oD�0�s�;.��X�eH?��S=�����0E+F�6�x?�ߌoq����S�%�i9W�g���V��2��6N�m ����ƎO �]���!�7�[�r5ծ؊�-�V�������Ð��!s �,���B ����98'̴�����`܂���w]��˴.�Cͩ"�K&���1�� �u}��[��]��)m�<Q:|9���Y��"��>7��:�=,F*� ��T�hJKO��nQ_D>��\�=�6x��V�Dy\��B�PZ�g�����盜��̋=̈́���Si+��dq�^ayV ���fG�_|'/���cS��n�]
�(c ���hO�z�Id-pg�J9�N|K�]p�A[-Dԕ�I,�ۚ�h���7u��~N���N�	��>�M��Q8.	��PK�Ѕ#�*��61�7ջ�!X�ϣE�"��y�8�^��Jq�3u ��{�s�{ 5("�#�
���m\�h���h��� �[wܥk8��<�n���CoN~y�>/��sQS��]5^3r�Y��vk�&<7�j�"�-�[eƤIBU�� (����"�����o�1��J�5��+aM��NX�9�	T��o�Yv�t������P+�ÞmJ�ܐu!u��afM�D�Q��}��m��r�Y�+�A�G����]�M��+��(G�A���"���w!Ѩ���$���T���q9c�W�a`�:JV3� ����c^�l��,������g3�h4����Y�ч��'� ���y���?Y�R\��+�em�Ƿp+�E;�W����JJ	�C�����G����ou���pv�Ȱuy8�BjM;15�l!&��1%��7&N��d]0��QW��$���S��E�C,dvGj^ޒ���:o=���>:�ǻ����FX`�r�u������BJ�6���K�Ai���<��Aʚg���W#��Nr�����f)��|X�|�fe���z)�%z�6��x؍[zҮ�vx�~5�'�ɞ�����tE���
2UF�^��O����ۇÇξ#r�6MccX��^$�BA���m7H�JW��q��D��������+#�I��4��pYB�Q��R}p�ՄSɎ� �Ք%,�²֧g^d�30�\��v6l��7��X�N��*#~�Y�'��?6Ø2ב�%W�l�w�L%��}�@s}` G�`z@W����<�~\|͢}�෎{]�OD�hgM��@�;f���ho�7H9@�iT؍R�����{���ࡽ���;���z���:#�deٝ�ӷ��������b�Is�e�[��g�ԃ܍�f���':�Z�t����7�Yَ���O��J�y�j�>�<�DV~U�C�Ԡ/����$�y��H��:�/y͋��&���&H;�*��{�r����eS��Ac�A�$5��: ;���
�Y1���r�C/!je�R���7����C�W\�<(�lT�#��� �'�C�ꥱ��)�)k���������x�7%b�>�֍Sne�S�k���X��(�l1�w�I���5}U_�.>��q��Ȉ�[�Q�2�MM���w�.�x�-��a 
���M�︞��gC�G]h�J%<��QB3n��Z��j�ucCH�ⅽ�<>���ѯ�^�7v�LG�dhN�Dg����V�g%`��TnzfH2Ûe.؍o7�9u�����'�A�4>��	=n %�U�0��o��+���Ъ��P�	vD�1�L"š13�J0J���u��fr�����].�E��"��tǘ�#�����o̾�S���d�S>}�����v{_�k�V�a�m�o�ޫCY�?U9QH����)dJ3lb����Ǒ)��ra0���@%(�(�^h�~�^@��se�q"����!��C�'�"��wq�2��>ic�E)�{Cm7��vTY�v!	��|l��dC�'�����^k'�	s���p��������gϓZ��ͽ�B�m،�h�;���6�꾽�}����4]��YY�W߲f�RF��F5���/��?�B��߻���S���kV���k�@
,��80����׻��OJ��9uu�Kͼ�`�ȃ�,��=�T�X��-L�U$M󉶐�&V����^,q�:B"?`�g��%� �)� HX�fU�C,U������W��޵;͚�?��n��p�6�2����s���/�qcgԁ�bź][�
�Q�hC�x���rP����.�b���>r&��E�z^X�yT��{_��Wa�G|\?L��S�]�0�u����#�HŲCz)S�CY�����`��F/<�L�"���Y�����w���zH��#�dP������wO@rd�~�@��>�h�|�Zqs�w�����J�+q�Γ\�(�1�9�C���O8n?��d�.�3X���o �zn�������SrЯ�R�9�Q�~f�|�uIl��'�ɢ�p+d�W�M]�2�M��d�>0��:|�:Y|-|�>>J=?N��VZ	�z>���z�l�5a��a�QB�"��K��v�䤻��)7�L�:�Vfy���Y� r"R��.�ȵ���r97[lc��K�h������6=t���j�S�I�丈���7'�X|�k�wqNၜ��.��)p_N���Z5��|N�1[P�Z:~���]��،�y^�!����V��������&/��L�14g��mrٍ7��t�����8��h�f��3��x�Ҧ�=���zx�!ė"E��}
�QpT���ƙ��hteZ�/9܎J�6ʤ������c�A-���դ���s�7$!+����R��^#�M/F�����e���j��%�����>y��oBǟ��j��}�]}ѕ�s�/	2c�����%�(?a�'q�����^EBr�����������<,l��vb�F,�����ش���b�Hq��f3�?IH"E�e��7���Lo�a� �5�OxSVW�	�6��PX�r3�J�1��Xc��(]��9p�����~1o����g
��a�k�������n�E=�:r!e��*	l>H�፷E|_��<2{��ߖ8���b�Jt{9D�翣(��W|9�{&��>:�d?R���/�Yza1�It�7�Ec�5� 	k1�7fg�㼑�C�T98ݍ�_���vtH������LQ�Y�=x�{,�|P��;#��X*d�L���0[��P�0/�`N�ű��I��J�.�B���w����L`��(��^X��k�L���ډ���U6<�D�8�k7���e����%t���<� &�o�9-%�0V��bWh�ӌ���+|ʯ�Z�Za�R,�� B
p��OKS���^ ѝW�4����<��
��{-1��[p�\�p�o�ob���2
t����5?ׂ��I�+g�&�
\ϸk��|�b���`&����?���	C��儌�����A_������Ս�����n9U���;�d�����pG|,#N��6�t.���]c��0{�-:'�?`��!���iG�Q����f	��	�nZ���rhG\!k?�dN~r�k��z�^k�9�����T�Y�!G9�Y�\��:�,�[������'�C�@q��G"�c�;��D���˓�E���"����y�9��P�,��j����4���wW�h� �]�Om����RT��<��SIn7��v��0H��`��ȯk���z4c`n%7��5^wr}U3_xM@0n1��}���]PųQ߱�����F���ȥ��S(S#�A�F2qs��D�[��9a�N!�UA �e"Xh�+"���A��+�$�1�_%gȚC�	�pK3�bt!i	��I�+�F��?�Z���"�%�B�[g���C�&-%�-r^~i�W*q�;�����~��-ŵ�*5�J��VJN4ֳ!��((�(<vlH(��C�>�;Z�h�EgP�P�g��ǔ�7`�ã$�M�!\��x�VAK\>�>�Z#�܀^N�eõ��2�;��H�����q�ގ�u�N@Nד�jf8�}�� �L�@����]�C-%���9YC,_�cqK#9.I��x��[qg[��#C���:�X<���c1*	� ��������5W#U�Y�~��6�Sm�(�][�G�e�*��B̐e	��˪��dĆ]9 ��;r�^�����`�������ڽŘ�*��?ҕM/C�@eG�6,�}��x�ioQ� �v�ݝ1��DD��?պ��_�*V�/.��eK�c�<�v�9�u��r=�d�=�ϣN+c�#>���n/N�+�'#1���=�Xi��D?:67�f��_FK�&���@���**�"`�OQOov;R^�9�D��x2� GV��i��&WW@�:Wc4�B�a<�4X�;&�C&��/�=��q���5
{yn�)~���N���Tx��{��(����KR�g��vJ)�J:�xApy'&L�k�?�l�(~.�da����|�h�M��u�~܂�&��j�o~X}5�TgvLµ�����'нa��DYϏ���� +�B�p���1��sm�<흾z�j<�D�|�ꈝ��_���kuo�6ه?���>�d� ��ςp�*��w諭ۄ�-�S���0
΃�2����}D�B�(��r:N�p��uS���Di��|L�sd�E�3�̻��,5���nsl#��S[�ގ39����2�1�����B����U&���o朄��읱�`���������q�,X�!vE��m0�\�o�����N��̩�r� ��p;%�b�&���^����(�ʢS(�RE���}�h~��֎8�c�v�i1��@�6��nd�*l�X^d;)`t%��3EL����U,�z�4{ֽ�B��У˶����8�w��1,F����Sn�"�X��q��ƃ��Á���_��K
YCp�t�`���C�X�����x�})��λ��28�W EJޡi9�O��p]�7�u���d�]�g4H�+�Y�
���z>�Z��g���k.c�ʕ�0��S
s���`1����.�, �нN��ҙ��Q߯3x-���Ļ[*�̰J!��D��eR���l%�	�C҉H@)�����;k�,�d��2���	h�S�������Z�Q�Dߣ!|RnL�ǉ��ۯQ�E��`QK�`���P�>�zF�X� �{�G�Xzq>��(Eolǉ�T�Z�ȮȋЙ����:8�QkH1�=�t�R*����l;���JZ�tN�S��ⓓ��"��W&ڜ���'�|�^���G7b�� �F�^�[I����z���h /6�[�v �{��%�gh�xqx��Ȃ(ov!�җ��������НΔ�d���ǎH��Y5ޣ6h��7��9Zf��'v	�+�^B��0	�Sp�� �&�k�p]Yha��G��q�)���9�����~k�]Q��<�3�.TgR�sa�SD7)�/�ь���n��q��|���,�Jz\�,�?���O��M'��ֻ`�$^��7�GR@.�1h_�Y,�����C�(�Y@VtBߊ*E��~��Z���1��1id��f�:"&6��~+v�T�Gb`n�����;Ja����_`�p���/��vo����Rc��$����l�M?�߮o����V"�܃-�n�!q�ap�<)8����\�Mv,)��.x״�Bq�����Q�p'���沨=MU��<M��$��SpW!�n�����]Z�1B��'���o~c�n&<�@ ~��܋�P��N����3����+�����Yn���'jS1�2������~]Q���ZK��XEg��}�)���V\����|�l������ī}d� L�� �0���K-���'Kd[���u��Z���*��}�`A+;�Y-���y"�_p���ϡ��|�UyE�Ըq�W�g���o����I	�y4y27Ex/�w)T�Ӊ9s<�H�k)c�2�����j[<6el>S�,�]�nm;TXnpC¢����Gs?k��� ��	G��Y���d��
(-"y:r�CL<�&��
7lc��<(!��(u� d��V�]�H ��u���XJ�%T��S�1�)��ve��*��F֛�ϨĿ�m�Ы'��=|D��V-��,XQ�o���:ɏ/�;�(fO�0L�BW_��V�A��� mz��*T'U�0a�3�s��J��4*}�3��E�r۳�4��J�����4F|�J��	�D_�fww9���$tP��U�k�s��N���Q��z)�킥6s'�wu-t �m�-ž���k��s�@p�Wț�Ѓ��4�feԒC��]�2��fU�8�Fي}�Ս�9���5'�a�FM�f(+!�=�����\�{- �|jq~�XJ8N��&�>a�,��\M�*JH,5|[�ǅ'lKV�!�@,��� ,#��/b~uyhs��<�o޶�;5 �$V���6�MTX��Md�ƅ<�6��m��O+��� O�\���2׈%�P�q�}}D��50����?�XϮ�|F篱�/�a{���`���Kh3�4?�xG6�!�l��F���
(]R��ʉ[O��3�[R]H�م�����KR�N��ax:FSN/�zT�5�C�G��mDǈ��n�t|�*>nL�/l�i#�I@<bL�f�`�]=�y�I��+'�\�L+��q%�9�ES�9�T�����V�^��㪸芵I��pI�*�5׋@������J4pb�A�b@ὣ��t�A��x�߃l��U�N��^� ��۹��,���)�U���o�>��#���B^67�0�e�c=�xKh�v��L�yK¼Ŕ�߾�����Ma�V�,^�)�#U�ݺ�	P�bq��j����G
����>���[�b�L��
���*�g=��S�^2�^��=U��WBm����$��u �F������ �͐%1=D�!����>K���|q̀P��]V6�����]�����Ro����h��qł~�F�\Ga�8��1��o�~^�B�O��k�t��Gc��,?Lџn,&�� �V.���]Y�Q���.����F_�'A�p��r@��z�V���r��I�s3�ĨЗ�d��?�8ܹb����T~u���|;Lb���d�#�V0����h�ҧ�>,�ę���~³�::2���B�%���̲���p�ؾ���Ȭ!}���U��hƾA#��@
	GO�:�ln�ΙU�xDj|FM����&ͷ'	$�ċ�}"��d2��{��k�:����ɗ�R*p�h1g
w�oi��}|����-R����}Dx�����ocjֽ�9��D�V�9��b�$75z�]����%&\�K_��ϝ�-�8����u��K6���&�ߛ�tO\#�`Qa�ǃhy"�X��6��ǣh���f�#�gҦ*����s�DR����Z���U�s��8$o���Q���>����SNU�]�9w���:�+]��jj���D�韘����=�}A΢�_g���W��k?��m����}솖R����I4u�]'��X<mϼ8�J4�k~�o�T����e��?�@_9t��G�q�Ӫ�C�p����=�7D��Y�5o�����k��>�7�����k\I:�$V@���JgN��݂@����fFS���@��$�z�0#Ħ)5e?%?`����&�ţrP�OV�d�y�3%�MĴ��Zh�d����{� p��HFư� �&���v��z_��}A�u��k���$�^S�f]��0f��e	��t4_�����N8Jo�9�N��=L�ru5'�r�'�}�7��f�Pp��ٷƾ�쒰�d�������+�w�J4�#�,	Nޔ��Gn�`&��N���MP������dpqY�gjN�G��ʮ�GK��8m�D0ّ�����q��9�o͆ݩ4HyW+���+YI��#��h��QN�NVl0ҴA�*u��y�]�f�$i�ab�Й��P�2S����%H������Cіi|*�v5�6$W����x�=DgzF�go·��گ@R�Y�PY,rQ!�P�P�M�����y�L��@"^ݤih��qC^h�����g�gY�23�ѓ냻 $J���ʐ�XOo�k�K�0���J�S���V�{�Ι�2���^�IY���oD.��O�Ng��;�艗[�)�Թd�͆!t�l�=Å��$�_�	U�1O?��C��]�h��;���%(��5�[mĭY%�j�w۫�
���X���$�
L�ɫp7L�Ih}�߉���-��\p<^[��������[���iҺq:3^��'�}���}�t5�`����0�k�nr��h"q@@rf�7l����M�l����I�\w���b8�'HB�~.�	��b�&�Y�/���[z7w�X��ee&��I�"m �nnzG�k����v4#��4S�m/$/$�߈��h6}@�#��-�R�����5�����O�c�5b|�Ù'�U�e�F��!��2n��6�tDG{�N�tq�9$�ޘy��G����MK���G�Mɀ�#N�>���ؓĞF�r���qG�E����nv�V��AEM+c�N��mB��{ j��^`�Т�-��ɖп��������Jkr>?0��p��.�,���%S�����C���կ�Y(
������ᗔP����M��VႴ��@uDCʚ8oo��f��fm�6F�	��vu)38�/���dM���@m+<���r� R�?Z���*	RE��4�F�>ʢ�s4w���H�ߪ�u�\����zd�66��̈y�:��C1�v�G]�= h���͑�*"����*f���?jC�)>�r�@�����+��S'��F�se��J�Aa{"�B1��n��U�gW�Z�7�s�X� X�L�������Y4�������}-�$�x�p�@b��Na�6�%fK�jVZc}�W�g<�a�7Zx�z�C��Ђ'��Z#��9]��aW#�����<=�3�����3a(��p7�qq���S �Q� ���qω>�
�u�*���皈��|��op�Ћ�G!s�e�g� rCI犑%�F5�|B���&��_��̫a��w���$ś9P����C��y�����DI��nj�g
�z��]��|��H)��;���r��%^s��_����-�s�]���e)�>�I�bT�,&�k��/�g{����0l�S��q7�-32=��/?�ӕ��I��ۜ�	K:�]e������X�Q�ˀR��.�$��]J3(,���|����DS��B����ͫ{s��M6��(Z�r��{��<�Zm�[�R����OR��R{K��0"o)��?݇���3�N�	�,�U!�8���{�!���7C�R!+����Ԗ����>t̛��<�џYΟ�5�<���xp�UHb�q2�T�Y�pWĹ=��Y��Vt6n�4��S^�k��%�:�,�/��.���#�`�EP@9Ś�������*�B��A���n�N���뱏����Z��#0�T.�r��G���������B�*R@���`p�{�5��ɲ�������� z����e��@v��0�r�W@�π#�W\c:׻�T	W�/a���u"�d���{w�����P�>�]��펄s-[���&F-_�
Q�N��K������&�����!Ur7��h�_�	����،�wժ��Z%�G�b�ӫ��P��r�]�L\<rͱεn1��,V� ��,��,�e�z
`ʃb����oڊBSj�mn� �ጋ��;�X�c�L�9�uM���_�o��܈�pD8#�v�Ic��q������3�#X����~{	l���p2��� &�(�
<,��aOA�>���yh�0��9y=l�	��.���{h�=>f$Eן5��o�����H�;p/q�o��2{�/���>�>�d���!?e�;���}w*�P��&�95#v˫�Q��c���/w�7��aKl�<���|����.�n�mObF��_M+a���3e��1���"��;E����Ѯ#��>���Ne��1}^|1!6s!
�5��z3@%�.���Wsn� ::��p<Q�~��TYA���l�̡���C��� �Qط$��P�! ����#���f̳,��r��-�%ש*��g?@K��9�`�W̏�Ы�\HS��2-+��ɟ��sV.�`%#::�F=l�T���'g�gf<9𚷱<�Sط=Ŏ�4]��{ K�\S9��]�<O)��|����g[�eE��pĆZ��G-�6*�{� ��
�ޑ����-��Ul
�.���Cf E����_�K�M7aCo���g1t1���Ԛ~����ݚ,�c�}ɰ���������U�9Ո�?�y�p2���ѱ��FGr��0֒���L��tL21�$ZZ�@F����I\D�j��6[�46��]�zs+QΒ�S`��<U�N�M;��u��d\_R�.?_���̀��$@V�L��G���:Њ��c�&��M���\QJ$�&�W\�f�n4�A4�!��	NQ� ܣ`Ǆ-��-�(Z�7TX�N�.K�p�R˧�S2�jX�9Z/�*!z!x���q���p����s��?�� Y�v_�����ϒ��%4d8̶�c�t���|��G�6��*�����4�8~�qD z���z.���u�\τ#����c�bX/��r�o��?Ϥ��
~xb5�uZ	T�.�>*��B�Y$�/������m�O���8��$lY�x�fG0��� f���Y���1[�`=�fX�N_;p+���~��G��,zM�<rP�r���6�N�xUc6��z��`+�/=�_,b����:o�O�l�Vk@D����Y{�umc����fn=��x�`�$C�C^�6t�˧t"xvI��B���D%��f�X����'ȣ��������@
5l�dl���O~���68�����5ke�Y�8�d�oUS ��gy<����[�]��N�L<��S>R��{�$����|[���)<�6���S����ѐC��	�
C'�oy9ju�-g
v���u<�6+*&<:��`��5��s`��f+j&*�߲���S�c3�p��a�!E,�u�mkve	��,=�Q��2���� ���?�7.3#�nW�z�5/��3�MP�7rM�?Co����&@^t0w��ڏ�w�fo̲���E�{�R�#��_����K�`���]�H�.9r�mZ���W�@��W}芘q;�D~�n�����+�B���<� A��:�z==37�@1�x�RH�6 �]�oP_�ܡ9�-��ѯ�}�5�e��Sz	��ê� ����g�����c�f�86?]��%BP����E���m�(��3���>��I	�������HL�/`�+��_n@���-��K�Μ���t����A(
�܌6JJ�77�o1�C��aD(�8�	�-�E!�Y��^-TA�zM���^���תN��eAZ��+�w#}Li�F%/%�O��U�f��J���[� KmA$� ��?����xO{j~&�� �ړ�i�I,R����o6��`2�N��ms"6k�iC��˒���w���&���zS:q�i%�N��fa_]�`4k���E!��+i�o�|ByhMH��ϕ�B�y�n�g�^����q�����K�Y�RX�h��s�/\s#x�	�
N�0(��L�K�1�v@ʨjk>���7aR���oh�a
C�c�*<�:6m�G�|x\M�%O�mɰ\}-h��#7G���
�]�߁.0��KH��hX,n����{&&{v��9R�OAi�����e��� EØ=h,F&�M%�3!~M|����^~�ɓ�����b�Jw�^6�c��t�4=͛�oщ�wuv�E�+�;5B�_�7�b+�F$c�BJ���Z�;I�d��92�� ���)'R�>nw������0p��X�Av ��?_/ns@W˔yӇZ�k�/^�����3}�0�_ì�QV��Q�wo=��U�T~�����E�F�ǭ2sr�W��N��]<� .F|�~��4;A�dZT�`}��'�Y�X�/;ry�C酫|�w�A>�B��>l�[���]lCr>�=?g�bp�m��Q0lۀ Q݉W"��a ��>���R���9���_����s܋�/��&�;,�j�Jh��udA8�6����l�g�5%�=|v�eSh����6��t?Y�dI2�r����=h�֪o��K�-횡G���B��t����e��{�J��V`R	�t������k�=���e�&CT=�x�C8Κ�h���jZ�p=`������f�B�UG��n/t��B���x�z�Q��8�S\7�I�ڿ2�r�AYM;��gQ�x~� H� �@Z�j2K���%=�N�����}ćZĶ,�
�A�<��\��ÆL� �7>��d�3[�����q-8�-��R<�y��O�Þ��*����O���{Pz���;m�R*T4K�@��̪�%���z��۳�?�b�N�E¹�T�g�e^��V�<�E	��ئn1�c����	ġ��\�-���@lP��%�E^��I&FP��=�5tf�mm��&�}�ݮW��d��|~V���E>�>·ܽձ�Q(��"/�^�Fa�w'YnC��=��r��Ɲ&�KGȫI���LjzJ�I�Yw�>�m��|��\ɤ(��'�O�E��q΀������@MK����f���� g��_ו�3�;8/����;�����v���Jf�o�n��K��<>��;�	�x(��j!����I���@^%��l��蒓�=�)�I�q�L��`�A�~�H�c��v�3<�V�y�1���K���'��o�eU�<kqv�#�[&���u�UZ���Q�D�M�ٳ���g��dM�ގ�f�IdpT?/ ݫ.c��m<�KUi0�!L�nTE�Q�oTi��y�ub�YCyU�~�3ؾ�����249�j
�TB6(J{S	�˶��槐RH-��$���)rbɘ��(!7N�{O��\��D&9b�ο���$T^�U�㹛&����c�
�;!=Z��͞�s�`q5 -�s�v��k�n�?�X)���z낣Y<�y�.١^<ϊ���j�bOdɓnL�@.~�JS����[fM���|�t+z�<�G�:�-��;�3K���R��&��훐@1̹�D�����K��rp�'�����c���̯�����e`UKWrJ���K�pQ�uG�h��a�DG��ġ1Ķ�-�b,��ⷮJ�%����J�jgώ�����LZ��:���QD����E�������n5����A���y3���G��c����zN�؄?{�^�px���jdb^������G�A����♢�M��4�*�R/x��Ϫe��4��Q΍U0Kb�S󡈩���A�f��������,��i�ĵ��.G)�w���ʚ�[����PG��^u��z����|Z��ls�D�m��(��<w;w."��R����p@:ݝ[��sx��Uv��z��0J_��	Y�~=/m���ĵ9���qƁ@�s��)���P4��w4]�, ֹ0�f��,��Н>Et6$}2ј����tbz�eWN�	͆Y2C.��e��?V�j��B4�؄Ig�l�����,�8�Y���\
]�3;���zM�ۮ�����fE���6X�"Į���r��"q1H�ӥKP��jwc�- ��Ȝl� L��y�O�{�q�oM��{���W�J}U��C�!*<��6�CS�Ǭ�H��۹N� K����|����BK��G�v������;����z��|iH��m�М#\h0�(_O�b�G���h�d W��%�r\D�ă���c��L͓���4Ptm�2A�����窫%o�h�v�ݘ��iK
�F��_������#"jl3�-&�SG�v �wNI��*��(S��;�oR6��23M�?8ބ�q��t0�"[�5Ģ]�� �ŏݩGb�\{��D^�����H��~S�,�.+b�Eg�8�Ƒ�F[X�^����T�.D64�{�����w�z�h�͐2ǌ,�+6v6�y5�Z�ǉ"C�ޙ�; q�8����Q�$�)p�`x�h�"����a���-�C5��YQl�~�q�_�����6�~G)1�XA����V�TQ�M���k��;��
��w�P�S���lm;1��Tr��:� Zo[�>���%���I׫8Poyɖ<��&���F�efY��(NR�=[��mI�|6�gb�X��S]�&�p
�F9����i�����P�@�Z��3sGFd'���e��?!�9��8�A1��nҼ���ѷ��Ơ��Ap@ʓ��@��]��I,nu�Ǖs� ��!���z�N�����H�O�E�M�kp�|Vt��\}Up�Ya�L���_^F-w��k<���ڎ&������Dԅ�2��R�"�/>r�&�?7#M*��E�<��!�����Kβk�>�$�d�6c��<g��D�$�(YF�(an��*i��ȉ�h#��#��aPPYoƠ�W���6ݗݎ��}�~!UZ��8���Q�s�ʜ[H�	x�F�Ѕ�;�f��n�>ۯ���@5�[.	���Hp-c/���}��h�n���!ۉ����x���2���P� ɸ�����>CAieCL�~S�t3�{q����nR���=��f^z�j���(��=�)=R@�����Ÿ���̤+q��$���H�(�h#u{�� %��źHx'|.�˃C��D2&���������@�:�|�Z��.�wЧ�`Ulz1ί�j���U[�Ɯ)���7i4�T��s4�_!>tyB��h�?�Xw'�1G#!��2�9]��ʧgh�џ��ٹ#�P���3�c��<F�и,tc݋@\�ł�]��$��3�:su�i�Y�hC�I�F2P�ZѰ��Py�ƞϽ,.2Q�^��S��h,�H�Eu�ʀ���I�N��������ę�����;���V��s��A=ZTdM_5��4|�;���-�洔��uB�<X��(����+�[VO� 1Xֽz���o ͬ�*s��7� 7��x[J������,�PI4;��������J����˾`C�:`�!`��>&��d�v��ѹ����K��7�0�	��_���ͅ�e�I��Z��\t�����n�:��&́햸�BP�|[hx�
 ��??���LO|�h����/20��xUi|
mw=��R1�BB��.�>i��ڴS�n&0;���QN�7�G
�%���w�^{���=��j�����0̪�T��N��?;�����������E�$DЌ���A�i��-���I���IL"����4��j�|)wX��88j��G�[D���̾��#��\M��u��D���Z�j�"��=�껹c���<�Q�vf�y:0+�q��a=9e�o WV���\ىY̬rz�h����v*�c�F#�ֺ���\8i�bF"?T��9lO��o�+f@�I���O�lnfT�8�~`��.��3���&{!�c�u(|�g6���2�m�����%uV���� oK+�l�7�t������g����,�v��bu��Vm���LN�#�s*�;H���\z%�AEI�j��
�1"�v�"������{;��إ�Yn��F#V��y��)Ȟ�7��E��y飦.�m-��cQ��Ԟb�׻�Ō�ि���r#��>��lؓBf�"�@���I��O����X��qjϟk�@����$��`.��K88M��%uU��2����S�g�b	�=�� �.4B�0�:]-?p��Wd�	ea�3̗Xע�Z��&š�@d�2�X��/ i�/�7j�ON��kq�zk�,������g��E=���&,��n�4�B��JY🌪������A)��$L	kC'em�=��&�e��7~�#��+��C�B�T�}� TP�U-�o/C�d��,$�V�sH�Zq���� `#�v8�Ӣ�V�R� [�bY����dS�k��=���������X�6��Tn;�Ƌ���QqA����'V'�s��
�u���ɽ���G�3p#u1ޛ���� ��]7b�E;O�E��`2\x�۞�����3WP�w;�X�=�c ��w�3�6!Pߑ<�1A��Z^�'A"��Owr'����X�.��05s܋��$��G�ڈ)D�f�b��Gb�I<:H�$.�tF�i���~L����o��HBv�Z��,�3��c���II��y;��ۿ�j䐒���'�Ol�W������d64�nw�68���-���F�d����� ����s i����4$�ْ<u��߳׋B�I��*��H��r��K'���{a@χ�������W�b�8��,]+��4��Bm��r��%�@�ZX�"b@�I�F	���j?���f�T�?J?DL>(�ӛCs1�����������
(UK�9��j�J�V>�^=���|���9l���"���g�'��+�g��_�}�Q�+��B�M��{�IbN�ޒHT<h�B�O�uq�V=��BVV��K�Μ��w��|�˶_���t(�vZ;�n$7������sN���w����}`3�2(�@'�u�sڨ��U#}�N'�K�h$	�ͥ��K"n�����HZ������=f�4O�+_��Y�Y�լ�\�h=w���8�7,$���ɗ] �g5����^��F��)�������gm��q1&\�� �&m����S��G�W�%e��:E��1%���Y_�u1��q#u@�>���P������'�J�~e�Q�����"�b���D�`���B�V���)C+�����x���ne+���)�K�	n@E!����rV+J�f\�8B����h8���˅诓rC#HR�⸏��ٔ���{� �Ŧ{m�LE��c�o�q2�>H��ή���p���4]����*5R�2����/ح����)�I8����R:O[g�pS�#O?�����uC@@j<�t۩�[�o�����}���I���{�;��MR�+�iX�I�
Z������D�:Y>�=�q*r�����a�,��
�*��
��Q6�FfpLew>��	(���5��/g�#�Y),,O�U>�ǐ����ؐ��XMGD�>+ �C�r:�Q-�3��P�CJ���;Ǘ����:L��� ��Xv���d��y����P�,i5v�ڵ$Sl�3w;�?s ���[K<M7���M��=�%�e��=t�~A;Ѣ�b	/�$��qŋCqn�>�CfID�Ť�uGC,��n�lR��>,4���:���lR��&J��S��������OJ����Y��Y��q�M��і[f�~��3Iy-��C12���v��P%�f�Q�����R$r�"2���贌;i{\�h3	nG�׋��+,��t��n����~1rHX5d��pU��xg����o�r��P�ǔ'䞮2F� 8O�拉[��\�E��O�"{\']���@���W��:uI'��7.��u�p��]�	"���lBh��e���J�c�E<I6�mM��K�RH� ��T��7�o��\ݷS$*�y��A��݋�Ur�~�􄭝�߉�#�9��A9�
�si���!���#��*����˾R�p�2z����gT �G��C�X���4�,*��r��s*��CM���6f��пj���2IE�&��1�~�W��_���}����ì���2�K��UAߤ)b���S�VS��)~\g��"��̓F��*� T8o����,|R6��G:�`j�*C?C2�4rв�tzﴞ=�#�H��h1�$	�^<�+��H�Q�F �7*d�TOKԔ�Ʀq{���,���k����4m�jE;y�>͹�-���F����W_�H�v'!cS��~$s���g�Lڸ��h�s�=����R�(e6�3�wȣ�H)��E}ۻ$CV�[�e��a/�[Ki�f�Fk���*����s�|Y_qV1���A�����)w���ON�@V��G�!���A���cWm4pcz}�$�U�C���i+�t-~ �Kλ��S�5��� Ф�r�"�q1�>Z]D��֨�?�̱�o6x��ch�����vJ��P�K�#o��4��(>�"Z&�PLw����~�T�V[68MK��F�  Yp�� v�����)�^f�Bc�q���0��]8�6��(�W��a��]{�uI���}�'�g ����~j�2���%�1qç-��0y�
���N|�����%K �<<鎦�#�v1=����]�?���D��eU���5o�ă�|��>�2(��G��ܓ(z�����L	�i�j��Ĭ0������*f��~�F�Y���._��O7&I)
=7/[�+�Z	=.���4#c�jL=�?�@�ɧ�o:�!���1U&�z��K�b<�dț�*i�/�@�F�>ך}"/.%?���1�)YC��| �������U|�A��-�O?���?K��G$��[F�B�:�ɪ��:d]�lu�ꛟ�P�8���9��s3��O�d�JY�X��㋋�Ս�]���6��Z�̸R�_A��I�^�����si�T]eJo�|n������?�>��n�:1y`m�K�����6�����6�Tօ�[F�C9"��5@�����W]�̾HI��F�~�k��!f��o�hH�	ƕ����M�R�%�`���j�y�#�ޮ��!+�GPB̯z"��$������ʋq}Q:������V��6 ��X�vy�K����h�F�a~��sدl�Z��y���M�N	3ːG��D/�¸�MU������RmwtZ�ġ�_ ����:.E�P�'���ٺ�P߃�ߖ?%F*�UQOW�.�ƚkf8A��#gH'���k�*�
*�B�1���L@���o�l*��a���!54y��{��L�%G)�P��+F��*�$m#ŵ�U,$-Nk	��Mg�[X�֩�7�@ TC�d.6W����'̊"���~X��I�3f�{�_� ����l0�ߜ
��4��q	��x2��(+jӆ$�q�$� �L��!�TD��Uf�/G��N�ڿw����X��%�A�CFy �ɚa�H�/nJ�%�CJk ��(�Gz�2�f������x�G�q��S����dl=�t�$hi��hu��D�b��&�)�9��D���ن|�������+�3��ퟐ4��ԁ(N���C���@Ju��5���L��
`��:{!�k�������ǒ��o�����_��G'��\�[dyǰ"���n	�i�Ӧ9_��h�����D���@�5�|*�5��}I����u�qy1�=�l}($� �J2�4IU������)�^�Э>=�=5���E*2d�72�c�������U(������cKu��8O�<`�{3�e�Q��w�YvxCy�J���c���qsM"1S��@o��\��xސ�ֲz���9���2�4�0\:k��B�6�� ��#wc!�([�0pa>��)�!� �����ˈ��Y���}������_�Ҹf�^��D/�Q��u�:5f�ဣ�o�dJ>Ek��9� L��]|��b.��>�8m|�1 ��/%�j֨U�E�J����a��	Hw$�(��g;h��D��<��ȀLh/oW)"
���+}�#`��&�M{�����"!V�GL�4�7����I]�)�e���&����ַb,����<��қ�릟���瞀�B�{�[I���1'rZȉ��x��v�3��,��C��Y���v�@d����"��mf�X>A�7�F���Ú�jٟ��j���%����w��k��r�׍O;����2S	��Ec�61>1U�{�����MڅL��oG6.v���`���#
���B�:��c�Θ5��~����q<J=lN� }�(�b�� |�� *�0:[�ca�up���T�јY���1V��c���H�%9d���Ѽ^��R��
n�����s��Iג#� �r�^�`��}�'j ��]]-# \E�-w�j�v��s�.��#�4C	�U�����6�埃�M��H왭���U��E������P"?'���v{��4f�ʷ�2�o��]��F�B�� n�e��`���q�tB����Y�n�E_^�r����s@���(q&E�P9`���5:�r�v=���up���	���6vp�6P�W�$�L����m��tD���[;9קoy��d-�.����8��s�����.l�Hd �h�GG�RkB�E��pm���YY�9E[���E���* ֕ɽ`��T]��$il>l.���h�>
g�s"nܺ�Z�"xF1L�����i3���ϫ�?�n�a���O�x�Q�Y�v�2�8�����||L�y�q��� )#�w���@J�ef�ZlH*:�}q�X��}�}��q� ���\�&����
��alt���uM!\x+"}	�t�eJ����8ڞ�����i����U�g�|�t���b�c�}�6��+{_����~%@�#�F�7q�o���J⾻��	�����E�|��kFf�\{ز�g��U\q��zM�$�җ���g:�n Ս�Sl�0���!���� ��a�ܛ��Jl��-Gq	�ag~2���WT�b4-��В1����ޛ���>'W���>�y���`s�W8b��-	����o����@�)��E���"�ܾ�U�~��{��	=PWC�J��Z�ae
ʮ-ưq`�%�O����_*���di�Џ{n|�K��Dy�׏
����.��AT�Ź�T����7$�\�t�<2#�	밭��z5t�A95]�O����)_�#~���P��s��毳�dM�	&Ҵ�lf��o6a���?�1\���e�1P�x�~�Z\��BQ�=F֟�N� �V}�?e�4�+�:��D1Q���>j/��}����1��hώ��?B�0��,��j#H;�!F O�D��T}�Ĺ�;'�_�ς�/4��a�&vx����ş����_囪2R~���F��c��~!�����i�}���L���^�w�^�?):��S��(!S��q�Х��Z�i�M
��Ͼ�F�'�4��=|f�
� �l�LȜr�����
a(��|:�F8>Q�4~nf��#sRK�ĵ=�{wpK���w��&N�]t��ĺ���:s�����;�_W�3��7�|�� �^N�N͝a�/:d�elk6&�!fQB2њ^kU��v�7���'�m����p�.X�'����L/��zs�8��E���E�:���Ώǩ�LX��	�^��(�>�C:��r���]������:;�PMNz0�'�,p��"=8�47��m|�j��e�:�&$q��곤�;�}�������%v���$��Q��҅07A����e��� �D������렌�u�͠�S���y�)/��
�I����(����r =������H� U��7[BQ���=��A��{�T'y�y��c�?�b���cFq��F�,Ldl��D�6�Ef2-����d~w��r8N�N��Qy��� ��R�Z��M)+�z��t�E{��WhI~+/�j] ��R��B�R�f�����3�B�̿wV�L�*��G�L�����	�pFy�	�U~$�-M���2�!Qix$���D9�e*c2���,���f���ǀl�u0�N�����+�-�aX��0r�˽��Ěe[�<�y����~	H��	<5M�7�M X=:�]�b���*>
!T4L�;��@�T7-� �r�r����36~�?�W��,A�w�f�t	tj��e;�!3�$at�����#���m�^��_�+ƣ4�H�.L����ߐ��vc8����,iRA5�a�?`�Y&/��Zr��@�S~a)��M�X�Q��1m��.�׆IҞ� xp2����O��q�@�5��O�����<�h!���4r�����m��+Q9\z;�@�:��.�?��7jd\K�"�O����Å1�V��WRj"FVtI���Z����dU��Ĭ��	��]��d��W�o��z�o=��i�0�2%��\nʙXs�ơ���v������p�#U�u�Z�a0�[Td����Y³�i�/���}j8�����q��~٢�Χr ]*�w�f�	�)�>������L�Md�!�`J4}A���m	?��P�E���X�m � d&����U-�nң
w��(����*,���DX'o��H�����=����1�X�[~x�FC��IU�b��N�ܧ3�����nM8D�/����O���b� �+�j�E�},O߲�z2�y����¡��b��4�[@����?@���w���+�fI�щC<��(�w�2��
��e�T���C���aۢ�'�,��o%��y�Z� ��)ǩo��W�M&��R"B�q �T��vLI��Ŀ��M�u��
�+gh��
Q
7��n$�|�.Jm"	�B n�3J0��a�8<��
����F�)َ.�6P�Nq3��GkR[P�O���è&0~���׋�i���$�k����I��.��2z� X��O[���������C,��{	y4��|��9C� �ƯV�@&�Ԭ���/�#O1G�{Zب	��f0z��uݪ��Q�C��N=�)K�md�V=�a4�*8A�$K����4����e���mg�������Z�,����	�:� pyL) �(��~^���`�	х�0��DS��r�B,��4�pX�%%�_<� @~Ӭ}��W9��D���q4�ׁk���H���	4y���Xe�G��1F1����4��A�	��m��%P����Uj���w����aå�{�x�k�ۧB�Ae/r�2Z�`=��y?66
��Y
AoD�u���~����:�,�,�.���d���C�J �~���>�툘���ϛQ��{շ�L��HJ����J�g�p�/��:,�eꢀ
3�jaK��57~�_n|ïO�� ����Dcn���vΛ�njVQ����ǁ8��� x2�Oe1}�6?�1�Q
��c�W�@YK~2c9FP�];Ym�'*��[��EE�.]�pr��_?]S�nR������\��U9�oq��}^��P#�5��+�M��D0bw�ǚv���gÆ�#��\����ŭ�G�m�8.�}󍫫9�Cc��ճt�R�h�A���g������x�w�\(y�)�j��m�)��8��|gm ">L&��̊'��wg�U��g��Q' ke������28���c!�QƳ��X��"4״A�7��8�镧S�W���L&0u�?4�Ari+a8�ִ)��ޖ3�����e���c%�`�&&��ڳ�_�!���k��S6�ګ\%�5��<��ͳ��j���6�S}��>�����S����3�Јƌ"�b�D��Ƅ+�]�x�|�1��,V�O6'llz�/���6�J�B�	=�S`�R��1:�:�jB �--�Ǐ�;<y�y_�=��+K&�Cj#�s~_��������d�{��HoO�#��3��:�0������>xV���>|���܆�y��[��B^��:��������M��( W� ��<>-4�W)�62ͺILa���C�?δ�DG��=B�[��Z��$I(���cL�>}>��j�� t�4����Q=�5�q��@��8���X��Z��d��%1�(�&��1�E�X�a�
yʱu�0�k@ʷPj�)��r��xQ��"l(!�U�K�{�_���$��r�P���&:��I����<��^e1��fՙ�8���>�e���I�[]�j�0�M�L�U�s42�I�򁫻Y���_�	����\i����8Z_1�F�Ga�k ������$��JD�@��( �o	8��@�5�7ɈW�;��m�ݡ�t�bzKd��6�;�p�XW�`��	�h�=���S�����6��S���F��=Pc�ɯQ�_�06�h��r<,������n*���N�ϖM����PE|�Mn}�� H9:{,��8�%~��ڰ�֓Ciƃ�9��,#1���'vĴ�P��zj���a�Kr��]r��T̙��vSl�-V��Z��oT��U���3h�t�H{��Im�<�a�)i�g`��{�$eV|�a�pi*˾HQ2��:>^�q�,�;�17P��/@���s4��D�P]�؜������Fg��-/U܂��Q6�A˅�3TH�=d�Y���>	ɀ¹y��6�t;k�ofZO�L߆_�a>�!z�$�b��A�\���z#��+���˒KeR�}y�	X��C��&0a��Ɛ���$*/�^��H��{���Q�_�D_�5 �b�?�W�q�O�9E �.��*��%Z��u��*�k�t/�Y*Y 10�>����hL�$6��Z)J�R����:f�wc�����^M�uR���H3O���-f)��>d@f�5$Qc/Ⲍ� �2`#���7/mma��z���7�I��Z��,����w(���'=鞝���Xi$	��.�+B_�ʞtR�W]�fg&p𜠍��㼆�}�_
�`���5֧�����^����U�~��&��uX�fٍ{Hݑ��?�WB8�c����L&$�Y�8�^M��HZ�T�`7RC��3��c�<�#x��}b�1ʠP�r��JCyZPĬ�v��d
[�)/��y[ד�q%}K�E���qN�"�2���ҷ}]���o;k�Fny�v��/�.��z���5 h�		j��}��'qi�VtH�N��f>����>��8>�(G�����l70p#�Y���1!��a�m��ll��B���ܴp0pu:!)��h ���k��&�?	�Q}M�iR(��ŀh�+սR;�o�pg^N�����y����^�̅x��>V呭�O$#�~���$��c���Tx��J�E�y��t6�@��U�L�.����~�-9��4���ԙ�m��gԠX��>�T��Xz�n������8q�f_�k����}���,��9���:AqϋY��\���6@�b-N�G�o�j=y�R�^�+n]������o�<�\��SO��6��\�*�u�T]�D/\v��ㆂb��q�Y$qr�5H�I��4�_10���|b�\�!_-�gq�`�t��:\�KM��v�JV���]�9�;�#���aX��`� ��;"�*o�#?�9m�啴��~�E�˾�,o�?�I����c�A�A^n��:6J�v(��`H��<����J@v������L��Q��d�yf�O��=)դDhX�����qs?m�h5��~��>�;=Jm߬�'�9�h�G8�6w	7kt�����t�}�7�%��:��&��:;ς��q_>��E+�~ߑ ��-�Grى�hn(�ܖ��լF�0�Ax 7L�˄�5:���{�����M����N�ˬ,����cÏ�����N�0�Q]a��5���S�c��b���Ha�O�����"���N���1���uӉ�nO��j��>���Ļ��n�Do�;��0�W1X�I��z��.	� �8�C���%����Q8�T����\�Or�=����;Q�0����6c�`���(��[����\g�OA$�\��7)z����֞
���m.�H�k���c#\ۅ���u2��o�XR���@~�Oi	`겪�t��q�vA^����
��fY~��MRC SOңěޚS���N�}��R��?c?1(�Xo椤݀���./Მ��/��I�!1���3�T��>I�~�*.x��h���v8z~$8�U
	��U��_�T�"�v% �j�z�~6��/'�y���p�Y8!yZb��G�6t��|�AtO����'M^�,l�ӊ��h$!2&(i����Ig�m�t���9�ɗ�0nW�EI���(*������K����32GFpe�#�����?hF��n���D�J����-��X*~@��)��,�@mfsKa{N6�\�0�d`��sT���am��J #�����"K��AEQ��]��<��k�O���(oER�q=��/�D�C��ٝ�� =� ��R�q����4�ܛ�	X�
"پ��p^������7��h9�߽¡(�������"y%\k���˴?ʙ3�3���g����!y�G1�:���Pnj��+a��q�O6�1w@�G�;�������uѝ�M��P�ϼ���-|Y�^��f�S	S_�|ɮ%h����Ci*��b�K�ѫ�rhnkR��{��ce�G�F6�'ouuz	z��#�-���ٌfԦ3d�@@[�,��~7�J��9���D�>�d����� �}8Y;4lW�A���$5/	�O��;���{ݻ�%p����ekQ{�H��e@@����K�ja��W��^w�`	2֔���D�z��X:n�����玲=�y ty��#�
1�f3{_WnEV���0D�(#�*/�P�׶Y+'�n�����%�7�=�u���IJn�"bA�)�m�{D��*�bo����P�w�]l������ ��x��p��~�s���%���l���{��^qץ*�GRK?�&穼+ݮ�#��j1�V�\��@2�����  �+Ğ���6/��?�vt�˴����/�Q��~I���pp�M�K2�Y�A�|] ���Qm�j�#��E��E�k��G�jeF���j��!#9����� �%֍��*ڏ`������U��O�Zv��[����L�-�+��mvȫ�ƥV����V�\�ÿi����$�j�O^�tx����v�����?d�?�$D�v����*�2�e�L�%�����Cl�w[#� �ƲcУd6
e�E�Y8n(�T�rf��TI	t�E�P��i9�(����9�}t v̰=KO51�}�8�C����?Q�cBR��쥶R;�Dk����^�/���tcУ��gҿwXC�����5���� ���ݫZ'9��4E(����*l9a;bM'?��{f�PɂZ���	��ގb&;����pA�]-ǳ����`	ʥ�g��5���)&b v Va�G0�.#��<lR���=?���O�Y?ƹ��n�z�&�۟$�q�D@�M�׽MgYB���z�QQ��/"z-��l�������h0��t��	��j��S|V<S\'S!�� �U��Q}N*l�x������":@�U�tç�H-���}N�yE,,
�kH���Ã���`���b�2��tK.�3�Y7ړ�q���T�i����>�A��#��J;U*���F+��W�0�'����Y�ʼ#^%2Nw%��%S��L��T� �?�<�-����r���H���?{oo�؎`�J/�3�P@��G�+���/���UZ�Hv���4������;�ȩ�p��3�����u�n����@��F���&��O���:�,X��1$�<�%���M��NG �$e�Ip����T���P|G��L�$�`���2.��p8]"���|A��5\�?�N�а"9Za�F[���Y�� �5xt�11��l*����k]e1�x`�'�!f�t%jAs&ܲ�9�<s?�ȝրs��{D�-=�~
��וm��B�;lp9�ki :+�Vf�>���z(#�=�ћQ�ݻ���0M(�~��U!�Z=r^��onglQ(�� F�u�2��k��
N}Qo�+e� hYr>$����k��,d%.�9�/	�S{���O��}:��Uq���f�YsOCPæ���6$0q�	
Y�8��O@�Թ���P"������UA��+�����E]�?�Q��P�Ȏ *�IT�abJ8,��8�����&���-s6��ب�1>�ۜ~�>��k㽴�u�����Ѷ������f�g�F��X!��`y0$��+�۬�b-�
�677PvK�w�y���L�,�ο�{�b;��PP�m���]�9	;26Q�p�p+*WF6 ]|ɹ?�f��8�2���<9sm"�wP�|���v	�c,�8�Ϥ
fӌ���������՚rb�5@D��,�D��Up_|���`JCaTI=�`{V���0���Bn�O�T�?QiN���#ѐ*Vձ�շD1'�77%�"TW.�P���c�`�#Q>R��Pc���a�-�Q�	
�3-.���I�~�Bk�5GyJl��A2�,fd33�A���Ds`�p
�E�0�i�;��%O#�Dt���߿W�(�����.����GG
T��yPF�'��a�k �a��@�	�)��8�m�W�����f�8@�6�E�h�df��եu�o!�캫�߄���V
?������X�𤴩�nW����ck�Gaü��8O+G1�V��"���.�χ��9�p�Rz�)��3x}�)շ��1���	�sΰ�6
��E������ǭ������݅�z�1�K����2w�4�Y
�+:�R%Gp�9������<��=�Q��� �[�3��L���
�e��d�9c�h�x���ZL��6俱�
O��`>h�IM����m��	,+�: ���2C�Rq<8�/���~KjU�W��B����M��֙���Ѩ${������HA+Zpc�Z��$oʿ¿����A3���S~J���T)���<M�duG���[_>����AE>�Zߐ췺�Q�+1,��n��i�H�%P�Qrޟ���&ߏ6r�
�RriKJ
G��
uQ�˵��0�1ϣ�NW�	p27U�*�����LV���W�K�y�Yc>���ELx�y$|���PY*�)�۩ٛ��ɚ��`���0C�T���>^�}KJ&�=;�UF�<Ӟ�����.J`�2l��),cT|��<�1l{�,����]�#�+�*3�<���.$'W��6㷡	谸t��<�ε/&��׍��R��}/�>o���!� ����\ahvwD��!\X=:L�J/��Zx:㬍�����D����"����<,�X�K�)!��j�v�b�w��yч��zs�[��rb�$O�A�{ԯ��)���JTb_�+]�5	BؚX�ۖ\�#{�Fr���MCD�)�i��
�Q���e�$�)�楦�����>�=�L���/;�^�t�0��8�Vi+
`�7l£6��A]k$�q�Q�o#2E��	�mB--
ٴ��L�N6�^���N�S�fXe)^r֠~���F��g3���.-9s/+Җ��FkM%�PY@��k�+��EP�|�A=��� GQ�k	%72��|*1O5�[L'j*s���4:�����d��|�]F�5�1�����*'yvQ�o���{|/���9�>�?��v�M����l��)��E�]�'���q�e �'�Q%�����SC-<1$�10��w.9��#��1�Re��-�T]j*�y��C��zZҖ2Q8I��`r�%����#2��?p|:ր��k7�O�-���I���/�gYG�f۳ᾣ�K�p�Ā{k�U�B~=F%z���-xYZE+�b<�� ƣ����i=� ���C�a@���8K���|7�K��Eӏ��:lC�[;��0Q��߀���#�:�����̚���z���2�^�5q��Y�Q��Z��)�L~����E�;s����BK��ZU�~4�ס	��E��_���߫\3�&���R`H1�cYf����x��{����C�Y�3����;�h���24��Uo���lgd|��Ok*f7��=b���߾���A�U�u(�[E�4f}�.��WlqI� �n4�����Ƈ=�����"ճwef=�6�*�u[��'Rm"��m�414���)S!Qݓ5KM.Yd��-FU��{c��%�!L˾ˋc���Eßcڠ��g'��H7]1�@\y������,-��gw����!,�k!8 �p;�vo�̆�	x�s	�*)i�0 �4�W��F9,�!fi/^�18�ð�Is��#�Fn�Qa�;��>U;O�c�����e�-�d�� ��)��vҘ��p��[�`!
6w��1�f����㰊����*|K̲��e:�p��h�o	t���h�}��5��B�X̃�1���쾬F��Gz0�T��K�>�ݝ�zh�ʻ>J��W�;s.�&�>��W6xlZ�Ъi�	p<�ۈ#M T�i��b'̝�¥H����PF)y�r�CZO޻�ߚ��0�0
7$C	7[QO"���)��G�>�BB��E��B��0c}��Re�1�Q���4-�A�5_���d�ｋ� X���Mdv�J���K��6i�d̩hW������3ǜ;	��-@�Bܴ�u/��w�U�Do�� @��xXʕ��İ�|7弐l~8�mF��W��ƭu�a۔=�32XR��^��b��ޣѰ�i�[�M����lw[vՕ��U�LN*��6�����^�'礸�{����KZW43�ze��1YU�۬q�X�;)[����*}U4�V!�n�t{5��t����V� d܋����.7��������h��=?��s�g�[!1Gk,��Hwu]�9�l�!ֵ����Y揸Z��<-�y�E��j}���+lK44���,�ML��Sr��	�E(?�&�t��kw��~YI��Ĭ"o��LS�fc?.$�Dg=zt�N>xc݉���9ı�c�e
=T1�
�  ���c�y�2�W� ��\(V>m�B#�i����5�u	-[���svŷs��w�	�i��e������/�[�ep�n����
a�qIe��W�~�� #���.H6������B�]TCI��W�]��{��ąB�4���i#�^d���l��U�� 
�Fe1�w�����>XN�xN/��?@�K���N'����=�b�yȝ$���y?����T�5��%���_�R�u�����2�.jM�W���Q�h�h��ε�j�_0��W����Od��j9����r�n����� ��=���hxczm�QkC��W�םA��~�>h5`�r��'J2���Ę=���_�p��Pb�H>���35�����F�'SX��l+Rۓ�GA�l<�d��nt�[�*=78wY��GO���$�ɴ���&�qG`�e:����%j�hc�
����t�<cXC8ω�d0�⤪1/Q墔V�Y}�����w���d�c���d�݁V�ƍZT��^����W�dtb	('�"��]b�3�\I»���N{%9Q�a9}#���ءMbLm�I��9�󭲛�	�i�1|��{|���t����;�H�,)u�~q��	� ��hQ�������� g�"�+��/���o�>ȓ��=�2�8�?�����t�5�O��_�M�� �Q�:ז� �H�����L�+���bV��b��%�s��\��k#�e�@��h��;�1���+�COfy ��q����v��WC��z	�� �[/R��$Y&��UךɌ�')�j�e`��^�lR��s*�������)mraJHb ��pn3:=�a�ӞUzq��=b�ʇX.�y������б�ʇb���P9T8�۬�$:��h]�p�O�s$-+��S���a>�ǖ�����m�
LÃ��d���s2�sn�c��%�*4�%��l��;]O�������FQ	��Gm�qdH~��N�x�
0����&:�=2F�UESH��e��e3�LEo��R�h��:��=��2Kr����כgp���+^�ʅ�W��e�Ӑ��i>̥�����ʱ;��j���u�����0+�Cv� S�]���*�ZW�Kz�:��*ڕ����»��Q�<�kR8��ju%,up�xj|��\�-�ן��,~ޖ������\�z3��P�W�%N��:D���E��wĻ�\E�x�>&�1#��e'ő������2���w�l����)+K�
����-"�HJMvOY��/�b8�s��\�[�d�Q걪�e�%�7fO�hg^[�EK���*���TӘV�S��%��[ \��c�}�cZ\�y��c��G�ڟ�{\�5�������=g���L>4� ��=��h�<�"Y���+�>�"�3�j=�hҥ�%�O� ׁ�)z!��Ǻ��ڳ����i��G��օ�ŀ�M��$/:H���$g(��@ש� �H�)ۀU��PeטP5vAm���w,�Va5Oz3���c���pn)l�}#�<�O>�����n^��T�o��)�l�ď�k�nr��U96(SWa�\�!5>�ZL�����c��-3���}�$����S4�&j�k�(�Ah$���_�`gդ��L6ؼ��������!�9ed�{]��Ĭv��������!���Rꂱj��y�.$�qh��[� �gT�L��1�����c�?!J轩.;ڔ�|o�]����\_Vd�`�]�>*t�޻(/���li�(%g��vS��p(�g,�$T�ȥ\��2�.@�S�ʦ�*r!v��V���b� ��;F�s!4��Q�0�_�|.�/Q�>��S<�
:�gG.3�]�O��gY-�Tw���r��V���_|�<�ȃ�3 ���]������s���"6��x㻜-�WU�
I��˾f�f���$�!�G�ɇ������(h��=�f��Ǧ�)3����t�}_�G�g�
�u���E�����(��c�+�P9�{%��uNƠ�G���@μ�I;� ���R�ʼZ��(	B�s�=TO�%��ئ�8��k;��v����վ�X0�d�s�s��i��Z���X�5r��˻J�T�M��ih�N�vsm�&6kc��bO\|Hx�ߣ�elM3Ƣ���w��x��*�.f������Ս��}����IN<����Eo�^;1}�[�H\���΀�%??�f��<����"��(��->΁��T�C��^����N،�SwgЮ/l��,���aZ㧮�T¶̅��>�X��CǼ�qȟ��d��Q[9Gk=�-��~l�$��G꿘o�)�W)��(�8Pw�_��&�w|iۊ��|��l���m�#�@2K�-;�JY�_:"Ιǡ�6�k����&ԩx&����7���m�P��wfݬԃ�?]�4�$�Mb[�9���d-�y��W4շl�ú�I��G��+]����bRyL�o����C�'�Pf�RuCI��iZ�%9�1���q�._�l�!i��Z���-0��ߚ�G۽�'�ͅ�>�S%M��'�e�� Vc���p6'��q��P��U��=K�c*Hi$L��ف���c7�~KˌޣW�Pk��I,Sym�^����
`�A��7�Yki�=��0���>F��Ttfe�丿��yq�����e1jU@�KO~�f!�3w������K7:��t��K�mW�vpY&��v��u(UK�T���s\)�{�ϑ^�E�C@a�o��F	s�)�/�|bŷ穕��b����U��u� u$�<u��y���n�Y*e��9t�t(-�bJ���z��7<`<#.�\���V���F��+�#O3-�-4�[���b\n�Scd�R���{ЙĜ�)d�opuIP�kJ袤I}昷�������TR?�5R�w#3���s<+K/N��#�/z�*�k$���o����,P�.�c�"� �g�P�3�/���7�;��@>0��ц�}tUn=v�-k̞�:�5�E*j���2Q�����H;�~k� �&�M���Sd�Iك}dC�%�����U�Ƞ*��c���	-�*\E���] �J��N���2�E¹�;A㱼aO�*�;�.��3��d����T棛jsTY{�����է1�O�S���������w�������oh������_5���xEpK?=��<�&+�?{Ub{>Y6{}�H�Ֆu�f�6��$�@`�uY�3�B����=C�p�ʚ$�����@ط��~�;��k�W�y��rfi��r#�h��n�J�,~���z(������E�N�&�~��F?#��94�ٹ�צܶ�(�
Ui�sf��"�-^�ƐX�Z}���N�\;��J��k��gF@��
^�;��/������p9s���Z�TY͛�<Im9g�	�ǃ0�{��O�O�ƸbQŨ^[�>�騙VnXI,�>��E�:�-�0뚻��r��.���3^�*P(&�,5�iV��\CDn,0?�3#�Q�`�=�F��vFzҴT�PHJ�jǈn|W�갋����/Q=���{BNk��L����_����ZY	G;���Z2�ȸ��g�_-i�4^5�ӱ��sb�(K���'������{��@�i)A�x��K�+���ޏ����lR�ӈ��=i�r�3�þ��r"iG��(+�1�n����ze����0h2!��&g躯��ٶH��)�Y�b"���|�fg�P�zl6{����������\���*����<З�Q,�;��#�l}]�3NL�ZP������㕅���K�� ���D�ѕ��2�)����X�	T�%D�w�,���;[ݶ���-GC_���'i�UƀX�!�O�>X�wH�4��NV��λZ)Q�84_c�1�X��'�QK�P���ҰB��*(�����o����w3�10S�ԮP�I	Q��yreز�Z��6Bjt�����&���/��z+�#G�K��>r�&( 5~EY��㫭��_B���F�b6�%�����h�Seш���s8kW}:V�@R��68H*�<���sbH��rN�5�:�$�zm$%�:1����Z)����.��5~�C���1���N�C��\n�e����tP��PvA��1��&ܤ�Cg�-�O"��_GA�r�+��a�WY���"� �N�܌7YL�� ��w��
������a.�2��;�\���9x�B	�2�d���=�Ǣ?O����W��t�5��E�ӿk�V��AD-�WKU�`��?�c$!�	q~�!x�qm����=+��^f�[sK�ͿRKy�Ԁ!��'l�lXg�Tk/���G�P���d����a~Ǥt���V����G9Oe�^��:E���Q-�s���|�7C
xA��B_c{p="�����a�I������{�@fFNNrd2.$G��u^C��g�Щ�%*7͗g��o���M��fO�ʲ�\��+���:�[o�<F�
[tw�4�2�:��������3`[�|Q���D��	����b��4����P�K�����4��Jԟ� �D�?�:��������`�Ļ���]�P�ű�e��5
Jn�釼�瞶W�hg�L��]_��<��-$.�*����"����K���v/�OEm�m%�k]�,�^�W����C�һ��0�S���N�፤������%u+��F���$Ä'"�d4x��̋/���q�%�6ow�l��T&s�iVӖ���h���z�7���P)��x$Ǟ xx�[�~�}�0�����:"�^��m_�ն>��!��� /EsR���[��o��~�ٙ��\y�J�lϊ���E<S�%�.�����dh�������.�,�b$�(M�"����:_�
�8�Zԕ�P��/]�Vx�u��:f�Z��}��t���'�+�CK��1�eB���/�rt�3[�_����X
d����$q%�E܏%�	{��1q	I݀�tUm�+�)n`y�u"��*9"2�	��qC�D���F+�n�N~
�S)"#�dIa,+��(	��5��vI�AG��*E����O�L�D {%���H�wń�{Fg-��P�������d���H�G�C#�,��3�<1��2*��if��JEZ=�$Y@$Aۏ�����u[E�P[Gtr��ld�'%�(��eh�W��Ŀ��40}�Rcl�z��$�A�9�F�c�r�f>!��H6���Gd�=G�s0���w){V��ɾ��� �����􍥂R:��a���F�/h�.t(D{\Wywx�)���fR�d�|����᧔�x�>�>n��� �*�*Ijf���< �*���w�d����	5�JD|F"� �4�f�g������Xv�w�B�1�T, ,�oIr��1��U����&��W��\sib����꾢���_�SxϹ��s�ۣ�����g���C��!N���F��e9X3��=�j�"߁�����[��4��Mxl��>v)߿9�E�G�����B�7�/>1���X������<�����f�"tG.�ts�U�0�TR��T�k�G[F�y�>��p##զeD�i��v�V�oMUD�;�p�Gt"��V�@�����mQ��X*Òh{��*�R�㣿o|�.4c�+������,��ce�=����Xk<���\=S�:# ;@�O��X����:���,q�T��>�u_��Ig{��P�Z�3f�����9q\�H���8T�vm�Ƅ�1F��?�P>~Ѧ�S!Oz�S+��v�CoH̾H�ٛ�Z�͖<�v�V�1��1C(n�!�_Kb���QV�������2��|�s!���پ�݌���耜��l����N|N��!_[��`�Vݬ5�rm�;��`�t�'��w��t�1¹~��'J�&F��y�"����,r�����C�'�`s"�b�SL�W�8����� ���ȧw��l�6��QJ�{}���+M��s,)w0�k�!�ŧ�8��-��F2_����:��7�M������5�⯳�+���}���!��+���Ah�+A���(V_u�n�W{nSW���"t����<D��kQ���d��	���4�]�hc����Qڥ��L�Zv5�UJkb	�;�:�$~�Ҙ�sߜ76'�!���R�dG�墤t;�f���w��`���΁�������$�c�@�����9�O9�>a���~��B��^� 3+k��t��We:gN<�Ѯ��6�����͜�x���@lZ6Z�Z��/	W�IV~�ж��W8��h#���6m����t s���x��q�c�g���JE��tGǔ�1�j�u`�ޔ��	[c��X�i'vo���L&�ߖ:�^A�nXɟн�r�c���/���?vB0J���a&�"$�g%�.=w:�V�P��n�c���nS8����V&=L�$L�w
y�+8��g��%��+�HL��4������v�g�Zo�k���T�
j��M�ܱ�
|�0�8A���e��p�2l��K�ze*.W2����r����5��p��|'	��*'�C��j!*5�:=�6���*�����0�}�%��<&>�a<n�nNzB�K>���x�S��b4^�ɮ���+}�)'����9Ȁ�#P���U��V�֙7��es��Y���$�߈Fr�99��w�'D���K���2���R��ˆ�T/~s�4:)��/��|7��I	ˋ�G��` �2QgM�ܺ��ìI�����)�5�%(���,;�&�R��p�˨V-N41ݡM�>"Ľ�2�6���& >��^�=t�襤���X 9o�-�
��s�E�hVy3��w�ʤp���(�t�@���P�9�!K�����jb��o]���`*�h����.5{*�,���t���A�J���8���I��(�!.��V(B�Լ��ে�c��Mz,Uw�% *�=[1��1�&���]^����ڕlK&�ܧ�b�}	` ����Ä�8���rD�k(��Ee��Ի�=�  ��7�-��9q�~�]C�3W�7(ng�	5�n���I�&�@&\qr�w�B��Da��-��(@g�;S��d�[�j��	G�A�<��`-������rs�4���ikSm��S��1#�i�aЇ$���N9�4���WfjN�nǴ 4y�Zs�^�ј߁:��|��ד���ʋ�8^Ǹ����QS{.Y\[أ�8�g��趃z�~�d�m�d�iP@$�?�x��{*7��x�ذR�Y��y�uy�����P�6�4����%޲q�l�OH�'N(����r����������9�Q�ٞ�ډ��c6ف_[�1(�q��?5:�lȟ�Y�|H�P&�	.�J�3
��&ZE3�N뮩�+Ar ���`aNP�7�"����+�LY@�^��	\�K��0�K�����^d2V\�`'������^|�'a��7�'�+_cxP��P�0N0L�
OS��Tk%�5������ ��t�����[�@iF30B�i��]%J�12�vd�� l�i�n�Вn61/�`�-�/��K�ev�wy�'�Wu���-<�C|y�ʓ�ʞ8�?�~L��p�1����u
=�D�������jhX��㣾[�O{��
�>�^�ׂ�<91-�Wץ�P���"5m�}5���ăK����e2��4�U�1�=�"h���CJt*��� �P��C=�������ؤ�Y�r�|a��Ȏ���f�?��x/�1<�/�a$�tj��� �:��h�6ӏ{��R��c*vrv��(�@A�r�����2?+vs?`��R��Yb�bҶ<�_��X�����b9P�΍�ps$5,�7�E�p��4�s�P�ǉ	��(�bě�-P������%Ơ#"�- "ԡ�����3D�$'3Vx;�f�I���\��
8Qe����/l�٫	�['Z��:�D�f�̅�Z�y�;U6�B�]��~P�F���i�� �j�ݰ�,g�0�^�~����P�������Cc<��ki���^��q�C�[�Ƃ��?�����(�I�u �7+���f��ͣB���o��ů&���C��cfC�G�Wj�X���H},{�\�t�K��A���l�����/ḚQ��F�c�~������rxR#��V�9��1~�+C�{1�>���:Z6�:�0�o���E8_o;�ݬ4��M�R�UZ.�Y�NP�@UX��lLx�D�>�sT����aø#�����:Uw�44O�r�,��_bVt��Wt��!S�����«��J�v>E��9Nq ,]B���6��ts�:�ɶ��[mq��R�]0`�v*V�I���O6����'�a
<��3��SU���+'���Ox�!�x��S7z�΋�h�}g��|f�E|��Q�콀r3�?�遪9�@�$�y}��|8$�#�G��
R��%s�����hbI5��NJs\fR_x7[�c� &�.�|R�����-�T2�Ǚ� �e>�q�
�`�ujE4轓�dkwlkz!:z��>1D�ؐXe��d�®�wPc�=a̰�B�H�z[M��_FV�/��B�{/��27�7c
�M�6u2<��U��y{���v����sGwnk�dmJ�;���2����`�s��W�?p�ζ:��2W5�WN������	4�|�4@"���f�|4��뾯O�i��G������|��b��v�4}H<��֑e�	d���gU��}/�Q��c:�xS��򬤖��=�|���E$�T8B����K�|V3]Upi��Բu�s���*>�\	H���Yȓ	��,盄�J�IeN䶓���j+��S���2$�1���e���2�!� l��iE���K��B��j�m�y���>x ,�ё�-��^�؍|�OXQ� ��)a����iY���B������b����}O[���6rY��?@����p�R>��x�i�U[�r���z�l���>ŷ���T4�����O���2"������s��Rm��]�������WO�r���J��;�L����A��-a�3ю���@}W��Zh�-;�x1Y�8-���v+;)�<�>��̥2�tU��u�W�v)y�t��/-xO�G�F6t<q�����N.�B��xB��Y�+��K~j�e��1|~�(Ģ���%k67�R���R�A��^��ѥ+%�SOKja&)�2v���v���H�D?6ztx��4T�N�)F^�G�xm@�՟����MKW(�V�sHT{l��9P�
x�-��Ýs
��v�0y�����{t7S��JO[��3ǝ'�mj�{�9�% �<����	C&�3��n:�?�4�Z[a��ˆ�K���zm��5�W��!Q>��o)��,��8�I�acJ�V����Y�H>�p�1�\��W��Ҽ�P��Uz�f�[c����N���	z���c�?I]�q�ˌ)��6k����1�(`<�<	�-����s�4^�������x�nF��g�b9h4Q���(����ʐ�t��{��|{�~q��8g�7�:L���!��.�Mv=��Y#�7d��R�E\��BgA���?N|��*�uCJ���ψ�0Tg�I~�P�F?S�ëD+P��[h?�������I�O����P}���[�3�;�O]�U��ή�_��4�X�#�F��K.��EU|s��Ee��2M�\��s��R�R�� �u5��1�����J;<���/q����+�ۚ�sp��L�ŭh:~�n����s�WT�	�;ZgX>}���^�ڬ��@5F:�^f�_��/�V�?�����^e��(��M.�?�)D�̞@Ҫ�ZIı��,&џ�)�R6�&�`����c��Jw��U����z�~�V�A^����	-�o����68��)�!�\ʍZ�J��[�*�rh �Z��H���[�^a5�]�ʞEP���}Kߑ�\��OJ���}���6k��Z�/��@�w'+Z�w]�"=�$�P���%��)��c~ ���l���k(������B����A��o�G2D���9B�^��.�8�,慠{� (�䄱8��HK���� S؛K�C�D�y*y�`���� �1��#��=U�|��W�h(7)�p��~ʸt�J��v��v���o_}�l�VBEvۊq	h�Rq}����ֺP��Ze_u �t�C:4B�&r�@ou�D�����R
�@B:�z� �=�(����.��oo��x�Ң�������s|���))~*pC�,u;�e���������BO�g�h�?�(��h$�b��Lʢ&��K��:1 X�
����?��}d�y\{��9
��o"��̛�=`;��4��p#���o���_��%��E�Y�Ev6�Ld����1\S�B��&2�@��[B�`6��}��<��)w��T�N�%-�7!�6���TiS&uc���DC�]��"O�����t�4�g� g���*�&w.uŃ��<������ ������=�����bh��"P���<���g�]H]qR��&�Q/�Ȱ��?�<���u��o��&��+	E��	��LP��~��F�n��ԱU�0(��!����f��	;2��;;�@U�4�`�%�6T�ͦ��b��OC�?��f���*�p�����>�W����}��&��2
3��i,�.�R���uur�8���-���8̑;0�
t{Ns��S��	ةs5�(c5���ɠ�h�"��/w�n<�ì{�	��]�u�5QB!��l�L���D������[��cJ���W�|U��Nx5l�V�<t��`�"�`O�͏��[7[�!�ǡ#�w���oQ���}��~�1�S��k.X�0��f���.�R0�V���ʿ��j;��@;�UȆ���x�s+���1��y���Ӊ �9/y� 8|Q�T�A5L�Qf2و�lQ��brFO�	����XB�OGK���1��!��$}�iT@l4Aݤ	�ÿFr�)�`x
hI/�P��I�)��cwWjC����s�q��.�
�� �܂���잤y_��6����R�Rl�%��g��Q>eAu8�{A> QR��5�t�>m2X������߯π�� A����L�[�.�̴�2�K�,���|�g����<�<z����&$���)�����1�Z��E�t�z9�hj*�5���V��\��ux�2Z��U���ktV��c���E�蚝G P���6�iY�dx�E6Np
�����d�l����.�ߗ��tʷp(Vn�K�_U(rb��y�XwSc̰=�*�h�5��i�6�e�C��w2i�yC�x}�ctU�FN��q�!��ܪ����s]P�ٟС�C~�0�J�.�3YY� M	ώh^���|Y�F�Ϳ�2~�ĭ=S�Q�\�罋ZX�Z?ھ�ՏT}��B�Q�r�c	R��5aD�B=\.�3���pn#W8�`l�Η������rg��\z#��������;Pb��VQ��e�x�r��^�O�c{�;M���Ώ`;�HB�
����iXsHi n?���و���]�9L�ء�O��,S*,����Z�ƯM>n�ڭN�y 1c�D���i�؉&֢1DۿG���r��.�i	RPp�<�ZR���E/��?pP�B��T��4�h@V*�����dU�%b�;��~q���Ţ�"�v�q��w�܁����F���
qd���u�:�7c�����/�م�7/@�v(�B�ݤtF]ۍ�n  ٫�hU geg����Q����V���͜��.옾A���~Y�/�NI�M�R;��s�뫙��)���u�Z���{�?|��B�).vT��w��'Y�����M�#��
+#c��]�ۼ�c���:mOS�:;�%�hgZ��S�0Fs��Mi&�E�H]o�P[W3����GW��o�����{ŕ4��⊤*���q�����[�H�=�`E���d�=D,Z{�b�Ay+z�@r��K�ۆG�G<��P\��(-���J�l��/��6a��@$}EU/�W��z_�o����=�jc_R�ԁ�4�Qi����N��쯦�2±5�7���ƻ�m���g�U챂7H��(S~�u���1��6��*4K�~�;��.�\���O�{��G�4����Țgf���3�Nұ2V�0ن3�]�Cy�f�������������!U.dz�+z�H%�iV�PQ�J@������Ũn�&xT��Ԙ	5����K�H��oC���ZU��Ŵ���.?R��8�w$o�: �'�y	e�L�"?�D�t�|�_�����8P>��H
������Bnڎq)��`{�("��f�F&�IّR��(C�z�W�!Kl���.�
|��0�w��n�~0�����#$j	C�?��O<�<bs����*�@%�զ��=��2���-5[�/�6�>L���^AM�"�n��\O��kP�g��B�3����J�>��I*���oܾ��N�Ѧ���"���ige�2� Ĺ -V��o[I��K�
u�]ȿ�-��h�	�H��P�!���H}e�̩�q���h4���BK��x\�;eˋIhyc�4��꺇V:I+������vE���"0<2��%����x�G�TAG�̦X�輚��_\B�f�dL�0'�N��Tr��Ө�߷Y��f5!� y�{�p'D��L>���v���z�5̆��2�>���:�j��n�͐\�7���0�5�J��S���证�oa'-v�O:ҮE��u�"'�.�'�\��#�7	$21%@�lDs��]��!;L�&G�|i���r�y��m��i�U���]э��hL�t�C+��c!O\?��14Ir�n�z�o�8|n�:0�IzY��NHhyUm� O 1QTJ4�q�n('C/�X��D�/�rs�
8�.ί�&��~c���6
�U�y��z��qT���VU��iPU�+�mz3ʁ���I��{�H��Gg̯�^���Ԥ�&Z
�ŀ�4!Q���Dx��@l�-��ʭ|�-l�3P���3������}�Nc�8(4�nѵ�!"� 7�uJ
^���梼�X�e��rpC��sɟ5�(cԜE�Թ�;���&��#�ɓ���������������i-��-��7��8(ufv��l�~��<L�����p������� ϔ��F�q����r{ �H	��;��,��Zq���<��	�h��,&���Ӹ{:+v�r���Z�<a��09,eHP,P�ޖ�~9�F�d�7h�<����'�>�,��ahAO�&��])��w�&Wqkճ%�H�-	5-_\	q������P�GmMW�	~�9� Q���y=��$5�'���ݭ�n�|���6Mx�o̃Bl�_*r�@)"�X��)t����)�3�a�܃�3�M>�ܵ�t���ƻ��n�Е�9�up�U�a����#�س!���R5����n�.E�9�'���&��N����z�b���ͣ*@R�ݡ@H���זeyT�h�BL++�
b�="�(���b�����~]Tۋ]��um�q!�-V�s��_!(.e%�&��v�<��<[h�?�iB�ӧ��?�i�v`W&�V
�BSI03���m]�J�(�E|!z`��D�uS<�MƯ�ԍ�8`�����CՏ��M�u�(�>�������er����vc���J�����+r��:�m��g����1K�B���`}�Q�hf�V)'��8�LH��o�\���dXv���XFY���� ]��ګ�{�ƶ���i��5MQG�b�'��xl�D�L!�����U(�޴�KD��J���/�e���$�~�3�g��m��V���՗�^v��6%b���b�Di�c�<=g��5��{m�#�+3�?�{�L���0~Qnpۓ�rf�f�ZC�F�Kc<�����_]/Q��am9���Bà�s��A$o
h����������/.�Ȼ�̘[�~/�.)/��f�o.�[]SG(,�k^��!Q'�uhx��=��L���(8��Ga��-�lnl�;��W�����9�`N���) �-��"Նs/��.$1��)�t��Ax�t6�6�Ƭ�ڌ��
���D�>��22�K�Iyr�f#�
�sc�AK���'���3�q����Z�.�{Y�;��K�H�^�GDھ�ʸ�hL�3�]����!�x$�pxtN��7�:��9�����ۑ��k�(��� �[?�r��P�.��p��%�v��7c��|���{�Jil�Qz�Y�/7��y$5p��J�tm�c�{YT�Ͱ�ƍ3�6R�.���/-�X����&Y{��D$�SK$x^o��mɵ¸�NU� ���G�q*. +?�%���n��%_@rxa�s���,{RZ2�ө�kQ�iat>��� Ǘ� ��l�gEgθ���LC�A3?G�/�^�ivD�}"ig�t �jڵ�A�mf3��� U�����6��MI�������=��E�*<K�tF�}ͧ�3/9�<y��W������;NR�Ϋ�;(!a^�X>�U�^���ҥ�͡mS��{<��Cm���n6O?$��2u3��>���q�����4�+o3���=�E��fS��RU%Cf���!�J|���&e�J�4 <|hV:0+.U�}����a�ZSp�=`��Z�N�g��4��isU����aDPK�-7(p����ݗ��K;.�$���Y�V6�tQ��C;se!����mXDkި;3cȐ���M\�/-?�Ě�3����.��5cZ����DO�h�Yj�wQT�85�?�|��|g0ֵC����Vۗ
�r��Ί?�~q�#��v�.�ٵ� %�2�:n���J�9%���?6�ڴ;�k�I��T��?Q"nM��ZOV l�4��
z�&0T�C���;���,<kzf����wՇ�eN+s>׀�'R��WY'��OTZ[N��gR�Q͞gZ��B�it+l� ��Z"߽o��dN�Cg���]��֖������y�9�5<gb?L]=��<�*�w5�B�����5����DAձc�UǬPg���&�|�YQH_��y�|�C��0��`~<FH�{-�7�r|�H�#q+��I,�Ώs�n�I|uKnz��( 񣅘 -1(�IP��cw�����R�M'g��]n22U�/@h��� N��4�TD��#�V#����@�c��I\_Ze��!�{�Z�.��f�
�}��E�K����&c
��T4�"/l�䔀W�d*$m��N��ez��"|K*�ħr��/�+�Y&p4Lz#�P��zįON�2y�*J��G�d��r��`'s=�	� ���C���E!p)�mQ�f6f��܁-����+��� rӐ�4��lw�ka��W�Um������@\)����:C����0)PM?^�u/.��t�]`;���ę��,��0�p����_2)�u��6���Y+J�r�ܬr"8M!��ĤI<����4���0肾'HfH:��5���C��3�O	����	��$Gq�)����+�Ȱ�F�vX��z�@Nڟ����t�K��%����r���yҴ�1I���@xv\��$�Ex�����+���t���,�/ZX��j�r��gJ6s����b�<[����MH��b�l�&/DA(Ax�6͞��)��2(GkM41�����a�پ�ޢ_��es����I�R���*��� �,Y�x,W&2��q|�,P/�S:���(zWSV��|�s÷T����&�V�� b:�t���q�t/VkhK5g'
�2��N�̷
�r`[�J�]�r��nE�Į�Ϩk�@�!��'�c�F�Άx�-:�0�q�ã�����kc�E:�Yy�W&��%K�+�d]���q�ȵ���V�?�T|T=�r�jou� 
�uc9�.��9j����D�5�L��Gb0!x��H��cԕ�jT#���t҇A�跍��Q��:�Dc��oHi���կ曀=3�P3�f�7;e�0L��ed�K�b���$g5���7C
���Ͱ ͅ��ضV�HQ\�L$�m�
P�bF�����$\��]�Um�O`���/.�~,��=E+�����Q�'�^gV�������'�#/��s�;<>
�}�m����s�r���Y(nk]b��e�E^-�F�3\m��j���Jp0�0��ᨠ��/�WR*5:��`�����r<�v�<�J��'h��>��
	���3��I�hrg7<F`��i!i�}�D^���*6��|-��F�6d6���`���9�t.�R�u�_gB؃�V��w�[B^��9ʅ �/_���Ü�ԜQ��ʠ�z�<Y_�\$���ޟ`e��Xc�"N�]�"��11�t�=G���Xm�zz�JE{1�'�̉Y�n�H��^b�"��`%b��5�n�:۝��F$E��%�*�
��%��',Z�@BI����O>����]+�
pÑ!���/P8^=%�CW`�!��4��\i�oJ��(U	qwR�ow(�a|���� �ǙA�;��ph׃�-�F������VԻ�|?��VЀbL���
��|]y@v^Z�0l���`��j32��&�{�t�Hvr���XI,�5��G���1�n�	dU-p���T�jgE�*�h<��	�.� �P��'"30��ބCM��_?$���!$�b�$�ғዐ�bf�'�Y)�}���s+��4L������O�,Acui��!x�׮������dd����P�����"�pD0��Ƴ��Y�B�YYC7~��y�0�zry03�Q�� �hY<����o��@����6`$`J�����j	��6i�F�t��Z�Q�~��ջ��^���+�c�1�h�Vj��E�cU&��ӊ��H��f?
.� �!��:QKW�
%�t��d��BAu�4p��^�����J���F���(���I?�lk��w$�g�r��K ��>��;�o��� �&hI�S�˫<���}ŬE��J{j�,�n-��,��َ$�c{���i�\E���Bs���#\c�hv�a�%�5ߏ�����XKiiad6ಷ$�w9,�!<_9BB��Jy� �S��-������� ��H��5Yd�ΪD��T�eDʲ��}�u�Bv�x@�V�NgC���X��,����VC4ng<�Ҷ��;�uo �)7�բ�-�i��9ه�1�x���Z�����@�Y�2�}���[��íh,�y
Њg��.�L�J�F�F��V��gPh��:8
��ATv��Ȩc���2K{��Ć��C��&�{�����	
�v7���n"XB��>��R�}JE�^ƚ�t=��=l<�=ψ�柽C�>Iܞ`f�gQؙt�|M(H�B����ě���c��p"1:��N�c�� %G��/�	[����/�c�ݭ�NqZ�@bw�I�������X=��%����uۂ��zk����
13Ǐ���VΚF&�q�NN���ԕ�c���v(����}���U[���o<ٜ���pe@1��mj��<�c�F��:��?�����!p��.��ڿ�Y��g��J�cz :c��_�rvk���� �9������������ �R)sE}���WĶ�RVp���s��RdZ��e]V��`�ؑ���1�(>���w�ӼƏY�}y��*�y��(��\�\��8�b�����dF�[zJ!K���t^$'R�]��guF��V�0	o,&5vYu�����m�	G ���o��<{��3S������c��� �.݌?��DO��'�pV�c�(RNZ�cagHbMb���u�xi��d�]��O�]R�L�\lւcV<�M�Eb�ڡ����.E���[���ƔIW���J'����ot���$���{O��d���m��`yu�1@E�S���jƥ�������O" �_q-ԁ.0���VC���N���&��S�=�,�Qhf�G�5iu��9�e^XʃD��H7P�_j�ېq�t�)(,-��$*��5#+9�C`�W&q��W�q�r��|Ӷ1
�;|/�'&@��r>u���^ok@�k��b�Ù�ypk�PZ�����|GWϥ�;L�F�7MqI��X��t ��;��Y��|h�abD�M��d���k�P���.�`lޜy`�/��{��D8<�IQ��y�~R�U����Z���ɉ=R�5��	�F�v
�����j/�KT�Q�|������ׇ�L߬oXv��+�a2��+ѭ�Z�+���3��h���]�������l��$~2h�?z貝�\���QӖ!��"� B��p�p�6n;�Y�f�r�$p��P9��T�y{��#R���h���
:����ӯ���=��tym(˭��b�.+����Ż�[I�d��|��@�8���8���~{�@e����:fc��!Z�C���au6�O�Z�p؟�<�?�N��W���J�ֻ�sA�Ћ��|����U�e������<(~��O�n��W��K��eK��i�!�:������&z�R�neLXI�'\LA^��ń�WL�͈C�I����tW�+��Jوq����|�����ca�KlքW��ۖEn��̽;;)��"x[�?�Hk&!�]���J�(Ǝın��3�4��R�SD���C���]i�Q�o/*�2h���黗�Q�VѴ�e]D���SK TJTU�����I��}�kr+f3� ��1�U9l
��5�xo&�+����z<����s����\%�	�U���+�=z��u������d@��xP��+��W��=>�P�r0ydۿ�y�|�M�<����'f�����tWf��o�`�a+5�]�/����x��y�d�WƏN%Pه������Fg�D��Y��*�'[��&�m��L�C�/�}]�����hі�0E��<c�;���)F���' #�'sDK�>D��
>���95EP��_��_��TL�����Ǟ�}�.�dd