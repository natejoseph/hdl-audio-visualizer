��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��N(��)�A\k�{�'�&@?�<
߷F�lD���jg̮bW�ҚN.3�%ĕ +�l���?}`|':ʭ���J����A�mV�Xޙ���C�lX�n80e������KLZI9��|Y�j�띠��V&�Orb~ȩ��u��B�y
N":`A�� 
�(�,������{H!�ƈ�9�;{�g��`�+)4�hPR�g�?���},VX�+Y��;-_Z�]l/ܷ �_�����}ϩ�1���(�^#~��c�z�Dl®wC3�ꭦ�#{��8:�e\%�����I��2E���MQt F�k݀�!��bM~�{[-S�Y_F �5m'�����R�!�������q���/%�٧H�۟�O�ɜ	n��|x��$�F����έ�u���F̘S�<hA/�	q�+)(c�G����+F��U���D}+73|�q�y��ƹ��7u�9��S]����ȼ�t�y� �:��九����7��������-����*{�^ ����sU=�ׅ�A��(\�EQ�]��L��~Jw���D���n@�M�=��M�"�X�����>PLj+��ykL\`�6��0&��I/�����j�� �Uh���E?�Z]�.�&�5"�y"l)*� �Wq���$�>�`�ea|�3�E�e�>KV�����ao�R��F{���煫m���	���V�hkN<P����(�io�����L?b�e4�����V�f�m�0"��FG-�J�p�Q��%������Q�w�m5B�T���R���LP������V�_�B|<�\�%�穥�N@�z�fI�{	��5�I�b�)�' ̫�����h -22�$��OL|7m!@o�Xv v�����L�z5�'��ו�����������L���3{��^%-�G��R6n�r�6�A2���ot��&(�c�|k���&^S����E�ä՞��}�����K��A\��^k���#L��s�~�dwx?��Jv��Õ�NE�w^��h���Ӳ/� ]76�/�-��M|q����� ��٤���rxv}���gQ2_�w�>Sl}�\������+��=$ҫ�[�p��P����+�ݛ�n!��1���SG��u�����z5��R씺z��<�aX�85�F 
t�g�����D��C��Y<Xّ�7���L��>8�s�m��L�J7���)�S�����$B�k@���.-�>�XL�`�1e+0z�mw<L����L��9�.���>V�&��_�N��8v�LG�p��z� jDߧ��y1E��H�Ul�_7��ҏ[B��2p����UHAE�:��җ�)U�T�HG��������G+�^/��R��q���N�ɫ��\t��Sh-G�ͻ���nRɍhF?��J���o�+���X�����\>���}�r�'.�����w���VW)L ���[H؈T��K��Ɔ�ݕ��<+lR
q���̇%|W 8�t��~<[,�nV/�p�'��w��b3U��p��B3t�AK�tD;�3�Gf�ћ����F��t*���񾣌�-(�7hDu6����x
�'iO����F��Wg���2�ĚL��u�F��Z�S�=
��]2Y���Z��hoa���������V+rѠ��+4U� �|�����y�i���b�	?��-�%\�f1��Q�2q��F�� G�+�S�葑�䞭Al�'g�u���E�K�6x���d��x�_g5g��H>Yv�2K�&'��ZM����#�mg�56�#��l�Qj�)�:�n(<6�Aa9, �"r��,�eF���p�i[��J`Č��C(��f3����t�ʬh��#��B��l��]�K���u��7��E�'��yP�W��%�b���k͌�4p��*՛���ڄʬn�6�Xy��\&+�S�^n�{s��W˅Q�������˱��U��� �O����C-˅�M�1�#I½��`=-���j�cI]��Ϻ��uS�ǻ��Hi�� OXf��s3C&S�ًR����N��v��K5���斺��.~�����X���Gf�W��w�#�����}���(�7�Jö/��� '�lQ�_�k����<��$w:#�%!��gi������_A�G1�u�\��Pd����H
�Xb�\�ڧ	������.,�>�D��j�1>�.�<�J$�(��Qoٞ&����C�-�#��,FgX0YKbu�"'����#J�%c?!ț�~X8�����F���O�;_�$�{�ϥ��YӤ�߂�,ť�A�s�th�|I�9�8íf�n]�������b����%xT�\�5rO*I��O��oQ!F-�O7��<�4���V�vq۴n:d?�63��Pk��A >B����G_X̀f�:���H-`)�Ҍ_G"C@H_��CzysG!��+g���&e��N���5�'�5Ϊ�WQ��&�����Z��~.uPc���ι��J�%Ή Hk2V��C��봎Sj}4��ɏ��%��h� ��M���1I���sI�8l#DP�z%Rw�&��g��JIf}D�;�W
�w|S��W/cr&�䥐dʪ���?�R���c��JY�j~HG�d���P���a�?�1�e!�!UL&:�GX��RT�m�����6�Bg쥲˲�G�]�Ffҷڰ�H��S���u��`�F{��F�З}Z�.�9\���,���(=�D�h� ߖ�섦�Dso�x�!݂M�?������QCݩ��Y}$��J���?E�N$���j�O�ޔ�Vf8�������-�>{*��1[x-��%z�_b����rڋ��1/���ƚ�[��
�*b.�Bd1�O�_f���OP4z�@l"�F�'_Q$��e)b1A`Ws	z\�1�%oń�Z��ʻ�4��˫� �$Q2�eT�u�߃��h�U���P8�>��m��|���h��*��K�
��7��}Hׄ)�Z<�I'7Z�_�ß$�0��Q�)�剖�R!���Da� ��u�*[����{{ �І's�{V�� �&5��d��y� @l���_j��d��"��������]�5��5@W�}#ʽj����<|	+��Y����ڂ$=H�q��9x��[E��_8觅�c�|~�6��;U�a��LO�����
�rC���=|5���0��)�Ԃ�D���Pzu��V�O�1�[�z�C��\X��v��ͳt��
 ������tR'��%�D5wxZJ�Q��D���X���^��w��8�>gD�2!y�Nm�DT�7�2�E�bQ��/���-��Xo��4��\�S�G�_Je}����ޝ�ce"�K�����-�{Iُr��A���GS�y�;:g������h,����x6E���8J-�xb���S�� WS�WxB���&�����t�@2�l�!��%N#0=,QqA* a��Q���Mxj����!}{D�=��)�R�ڔ*"���{�zQ�Ƥb���@�
/i	���ҊX�"�x]Jx������\��	�G�)2��(|_��<h�(��E*�4"��8}#�{]��CK>^=(3|��AZq�� �x�"�E'Z�s���Py���7���6O��B`Zu��H���g����ewb�����p�u��C*������}bI��>NFf�?�	��X��P��m@΂��mM�me�_�ө
8vR�*U���d�}�P��'O����ww*;U)�&/`Sif4�^�N��w��0��I2�մ m��i�Ž&	�bn�nL�2d��v�1kc�xu�D��v͑ɱn~�:ʾ����a|\
�+A�e���y����������M{jVX%��8�Qnl��Šf�ۅuv��� ��'p�[�dxbٺz��A�J
?m��� �L�7?��PP�)��\
*}PѯA��u�:�Q��J�؞,'4���n�����57�y�/�p�-H���	��h��}.�\R�O��PY�<ߘ��"�R�;��dED��-f��n��d(���;�P�ɯ.�/������l��r�j�eI�&K�l{�d�e�r`AF^�f�qy�s�6Gn��p��q�Пr�Zv�D�ؘ����MBOmdSй��T�&�L&�qsHc�k㕀����[>E��Z/��5Ӯ\p+�1��۠[�F��89:"e��S�F2��ͅ���� B�F|W�e˜�NWGյǉf<ҭx����X9��"@H��>�Ip� �i��n£nU�8�Ł_m4^<*�ձd�k`���ۃ�"C�'	sK�J��o��G}����5�I�h�q
�����$ϡ��Ö���rϊ�W8�"-�q��F���믡��+�������y
r��/��k��up�K?Щ �&DTk��)_����ۭe��i~���x�K�V�Z)�h6##�T��dE��l�;�=� ,0��!�9x���l��8��h]�sW��,�T���W>&��O��Ȋ'����0QԶ�I�-n�	��l+�s�@�B�� � ё�tȁr�MB(�2#�P��pM˿ 1d	؛r�B �
�8	/p���X��#?:���E�H�oDE=��Id�������g��&:�Dc���M�Xܢ�7��}�v�����bј=m���U��Ʋ=A<�hWf$0����3��A�˺�8:�3������g@zB���#��&�-B�����C�y~h9�
b^��b�n�é����9��+��&2��y؛x`�zSd�F*q
����J���S�3��T����lq�Ν���B�t��[��
�S��MUf`�/_�>˛J�łM�EU���A�/��&��VQIàs=H,�g|�>aD2jƢT�*�0�؎�T{�;7*��t�yI��� �mx�Cl+��+�G�`��[��!���$�w2���S/,��d����"���({��.��m�WCcIq26u���Mǝ%`�C>A�q��d�ϵs}�$��7(L�ώ�-CF!E�#��v~�ʺc��2���|	���h%�.�}=�,|��U�4��7��j��&b��'���X�zc��"/hOj�@I��=�B�|�¶�����n�!�m�8�n%� �W~�(]ܖ�O�4
un;ኖ�s��;f�I�cS����uF��WF�X �����W�a�������P�Rk��i������)�걭���Zvu_�Eׁ��@���At>Z�r����c[��
�̒���D+��M�\��������k�D+>�I�X���Z��7�ᴁ�C&b��z�q��7��ʆ.
`ㅹ���pM���\�d��lgf�vH3ԃW�'��e))���_��{��H�����Q����W�� ���DIP���)Bw��ޡ�(�1y�J�Q�Dba�Kw'�-.E� �oa�]K�x�kp�xD�G�pnS�^!�wj� VgB�%�д≱0/��׷� o�K�����
�}L֕�j8\@dہ.9m��".de��Y��n�����7���.�p����������b�u}���.� +��D�l꛼48ʗz�m>u�.�y��S2�������SX��>�$��7��-�Q�� �Y9>��J��sʾ���ϯ�.S�xX����hm�"����:;qak*�y�ɐgB�� ��9^r����Ux��B�W��'�nxD����㿤FaC���p�Q�Z�~������Y0� u1�C���-���جJZz?Y����'.l��J�oƦL�%C���5{����J���'����d�5u%Nv�t0�[�G�[����[I�H�XM�Eڭ�dd�m�tؙL
�@A��9Z�q��9�Ǣd:3h��ۢ�ٺ�L���>jhIX�|�g�nU;�ȣ�r��*�䇊(�L�������"��M.e�-��c,�G��RƮ�hK�U�}`��'�ǽ��͔{Z�c��L��X�K�C�8��jki3�cLd�۵�G�EN5��7���|�g2)�|�71W����p��Ք�Ɉ��.Y��SA�M�P	�ȌL#��0-�-�]�đD�,L3�e��010x�~�N�~dѸ�Z�(����P�%�%�m�	��W�IQ��j���(Xm&��ݭD �O^<val�jg	�S$�&���D
�	o-՞>1H�%(��mũ��r��o��8���*�T�/$��q_@�溭P�!��9��E�U0���Y�x9�mQ᯿�K���:��=%�:�{�t�����.+�X�����)s(o�Q#V��ϮZ%�v{=���ϊv�"��H6OEE���^����h{=��f�!�(j	�����T-�Y�W3�Ǘt�1v˗H��X�~Kz�1�-�N��/[S�M^]/���3��qCve�B��J�3^b� ���{9^��ӱ��\��+w8m/I���p�n:+�	�:oA��8�U���v��a�5��`i2�@�^<%]��[9r�t��L��X�:m���*=��n}��O�t��/u>��o!�Y�WА%Y�ϴ��Ǜ+'�J���g'���f��GP���N|dzw����n��w�����t�F@�G���7�CC/<u�u���O�,�,Zn5�K~�g�P�qJ??�L�F�~��'����<'�u�#����������/�BV�b�s�X���<����������z0�_5��|���=Ö�rJ<1j?�b��g��9g��2��^�s:tj�S�\d��Z�'�z�1�CI�g��}
�f�hcO��/��u.C9�<x��@���"�����a�.7k��Z��?��m�_��?���\��~GO5��	v#��H8��e> ��_�F�J��$Bb�`?�P��l���<�m%Jv֟*��u�s�x/B.�ٗ9)F�.����Lx�#V���>���8Z�B6ad��8	ͬ(hv��)gr�;Č7`U�ߢKv�6߉Yr��,ψ��lԷc��OgO-�W�e�|�����_-���p&��;�ӑ�z�u���(�D1�U�T�t�a����
E�q���,692]�"j��ȉ��ݙ�N�8L�Q��A�uAr��.���C�/�UWd�O��ƨ�7�R����:���/6���+I{��ĂĒ���[��@ڂ�$�M��\�9�mڷ;a;�?q�&��˂n�'�5�>�M��x���ɷ�s��杏i���n�����