��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�v�-Q$]����n����9��p	�nS1���Q�*Q�	JbK�Ae���-�\�G�I���K�a"�K����Ep��Q�k��w�@~��f);��u����t~:��S�DK��X��Q	��f܋qgy�ΤZƊ�}/�r�s�V0a�K��jt)k�u�xS�I�Ǖ�����X�tA�Lw��K9�~�5Zz-���V�O]�i`,s]z�"�nE��0��I�Ϟ��:k&��)��ӎ��}:��R/�n0(�j��p�槬3��Q}�m*C��YfY��S��>����m��2t�8I�����L�qC-,k��h�X���c����/�Ud�+F1:����K�S�	!"c�q-���Pb>o�ȁ>&#f8m �:�����/��	h��C��r�d���¶@G�z�%����縟�)��[�|+�`�ä��� �\ma�����'���=��L<v��������$	2+Wu�5]��_R���� t�|�A_F���"�EE��t�Ay��эP�!k�2k^zE��o�:�ʶ�CŒ�\-��C���i��i��qI��EZ K�s���@1�@-#�$H\�r�=�^����gW�k�@r��Egk�� ��rǨ��gW��D�)6�`���M��]��x},;�O�۩X��j��? �?��e��X���'373�,�v$ԜZ>�;��n�k�Z,1׃.bPˣӛ�)��9�OW ��e
��_O�����E�'������a�8�m���2�n��wE�W�%aV^���F+�o��!lk���.r~�èz�O��]Ю� +�z�
mR���Hؖd����R 7��.jքg[[O�' X�#�py�0�����������E��Q���mp�<�~�69�ߞA��m7�`��~l4�H����ɟ����x�c͝��[�X�J� g��O�y����Iɰ���eT��������}_�A��6�P�L��D^-��Zܢ��`r4�Ӟl_���(f��=�d@A�C��we:3`@��<V�f&׭
���ƴe�dT�I�����o}u[��C�7r�#�j�<�aT+s�3wu�ud�1�)c����B'��,ϫ�W�i��x�����a�p���(�4����O��cs����S���H�
.�K�`�,'�X�:(|��Yɍ8�D��f�:ۺ��}�w�KD}�_���v.;`��<~S��?w�|�k 0��I`�!��z濝)~	kɅ�Ŷ�M*8�m�<H��3&���f$ =�M$�p������'�O@���/l6p�2#���]S�ߋt�@�ɏ�u�D��(�������Z!*�t���:���4:2��֏���f9����i�����F�g��0"7$S�6�N�ݗ�΄X���b����Q&y*Yot0�Ⱦ`G>)���*ܨ�鏴hؖu*��2�C�г��tG�Y�+z�k�W:`>A7T+�W���UltޝzHZ���8�LCwd�:F;�;�*��!��uۃ�u�ll�b�&�
Rß������o��gZ�Q\y�~䉠+��p��$�S����6ɭ �5�K�"��ƺ����0`��?ض-���cզ}��;M�9]�sQ{��xY~5�9B���5�.�����@&���{��$[)��va�uu���n������H��XG�]?@y ����+3,9��/�.�N��^э�$�v�(���&���GiC!�\@IC:
���x"� �4��sF�y_]���u�j�,&+�㕕Ky�,��;���@���ђ5_�<.g��di���B����^�¸������P�7��E�f�|pj�hu�X�m�S��6�L3>��٢��D�E���Y-x�z~4Ϋ�@�B�ba��F����ܬ�������~:����{j�\� $a*�l�ޝ��!?��G1�b�8KMt�[4�:P3<���=��:���a!NrS��iկ8�`���JɭyZ�X�bp�U��I�3�n��BP�B�r�]�<�,�J�Z��<w�٢%���Rz[Ss&��?�+���Y�ه���M#�'�)���5BI���B$㶳��b�s�^ތ #���b���
U& ��Ot�~��y_������@�/�0Pb��^-����/Hv4E�1f �W?��aպ�vb''v�G�:9�a��>�y��En��>!�p��-Z��N�4�RA�m�Au"?G����3�B��X-�n�j~�[�j ����g8ƹ�������J�5�l��0��<WH���`�Z#���e�d��	�"�f:u7N���m׊��2���Xd���c�e����P�~ ���������!7M�xꖒEM�xz,m�6B�4��*����Zf�⢌v��⭀W(Y�QW�{�5N�S>�B^�QS%{=G�e�%'�m������N�2���p��OL��'�>���ʨ��:}���-���XJՂ�;�}'�I�����V�-i�AC��[�L�WV�ҷ�e��c�)r�"�h�1�Lf���h���M�3᨜M��6\A�4>��;��p\K��Ga�g���G���t,>��lJ�Ph�
Z�y�mT�@;�m���+;J�"r�|����ò(Y�~ �06F��d�h�x $c��~"n�O!4[�����-%�C�$a~�>�7��lk�f��1�&�
Ĺ�)nX���T�<�y���?
� �D��q2�h�]=�yxoV!X��7al.���/qNX\�1������W���k���K(�8Ɯ*��[I���"\�9������=�׷�_�暖�V��HE����Q���_+β�`TXRd
,h�����[����ð�w,t"��S�[�7��o�H-�_J��;�RV$y�f��ؠ}W<�c9N��"������ʞ78�xԪA]��s���k������=O� *t��Z�`-�s: n�j����" H���©����1SAʅ){�����{gx����7 ݃�ߨs�+߱��r7��?^�h8B�S���xʦ�$x���^y�r%n�$��{� .��_�H�B=����h�֜n�KQ�D�W��Z�<2�	bL|<y���[�Y��*!Sxd��b�,��8ζ�7�l� ݩ��+�k,�,������C^ݓtc˵�ؤ'�>9�?�\OY������ L��ԍ=�+v�.�n�)�1�u�i�h$9,c��=�#:�t�������(���{�Z���}���Q�'�6�/Vũ���X�M�t��R��|8u�L<���%5�т�^F^MV�����3�7�#���(<�	�6�^V��6NJ��O��Ж�Ͱgn]�C/afC�n�n�.c��5!��>�p����(��-ǳ�1��v��������^%r	,4�V(��uIO*��4n���aCK���>Tt#BO�?/c��2N�Q(�	 <u��:w��H+q�@�]�C��
��~cI�+H�ג��[ �?����.t]ݞ�5i5P�K�'��O�Ԗ��˕z�TW�V�t� @񋙯D�rwf�W-�Ph�m�qt-(b�%��f4�~�j���@bY�)bL~��4;d��=��C0h��xpS�ee��r�y��@g"7e�\B�Vl^�Ӹ��&ű�Z%�j��]p~��C L�(�M`�2�48 �q���Z�=('�8�"��`k]�5�m���i�grvNƝK�O����*k�3��R�ָ�ĵ�&3��5}HЛz�4f��KNX�u"~��]RȞ	3�ሺ�o-?�1���A�w�d4��gVUW}��e]$���/]]ʧ6eF�ܺC�j���~q�R) ���w��r��E��YF��ң?MH?pG��!���&�W�ybk��{�j��AD`1\�#�Y��WU3ݫ�1bĚB���:�Y3����j��9�S�G+cH��><<nR-q'�s�Հj�=���k�-�ah��I�\�ae28�B[�&���K�ڏ�����@�d�C=��ò)��A�"?ss'��a���#9N�ӯ(hێ�Np�+�i�;�%U�I/j0#����%|�݊:o6�?
i��`Nū ݍ��<����,��8}u��|@*��²t��L����� {����>��UR�y�3�T�N���9�����ݶjX��α�v�r��U1���8Ł�	T(!@���S�P>F7|��drZsU�8p�B�J�cfⵁ&�t�t�u�[u6�o�a+�f�c����]ߐ���Pe%���s�X�4I����7�P�Mկo�%Lw�����CM�ns�e1��ؘ����j��#�<I����=�Ņ�ӷ�JA���^����wٛ�&8؞Ykn�	���^}.��"�"�M�jy��e�fm77xG��w����4]cL�j��~D�Q'Uw*R+qސ=���|�OD��?�Y���G����M�1Нi�p%^	��"�|)�r����G�	�8�=~�������k�cS��?�����yƖ8._OL�;g��b�QJ�D�@�I���0}�tc�0]��Ye�V��[Br��`�zֿ�jͬ�ɼ���ۣ��/jr@��C����]q&M%�|V�F�^>�b�R�q�HU��Q�?V����0>����{ X#��u,����5� ��p�/�z#h��%�;ĳ(q���Q7�~�쎇R�Q#�SS~�+�o�C�cs�I<bC0!��^��z�>~�t/V�����֜
f{jj��9]��Sط�K-��k:|�f���_1�_ݍ_{
�
�R��ث��1V�*�(m�m�#8�n�4T9X�I:������ɤ�!�z@ `f.jm"���"������j:��gq�6d�}��oz��G��K
�u�[�[��%[v.�lK[8���B�U�SK� ��u��0��N��mLKDtT+^*�G�ӫh���k i[��JH����I�\�&���N���Q.�:mQ�C����ڼ	7@g�Ά>$#�d���"��FY|z�B>w�<s�s�� S�}��B��T�S�Mn;1���