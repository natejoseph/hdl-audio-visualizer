��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N�����9�'Ƣ�ڗ_��8�6��?��(��*Jm"�_�kD�g8���L���(
q�۹?�>N�9�U"��1���R��A�fa�5��9̿�:���Q�z�'�n*#>�~ $+�C���Git>���� P�f�a�cTg�Trv �A�q����
x(U"b�$�-C{�w�Dk|.��3\�4k�z=TK=�H-��*�v���xi��P����i���a����6�Z���P$�hIlP��� ����)�N��,���aO�/w�M�Z�����:��j��CI�v+´�e�F4*c���`hś��2��	ԻE����\����%�d�TP�	��(�_P#��sV$��t��C�XeK`6�v���lEȤ�JW	ĺs��j��Ů�]�#�������b}��o�'�S�����?�%�=W�J����g�	y�Ь��̳���Uc�4a��4j�>Ȣ�/	D���ѷv}@���"�4yt�����k�� �X��c|7�+mAg)`݆�|�5�͑A����Tyd�H��(��0�N65�]�X䦁i�:�U�x�����	��0�bn%3$AB�G����J�Q~VԱ���b���h�2��hF F(���I��J�Ճ!�}����O=Pr�M�m��.!x�ͧEIٕ��Ą�x�|�jw��ҤK�2�ޱ���D�!�JwUX`&./7�\�4	��s��xS��W��7���,�1tR��*�oo��>P��h��Jc�$� B�s*j�KAޯ�e[��7/�;�veĞ��d׵��=I���7�����T-���;ܬ���he^6��J�ȿ-�eX�����z0LLja�J�c|���w�'��3urU���
��L�Ұ�po�M�� s���Xد�lg|�����Z=߇%�p�J�NR��&�_�&���=�p�����EN�Z�P���W���p7�u��V�B��W%���C~��CdE� ��c�>�A��m�Pe��sڃA2���'�E���}��%�r�`z�W>U�W��ex����l�q���>�]g��~�X��.3�Cn��-��f��)�ɿ�d��7�,�)cM� T��T�{j��1m�����~��%/�Is��\��dC�?��o���oj�=o�F�(��%t���f+�����v��o�Z�0�Ϋ�O�F��)�̯�md���׻����rI�� Th�� g���q87���X�o{���D�0���K^Ȃ·DKA-쾠go��F��. ={x]�0;�b�9����� �:i���ѕ�� I:��Q����|�:��s<O�T���k
���`�E�)7���]>���Č���-O�>I"u�i}O��	�T�5�������"���A7ޒ�Tt�R�g�y��� �2��O:���onr�Չ�2�c?m��a������3�V������v���K��·���z}��B!#'.z��jBkLc.u��8�\4v�q�έ�@�V�_bO���C5�T0,�@�!��@M��,̈́-骉��o��$l轧��1a�*<��ܔ
���lR|y[�"3��B`t�/Zj1�b�;W�
x�ܩ�J	=CZ����I6��_]���\��B�U��%֛Di���h""J�Pï�~Y�4����%����O{�c?0��&��}C�# [�惇!�8��3��c���eф���plգ����w��h�	T8���[�NX�,|I[uG�[�VJ�dSu;���uտ��-�m� ���\��M���)�Iч���VI��m?J�H쮡$�s�K��׈�����Q
WJ�h𙕺��7<� �|`n���Ѳ�zh�+RIO�M
�!��l�On�������bdq�H�$�@��
�G�Z}o�|�*����q�8)���`
	��D���Ѫ_(����A ��։G��?���Όq�H����u+�kЧ￾N{��%���ȸ����\Rd(9�=�- ���j�V�
��aC)���PF���Q�N�md���-�����]�~�-����v�?<:]�f�0���N���yB>;�����80�����	�9k�o��?;25h���hc�Ƈ"od��-����(�1TW����~p����5���Ah��Y���r1��@��x�K��fB;�I��Q���Uܥߌn�?��/���U}��}������l8�%J��.��*<�!nQ|D��6\�q��Q�ԔeK-��U%w1�\u��,��R��O��JPܳ�H�5b� -�b}A2��#�R��BP��H����m8��ϝ�HD<@��&��{:�){�R��ye������g�j��q��L��A�Oʆ/�K;ZER��}=�)�2��6h�Q��(<Զ1����@L`�@_}�2��&;b���t�S�5;2nT�2C	#� M�84E��}q����%N)���l�ʙzܨ�f��6�v�Df��PR�C�Ƣ}Pmi��.`[��Pkpr��qsm(���	�ǹ<��yz��y�`�l�s0���
3����C���@ƀ���i�f�r6[��t�,Gj��Z���P�d;�VW�+>��"�U�&��8���h�����x\�eYO�c�]+C����E��� ��inN2�t@cex�,&B~�d|Ǘ0
:ӥH�e�������"�,���!��]m��R�`~��N`��
�A�sל[_'?�$w���^	�6�_jٮ�9��L��v�z��+�N�[�8�� ��(<�)��g%`J�FU��u��\�V��q�^!���8�pG��B*D��H�N�EF�����~�U�+jî5��$5�h��sp�m�μ�Z��K#���#S%׎ߖh��9�R��j2���$�?V:��t؝O�u%a�)� vĺ�"_ ����;�T��E7U�\u������^�/�W�����0����d�|&�r���0�Љ�yʉ��>����AfD�q!1%�^H܈6��d���c���c��'�5�/�fj��bUݲ�?�I������|���g,�]��<|�@�jQOi��P�C ]Z��P���ʿm�&��H6Ƶ�Zz��6�� )�w�0��{�/�}�*��_yc�{�N �f�.J��]ᙗY��X�b��hM����ān3*�&�8U�����moW���ũ|�	zݳ��Q٭֤���2�]:�����g"����A2Kk�kfE��{AEov��f�$ĭ��tb����5
�N$�K�:��{�����r;�V���w��I9��F%��jF�"�#<o�$l"�l��缸��)נC�KMR \{�`.M�Ssֽd�FS0��
=g�/����i2x,$�$w+6g��賽鉬�O��{$6�U_��hp����so���)����E�������
��u<U]Kf��Q
���4������F�%�)�>�h�p�KV��ͫ���BK��3��)��K�I��b ��`]^(��SE�a&�#*t��[R�o�]���u�Ox��Wݸ�t�$$�#��7R�;�O9"/�ᚆ�'�r�P�K�9#@>ˤ�m��Ԩ�"t��,r;�0 '�Tוt{!2��b��'��g��(�!>$����6@����8"��'-�j�m�#�����9H�oH�rEn�a<�V������5����Otzr��k�C5`s�5�7L��qm����|p��N�gŞT������-�V��@��he�p.Kz�V� LJ(΂��DL�9E�sv-ɂv�����<�H�O+b�K����#�҃���G2�b�v�!)\�"�݇x�d�����S��)��%�^c�{l�*�P ax��Rp�m�ShD{���D2�g1 ���%�GOl
�����TVȎ1�[�J�VqZ�<�5��%�"�݋��1 �|f��Y^�y;�
ܭ���'S7�]���?	O��z��mu��,�Us���9{ck�,:���x�$��v:9�`��]�����OL����ڥ]|�bO�5F�w	e��ߖ�s�y��6����Y�Y��K,ՄZ�3Y��p^�zP�߁�iL�E�j��S�`����+�^p`%i�����)P!�R@��UU'��c�5�˓;��FgS@!��]O�� �o��DO�N�C�wUr�iB,\w�猥ȯ��|@InX�9�w+L�1Z�R=Z"����A��l���fh�����F7/�ˁ��٬"�^qqè,O�Q�m�]�#ֆ��҆k}W
����J�cJ�@ ^��1�я�ˑb�����&�a�)��K����k�H�,��k�{H�y�P*�^�TzJ�������J��B�Ry��G���=��f���!�+Zj�ۧ5=jT$j�)T��h��td*�k��9�?
����A!��%*�7�N]����h<y�\�L��pG���O�7����C^KR3��9vX�!1�3U-�P�=z����!Ld��"�.Z* �c���x��G��P����ȶ�t^� �5�?�=���
u��@"2\PVH�Z�O�o@�������&�,N��H/�N4=��Aۘ|x�uɰ� ����4�)O����.v����ϟ9X�K��\��s;kO�gU�?D�����3h����\�_r�5Q�K��R��gʎ��L���^�����C	��N=������W�*uM(Ln��%�l#O�	-*[��Y�?�a���F>�2gf:��N�U��[<:N���Y�M�54��ͺJ�S��q�2���$4^=��r�Jc��h��=��>W��F���`(c[~s�a�zX������M�0�e���F���;}�X?�< ����Z�3�U�s���b .��5��aSd�_��uё��J�tH�
��g����G+[�:���C쯺��XȎ�w2�B��������+�� ��m�� ��%�	kY�1�N�(�P�^
a'��"{�Gy��� ��J���!go�E�n����7=��N�8��\8���j�+��o���˗���b�7��
��>H�+�bƶU[�g9�����5��ω�-lMZ�+��6 ��|��q,- � �9�dl�`}7e�XL�_gֽ��ؾDPlGr]_`$";ވ�C2۩�by��s��:����s
v�ĵ�v��P������F[x����Fc��y­��I�"����}5ǜmn��ϱ�;{nh��"��r��`�:���i Q�$���CZ|2��# ���ZL����MC͹��`���L+7�iO
T&0�`��߂*.���`c;�"�d^�ɐT?5,D�)���*�X0�E{ Pc���0b k�F��PH?X���Ëa���q '�d�J�~�V�|�3}FزN�<���i��m��оfK~�/��u���L:@����(���Yͽa����å��<J����2��Y���)���щ�B��{0������<r+�l�~�Ϥp<�v�a��Ð��� չV`p�&��0�!
�n�v�:�A�4"�iQ��"B����+��*�H#�#�3,��/�GFT���%]��b���I����n�-�Nb��VEX�b��D�g������O�]T�!IN@o��=R�V�2�R��iiz������$�r��!6���õ%>�%�UQ~�0L���m:��[ױ�����ԯ�4�[��'Z�͏#ÓA��/�H�F#TzK���ȩ�`�f�;%t>v���#�~X��h�&�l�-.4��U����+)�+5dm��(4L�S��#���{��Y��%�`;��*�7/aA-��I�����m%v�q��2�L��x�É��'�g�(�_��8x�~S|Z��H�ح��-HgrHjE@���o(����"���r�SE�(Ĳ�|��G}����+�K�[�L�1!�q��M���mǋX�eQ�UU91%UeO��v��F�!�O�3���{�.,�>�8���]��R��r��)���Ґ����>��%;'ӥ"�&��P���S���xB+�SjhS��uU߯~F?��T��Y�ƴ����.,Fg
�5f�﯎���5j�{b3�=j�s ���L�dD)�(E�\C�E�ʍ�d҅>7�Vn���û��_� HM�m]_&>.�4�P��{�����U���������:��X;l�)�Pԋvzf�|d5}F>Oy��Eh�eG�%��*��I����-�kyo�T��4^AC�����p!_K����� l�4�����[�����\-���L���Z��Y׎�v4x5(ǜ�Z�o�8��^c���kVEdo/[�9 �W*:�:��b�0�h�7·�K��]ӄ���.�=��&�ߑ_i♟{�"�Gf����ŔL	����kA�:��8Ҫ�eɰ'��͝�������Ų��(V�ޡ\����Y�o���H1}&[-[�.�V�njR3��>O�$� �H���;�]F-{Ro�_�5�ۊC;n���?[)Y1p��5�Q�N|���4'��|�����>��#!g���d�*fV�i\��+r�j���]�b=��κ�|Ʒ�\�F�%�'�M����s�>)��
��5�Y
gnO/��]5�����w�hU��s.�Q�!��𛉱js���fW��*E>��c�@i�CC�.GB��K�@��g�����H�9�TЧ��J���"�M�]��/~��xҁ�H(�(�O��`b�0
QT��@,���v���L�I�k�)�֓F9����S�	����^����H���	���'��A3s�O��6�~)�%rY�>o�y�QʢW(cu5�2�騲9C,	/I���Ҙ�\��`2����,xi��B��,Z�fܩ0qw󹝰kY��=���]N�b@@w1
.k�M�{�S���(jwo?hğW"�k��+;�&��ݪ����e���Z~��l�a�Q�nV�?�%����\hǗ4�5P�E����*��>s���0����?m��\�%�ׇzbB��Uh�E$v�A�2s��O�JN	T�%��V�c�Z�7�㮥L�j��H�Ü�!�����7
�m�U����������8�hI�F5�&!� �I�RF�JI��E��������a9�e�ƪ��������b�!������H'�����R\H��[d��0'.3.�l}�bW�v�=쪩%����@aD�Zz26�D�-0�ǄB��8"��閅�9��M�z�Di��
�KΊ�bUj��Q�?�E%\��/;��?�x�+�����*E`4(�p�n��y��9dcW4}�i��\�����'�CS�6f�hC踉y�,���l����-����ћ�=�Eɏ����đ����{���x��;��x^pGK�Ҵ�sq5�b�����,�䍌���y�� ȅ���B�9m]����Q	�1�E�~-}Zq�0Ѳ�͂7�];|	o纃�I,#"��%k&�?��$5��?����St-�����P g5X����㖶�K�q yo�s�/aˍw�7����	�拃���m�/0��͸��7�Z��f(Vy��F�8Ͷ��C�xbu���n'�V������1�w�v  ���$c�'�B8[Ș �pY�>�0�y�8���6���N�?c��|t�C�N�@!��z����U.�:�QV�.�����o�:���e����NpЩ�~����.��}>�i,䂱	�ҝ6��|�f �̡V멇�r��A-#(M������}͋L@Ӣ������d��9���������`^�[���]�H��u��N��ϒ�2n���'�55%mk��^�:�He�4�M6�zgI� ��β�*��?��x��x��+,It5+�����5�E��X�-l��؊�����ẸG_X��ԣ�)w$pנe�`۴ώ��;�f`���@[�쩠C���xVm|�(�Gd�C�o�����s�[}�Ft����Μ	j���z��)M���G�!neE�������x�a�.5Q�|F�ʚ�b?x���ed"��B�L�OCҸ'��������Y
#Tn2�%�o�@A��F���Q>4*��Z���$-� ��^����o*�B�ae=��8�k �U8�b�揵W!�f�vv��}d�3z���H�8/�����'�(G�E`eMd�~i�h��ߤczS��
�.5�`������o5iG7�Э�tN&����5��d�$!/ �o�`Uԥ/�j�Th�F�&��B���ͺ��kNŢ9�a%�xJ��{�Q�-���a����� ���J��U��SO��9�ꎧT��٠ʪ�Y�$?/v�a��x[�~��a�ʣ��ʹ�zw6r\3߅M�����*A</l���Y�بX�zDN�E�5���5g=N��͇>p�ꄴ%�p���3@%,V'�T�٫�;s��b��Ѫ���M�f�9���_�e�+��auF��$���|��'_��.ۍ	��.��ʲ:�#��O>����IL9#,l�܇�τ �S"�zUJd��w���4W�n��Ǣ�6�E�ca�N�	��T>�u�J�`;[����H���G��4O}N>��5ԋ����d~��P��Xx5/��L�� [%��⤎m7<?A!�{M[���^Ұ���:Lx����Z�M��p<�i��i�k��K�ü���7��X)H�i���c��t)v��.���4��UԼW�
�B?GCk�� ��[���w���_��q�%K���R�1�d!����!d��Pء�V�/����KJ��`Z+
Y(>9'��s�c�B��(����֍5���Q��벍�>BI��~TI$�z�W_��t�������n�]���ٹ��CBp��<�;��ʄ8[�HB*��'g-����^�����;g2[ޱ���'�>��<��&,��Rra�V��d{��?��ynf�w��&�*?x��n�y�j�hMŵ�Vn�u���9* ��`��f��9��Y1�0m�@<���Ě6&��8��@���N ����R�Q��5s�]E����������0��UCȽ�W��:�Tʡ�[��J)84��))E��f��N�n�9nE��DfdViqΚ��D�M9Xg� n�0a�,z�I�
�4x��Ɗ��>�^A�rQN�>��?����������1:H��pRy�����A��ZI�[�|I+s�O=�O�*"%��r��d%��V��Q�o�;�ľQm��u����%!���l�R?�vH��m�+ø�S����gp����f��X�`�b�6G��r����9�����aO\aqz����8��d%�S�)�..J��0>�wq���Q��F�&߻���8�]6�s:��3���"ɚ�4Kv��K�w ����(a>}�^JVԇ�m"�e9��Mi�u9���I3=%�WQ�L��\��3�g���q!îAvi�X���h����~�{_�=�wm�Qx���\��>���5+W�LR�H>9�������Y!��m�Z�i��� ��X��Ug�?�\������k�j�F��_\��?��ja,�Oc1�3-�檘1�Z:��ï�5$6�*_����&��٠O�b_�5x�s�L�rO�m�\>��ʑ*�6�U��1.��h�����HԌŬ��bܷ^�#�<� ���%<F>�?�aAÔ�p���B8�G�b+p@'o.�/�! ���ީ1�W�y$���A�Ō���Z��Þf�P��)i9E��e83���Z{h�}��&� v�-d[Y�]�£��U���*n?��Ex��g.�6d=O�w��uw��������'����r�24�
`�,DѠ�h�%+,t�=mP��w�
٨��f�[��3̈́_
��v�8rо4�p�2�,��
�֛�4���������E���K5�M���>�HR��"LO��ʍ<3|q�s?e�iB��yK�"^�H<L�w	]���Z�i����O�C���GR��cz.�S���GZ]E�*&�S��}FU�=G	���|E���ڹp:'N+H�Z�G�#8�a\\.t�Vy|���?��JK���?�x�����(�c}���3��y�Bj�KU:�.�����z�m����5w\_���2���vϩ�f��c�R3(��&�Qz�7;�-I(>�.j<�Z��fd���SK�2��My����*4x-Mǣ���&t^����8<b�N�)����v���f�eJ��ǲj��� �R�#N�)�ɭ�s+;/�%R��}�.��Vso(o.�"d"˃�J��;�[V�@�O�?8���+@����s0��gf�W�"Ү{O� h'�Yv4r娉W2o�Z�\g��i����nr+鍩�2�������A������G��nL��[� P���Վ�m��� (g�r��چ 磗۪��U������0	�p�������n����K�;uo6v�~���S�ە%�����Dl���t��O7�Y�f�������`|���)+��v��E(r�Fݰ�cm1�B\�bj�w���Z�J%�n ���L�+}�zl_��,�D��ػO������E|�D�Ů����e!�{��0���|  ���w�lEH�溡� ���CaW�_:�E$�'��@ ��|�Frn�;��	����?y���j�>]�%3�U6]��Rn)��wm��s(9����4m��g����4�����L�_,'jA5ϧ��6g��<R֍��-��o% :@��pd�/_�Y�F49��aŘ��`	�T�.�f�wb9R9��;��Uǃ*��<����0�1�/�OBK�B��W���m��YO�c#(����p������h�H?��z���j��J��gg�� �;v���*�4[��L�5�>#��d����9x�g�J��:�?�9���4̎M��z�t��m�'���Je�m��jF�a���E�ۦ�>���X�/��ۧ���?��M��(T��u+�Y���q�X�ɖiλ,��=��|����W�;0�R՝o(��n�WgC�ZH� m;�8ғ�e+�/\�UE�$��)y	m��$�_gx;+�N_?6�0��d��n6�-E���]�G�̬�X�J�O�ֺ�SY��P���#��Z$(�oj�E8JM^�]�v��I�ͱv{]�F`���h�ex	^�#`�D��b��,��&���FM��G#]<��2jAE�0�\�緑�/G��l�	�{/�\5#�5t���U�89`��O����x�W�6Ͽ�V���5�~�17��e�|�|���V��v��q9?!�,�e�~d���nydry��h��
�o �	�Ƙ�䠪��cU,�#�G�� ���n�y�&�[Mjb�Z�5��x�+���t��[���YB��WY�*���s���s�� �NZL�T�#`��3�� �\�U��c���D>q�t���Xw�J�:�A-R�ʩ *���\ē ���i����m}��l�Ѧ:����&�-�%�n�,��4��de��;��h�3�Cd��Q���[���p�FW ���U�������Svq�jonۣoV��χ��c�=��n�_ވ�6���+�.Ϲ�lF=Z�f ~ç�YEO�\k����I�H��� ��x��O�U����x�2�y���?��',cR����eA?0;�]�"�*�9.�X��A�-CPR0��By�>�.ok1�&���(떦�ڢ���b��5���������΃=e���38i���G�~�+����A\��|O6��F)�o�����e�u��z��wX�#�'���W}���ȫ\T	.0�&�#0�8��t��uM��B`כ�M?��6��/�<k*��߰6K7�ڼ�`%��w?�y�d�
5���V6`(��r��(�=�ĈT#,�2�5�2���gQ`t�\��z3*p��ε���0I����^��Gut#�-�IT;8�!�Gl�|��
�0�Nfcc|/�
P�њl���-dg� ܃�j��ϴ!Ц
���Y����Ix�G�:bq-U�r�:����U���roO������
U�$���F���z	h���2�����d�P���ws�DN,�w�a]�,m��d*a�=��Q��ǰ����.��%W��������*|���m�>/=���b��6S��9!�I�&��揈�q�w�O��'��0)��	��|�����6Zs95�Wq����g��ѡ4ބ���
�ͯ�:ˋX�c��ǰ�3'�Ʋk�w��
F�"�i�	�!�4�1E%l�n»�N�6����V�Z����~]��$ϼQ�\�r�U�\y��]2�а��b@Gم��N��喢�jz�>um�ucmс��j�@��j�K��|�>�hdz�M]墹ɕ�8<��;��A	x��蹾�a<���/�v���_Ɖ�`~zi�DL"3�O�_r,<w�>�RX��7��ș"P�������$���\C �)��FlAWD��h���c��L�VopYF�.!���!�Sw�[(j �9ER�v|�lgo�<����UC����PR���	I�Q�Y�+O�LgL���-�^�;��b*˝����Ql�`X+�\�(&�,1 rN�v�`��g\do�t%M�}$��ADͷҥ��������_�������4���7��#,�R�I~������U��c�����������V�{0���¤�Pۥ8�>aW�-n�UX��xN�����{A��>�� F�gĕk.��L�7$�)��� �ۧ�<�(�\������z�+��壶�|��Xd�����z�u�?�KOGJ���*f��B�D>W������$��MwH�>h	�W�8�<��u���a�_��"����v��
'��@#���dK���"�C�m�/�Kt����D��Cm�¸|��u��4O�ƱK�rC���V��h�`6���G�#�jQ�#&tz�T�� 4[�*O;�5s�Av�ӏ.�	�.Yu���=;3��I����Fu������#~��S5��*�4�}$X|���,d4n3}%�ў�$��;��)��l��,��������'�޶�m�+P���(�X���S�m���I�r�.!�#I��Acp�q^�%Uy�P@�l�Ay6�e1�veH�-%�{�z�~54���b����~5#�����v򫊐��(a��~�Y)��?}�c��М����)��N�%��2�)A��n)^�|~�u�D�g���ʴ#�;6xJ���	�o�˨�>�N�)쐇�,��q"j�y#��������\v��B��T��,<l�e�R��bZ��Z鬣G		���A���:'N#Hޫ�Y�ۜ�f1����Vc�XXr7�3.V���B�^��A��j*�W5���op#)αL�����^��gd܅qh5YH�0�Cȗ���֔�i#U��}�G�[�h��c_�sl��Ņⳇ��ꬆ���"�;�֜��t��:�ۋ ���������Be�m�7+˺�1�6�{;��i9Z��A���^j2TUb� z�j_�w&�u��R�?T�`r����;e咷Q%�r�.�j'�N�H�{��B�i�i��!"*5��\��l�I�j�|��(�h�io�`̽�D�����Q��-��0"Ņ�WN��s���}��NX�R3ϑ�!3)�)@��4��F&�9q����ŧG�J`�R����v^�����F��Ac�Q �@Fҋ��ceZ�?�UQ=��~�o�h��; t	��������ew�� l��a*N`���펀n��݃G\z���y�s-�0C~\��Q�$�ђ5ڮ�.�����˄e�����7���;&t���V+%'G�Kg?�c����Rf��w�y^�_��4�Gf�Em-+Ӷ%���֮25�6���o]��hDM��ﯓ�Rv�馦Ld���w��̸����� iAW��1��"t�2"H����?�I$iX��B�ÌiԿ	' 	�/��T�q�Q��zE�����6=`�	�'�A�'*^Bt�	�2�pZ�#��=ζ3�u/�k�S��/��Q@8����ӊ��, C�@!2�$�(ܭ*���&�Uc�h�"A�����0�eJ�^8�0h�3�y�h{h�e�1V�>�R�u�d��!,��H�r���C�?�<'	o[���u���1��RG��L0o��dZi@�H�����RdX��q؁�|�F�N��/���"���f9%��˚�է�kq~��`@�DIW��d^�y��
AV�B���Z�IFm	䂧��P�	�֓���a�R=�r��?�#vҜ�'���n]�y<�`����'H�Ke��ߨm� �^�?J%$�(�+5bL;��"��p	a>s쀖#��_X�U���e4 ���q��tl�B>��ϑ툞r*�i3r�n�z{����U�lJ9��kU�ص�3���Zv]7RJ-)����jg�wֽZ#+wS�DkZ'*�q�ʆ�:q�Ɏd@h��az9�z�U�%+q�����(�}h�?�q_���!��D�-���pŁ/u�[�$F
�g��X�s����ńj�?���h9�����5:~�T�v7�լ�^.׿J�OH7of*������������,��e��%ܡ�E���C��d��-:Ǟ���R>����Li�@Im�� ��mY!�L�/ObU
��_%N*\�/H��l�w�7O�D!Qx��xg�i�Us���+E]E{��>RКn޼@"d��^���N6C��J����~ol��P͂=�����۳/+��X��ڏ:hv�Љ�������xC<�p�p3n9켖:Yv6Ňʊ`\�3���=�EٷO�eG8fo����L]� E�@���Ǭ��"���Q�E�O��x&/�R��@���β�k��9b
�Ǉ�-��/ ��0{���"�!\YM�����z�.��j�J��J����F�����K�چ���%��A���#+���o�"8���M���O�ٞ��Q'٣��M����ݳ�1J2���B��i���*��߼���G࿶
���SV-�)���Ĵ������E�B�b���>�P&MYv��+��_�l���7�WB�����z��5�e��,s�K-,�F/�u ��q�8�r?�Ņ6�J6,d�F�H�e�%Ac��z�o�@�Ƕ;�W�̓���C(�Xܴ���D��xLU-�Ϧ/��%�T3��[dV@Q�����w��H�~�0�r$�/o#��ަ��W��3�ąݐή����x۠��V6�� ��c<-��<[�D��X��w�v^pI�Ĳ�׋0��I]�U�6y��z�ٕ	^�<��5���@O �{�1��(�_�I��bgz�U#:�E/�h�����P���7���@:W^�#�+Qʝ���rLO>3�QĦ�Q����]BS�T�/���}���he���Y�Ԯ$���b�[�b?�5Y>vI"�6#q��U�!��UX�di�|��z�	���"��䬳6�%{�\�+����MR���r�I��a���+��,���4T����r���jY22-4���m�n��#��4Lց4��0P��>�Gt 뇡�n0qK,Fz�H7�%�	�����v`�#����mӊ���F��|~���|��V3+��d։���Ru	��u�U@f)6�@�ʞ��ݱ�~|�!ˈ�c1[���Ĥ���������/Y�z��2�`�W\��F���R����~�Ҵ�+�a��(�+���D�
Y��d2�$:�Nk=��R*Gͬ���P\�SؗF+�J,!
���ޡ������TQ ���	͖�c�^0,U~�7{(8Jy2�զ��8{ �X����8�u�q�S���%�Q�� ��]d������P���c�������:~@ǯ\-�0��G����^{1	��$v��I*]NxQ�����V:rݖ���I�0m?�� ����Ӻ�Z9�i&bm�F)-��0���M=�y��l.���p)E�����IsR��>�߾�Qv^I�=�*W��4������)�S�yTPsHv*U�?�T,��#�mG��3{2z�\�F�rj���)�}�����5|y~+Fz�a!FQ){W�;��a��m/�r �7>FLZ2+���6�צo�ݥ�,|���'�ќJ��Zn0�iz��ߢ�t>^�sV7�&x�P@��}�@�ueE�H��r��oc�n�'�n+��f�D��q�$������|c޻0��`_��I�R�vl��⦀�r���H3�_|/��k�"BN=���[-��ܵ�$�5����a�B(,�ծCqd��q�4Ǭ{�T�_Mp�
z(:�W����(��������[��f$��hW�4/a����,?9�F���S�5���+�����^ĹM��J���.`��T�zV�?Vzש����M�K{�p3���mD�O���U�f�h2~)�z�6cK?�3��K�&����z��`����8�㽗�+E<;a���]�%;�ME�c&�'�b�a4KT�G,5r��XƮ�Ί�3�ѳ��'���33$F�����f��`3W�˷/E^� �����D�f�'�g6;�heëy��;��h-�4�`p���u��[��qWxe�G�sKz��P���|�*��\}���A[ufu�M|`������E�!Xs�K�[�?OmX/�h|��84E:e�9m噫�W�/,�K� S��B( !A,�c��}r.@��̗{�8`<���l��"A)d���� ��-}�u��ܗZm=�{(��:9��ZBX1�R�ά0�^ٜ�w��a��z��v*��=������{*����xv\-�~L��*����#� `V:'�9���7�+[!�ӻ$|g:|Lj+�l�r���"�n�'I�s�R�C�NЍ��X��E�0_����uT�����n$P���!���;zLK����0BՆ�&�bӭ8q
۷�s������3�"���$�7���e��&s6��V]��<�d�|��f�Y�yj�G�GZ�	���W�h��a�0V����K�l}��Cʉ�	z�@��ޥtr:[��?�T�±�ɹ��^P�<.Y��U�q�/[|FM��Hz�Y�^�'y�j��
-��4@��MPcG�M�yݮqw�!�3�p����sS
�L5�T4������O�Y�밃�'��a�یʚ|^3Ѩ�>)hv�}E�0J@%W�ϗif�c�X���RWJ�끃tr�͛l�K�Yp���.R���$�	M"#D��B�-�	���W+��q�O>����1B'!]Y����em!����
ۻJ����!����7��vk�b��S�;��)�du��ݯ��.��x����������o�A`��ƹUh��F
L��*D��&��xb����%�/�L�*X��w{���2�Y��P�vI��|p����E"i�X:���q?�]�ʃwT���$��]$��P*n�φo/�]��*����B��Y>�!���Őa~��A9L6E�Gf�@F��tI=㤠�8u#��]-��K�"��n��!��:I�J>M���Vy!J�q�-�mLʱ�>��-k��8Q#��߹�c��3�h~B��>��
�F���Q������S�Ue`e�B85�ss���B��B�"�KQVO,��*<-�(�E�c<9R	{.����#�n�B��YM�A:��l_4W#�����M�xo�]G��}�5�Oѧ)>#����!��03J����ɢv��)�e�>bG���4�t�t�V���q%RG��C]��+T7&��b��-M%�T��"�x���X����D.x j��q��ը��_���$�?lg^�SY���% Ҍ�Jj��l�5��`�0��ޘk�I���x���!���C<��$��}���#s�
M`�:'J����Jܛ?�8����>ۑ�i�����r�8�c:e 専c�	_��1Ӥ�:c��:d�y���""e��}����=�O}�|��'��3�A��|P��j��%#ǌ�3���,�yF�;c�@�f���?��֪���7�������G��ԁ���5�������rp�Tm��l"�T��s��}=+�;ѱ�������A ���h��i����h������f���+kOO	N��?���x�2xM��d鸲nU6�b�7#:�X����$����f�?����[���m:�ۻ$���k�Q���1ÆeeY�24���� Bc��U2X�����5

sm��!WH����_��Ty�PsZxvePZ{-&�����3M�ͥ�����w�h��.I�Zp�:�8@�O����(1��ډe�}��<�J�l��	�'c��R���P�2`9����fX>��3�-�|yl.�S��Q���0�V<�XF�vSM���\	v�)[�����xS�[s<N.�Ԝ�Vdd[�n]v�yw����d��@W��u�BALu�;/8������9c�A��
�&��K����m(�;�"��
t9�b��:���<d�R�������e��n����rE/vC�s--��̎}�� 1\C��Qfx�FR&� e�G",���?trq22�*'U��� �h�BPO+{�n]�nV�E`�P"�3m��@��*��f���>�,e�K��E�� �������OE�M��͍*����Oi�F�8��0�ѷ�5e�$#?JW�������6[�	t ����Q%67�1�{MZ�zya$�p쒏?\0׮F�u�c�F�`4Kz�U�̻S�w�����u��l��7T�KQŠ���4��@0�&�܋�פ0YTo��F�>%�&���b	��Sn��#h�oj���� L�v-x2ǉ����p��l�\��C�?xo��| �	.V�����w�]7������0��R��/Y/��
L��Cy�:�L�9D�k{�n�G����C_ču(�)1q
��� �Tcf~��`�Zu^�>�9�䨌G6ykV�y՚����E�wB@N_�BH�F�,CZ �_E8k��ڄA82��LZ� �6��ސB� ��œ� `���j
"oT�
�QMn�4�-#��c�x�  F]���n��R��?����G^��ln'�S�R��/���~�9�6d0_w�f<��xA�Zv zNì.w	Y��g. ���D f�42A��E[�MFl�u��]/���R
h 	5l�nO.��]�I��+���4����T�����3}с O�V�����5s�M��ͱ:
k��E>ոmr�ZH���G�aF2���*����=��+�8��O�q���f�W�W=��F6���jS���0���D?�W��z|�����������R
0Od��.;���}�\���5L�&�sZ��@�r+P����U)��s��!6/p">�.�� :D����M@�C���l���3��u�e�>s�ǘrVG��F�+����n�S��r�ĭ�ߍ�Iz��\tͮ�eN��{5a�sa9A�*7 o�0::��	�<����^g�:,��ځu����^Ū�G�HǬ����)�1��wo�ni/���V��!8��r#��"��4���C(eG�|����6�>{V_�j���ܻ��L'UL�����J�'9�R���U�Z�2���IA9��������\�l:�G���J�c���,,��cx��k�g¼󚸶�j�)2�6�(@����{W�s��$�]�H��[����Tr	$�O���d�S����U>1[B�8Y��/y@܋0?�0��t�b�;�����w��uIpw����ֻ���̣u7,�'/���;IƓ��r�ᗔYd�*�fE�o�kK�Y�e�1�z:L��U6�v�d�:� �-?��L��m�5�l�ʠ{��x�/\��hPuc8��/�&��s�PۿR�΄Y-F[G��+MU@3Gg�56���'T�_Vq���X��-������`�)�*�Ӆ�l��h4�p����n!I8E%�j�F��)��zF����ֺ���,��]����W�[`ɦ��U�g��=��������yf�F����(R�?��}�G혊�M9�Ɇ���H�\�,d���ճ|i����Z��)Xk�#W�R�����N�ힱ��i�u��d3��Q���/U.Xm�Wa�&]�u�l �F����,�Q�r�k5Z�yw701��<!�iM�hD��xÞIjJH��#E �9��o�H�,��zc/iY�Q6S��en`���@_�}�0�ts�c�"����Ywp.	m���N/�f��msͶ��0�,@��P�a.��NVW�����X��i(c�|XW�HtgiGC���H< �3��Ó�Y�I��`�m�OB���]�	�̼DR>��O��'�J�O3V�@�W�͗���t7���O�N�mK�S�� ��
Hjʹ�������h����D�>���,!y;!�.�l0���~G��4�a�;N�gÖ���s�:T��2$2��ִ�@%��=y6�.�C��&� //L[�<P�H�]3�O�g��,B=�'�|w}.M��u��Q�vb��1��HK��VF����X,��m��F�'�Xk�o|C������T����X��T�b끿���'��8�7�$���㧉���bv���E���uvh�/��
�/�q�s>*��5sB6��R�B�����e֡��AD�*mI�lI@���z"�R��(A��pZ����0WflX�Gt��+���T��;���+E�ß&��-���w�g�Ťe�4�$�'���|�E�D�XC;�_v��,���k�SA�)�9������oYw �X��&+�n/@�;ۧi	��b��N��3r-�c�|�m���\����o�h�:� �ݞyUx���Z�@^�%�۫�wՅ����ڐ�{҅�l���J�dl�Z��Wy�{��{I�+�gμr�i��'�V�\&C�P�g=�#����Q5��4=�Z��lO��9'6Yr���n�Ժ"����=p���jkP�?�8�bzh�ET[�L������L��_���f�x`iE��V����J��Q����A�_^&��]q%����y�W�Iqk4HOhU#��y̛��:��Ҧ�&�i6�>pI���I2��N��K�7�v$�	�:����<R˶
h�ʀ,L��8��,:�7F/���{R3Wԥ������ʍ�I�ǜ�W�]乨d>�{UY���?;�o���b�w\p9�G���@�D������-�r#ة��e�W+`�;R�V��
-4(�@+��Z	��YXo��CA�������|�O
�Yc?��b�z};$��V��K��߷H�b-F���O��%�ɥ����U���й���ڶ����ȏ�5t*�
Tw:�NRH�������J��ѼR6��^4�!ݒ�̸3��\E�J��6���TcJd�� A�{o:]/���V��"��;�l�=K��iYK��b2�!y���_���,��ԩ|��1�-��rlX��Do�F�m�8(���8���rZ}�����O�z$
2R��̅[w�Qz�d�����Jp��W��V_���.8n���r��*kN���` ܇�a�z8X�MY�{���i��b�?�Xql/Ċ�,���*eB��-�or�?~��,��wփ�R`�HY2�X��$e�̰�(4��!�R'�'�=mfO��vMtK琾��5���֋�@��;��r�J9��#hp�X[�?"͏�݌|����>pR_)�{5v���]!M�G ����L�fqK������	b`��B���]���S��$�x�y��Eh͐�v���|om�%�+�]�Ca��*��\[9_SZ����QNk
�x�q��B����XR������L�R�W���TetO:*�o���>�7$�?�����bI9�T��	�%�I��훱�βt�"�$=CBI�n"�'��	*>�o�5r;K�#he��Y��bV�=�a�x�(5�x���	������Vr� �M�yK� �n��:B�G�]�����$�\5�Y�sfr��H����q)����h�F"���,�rf�6��)��k�R���Cb�����pa�J��$�(��II��n|��,�8�Hy���$�N�K�oU=TJ�9�>�X��R���c��?�&u�M����0�a0.z����e��
�5H=�\[-mf�w8dC^]� �UQn�`M �6Ӥ��A�5b���,	���@I9g��1�^�ng��I��̛��{�&�y��%	�r���I.PN{%ާo�[�KQ�Љ䒃,e�V�)VV�7&x�OTQ?�D�q�9�A�X�OnƎ ���5̴I�n��<8��f̛n��шA�#&�3)�T)O���C~c�P��E�l�J#\����C�%�tQ�4D�����ثzW�����P[�G˹!�e9]W5����H�Z&P��^�9��0�����g�f��*$�aG�@Dc���=��^��@�j��_f]�g��� 2�FN�V��?n�x���{f�bTy42&���@XHʰ�x�� ���V��)dw��_ߺ7A�_fp��M�Y�'�&7Zb�?T�1�w3ڨ^:G=�gr�a1���Z��_-���Т��b�����y��)�kݺ2N�E�0���_b�F��?Ҫ�x*������Q�=�6e&rl���s����Km���5�*�����\�Vk57'23h�s��m�X��"���"�'���%[Lѷyk`W�2Y޿η'����[��i�ϗ�N��7�'���V�����z�K�/�G����I��nGª����M��H��J���{��Tɧz�|ճ���L+"��R` P*�s�#f�&��T:)F9�\�4���S�X�)3òԧzJ����`��[�^<���F��S��j�i�M�0���'�)���bEh�%�i�Aa�u
*�E�D��o�Gas�$��r*W/U��ɣ,*�:)��Ө�2��F֍�׽9��ϒ)_=_$ų�F��S��W� <�.��f����9syP`��V�yYR~�Y��H�2���x7+)Q��_��\����&��2|�+ݨ#�[��ą-6g��D��>+j��{�g�|�)J��L"�*��9��m�랥�%y!�S���ք��}o��#|�N�ɚ���Lˣ�_>>X��=-�E&��!c�(]a<�pRa79���Y�ۭ�n�U�^O�R�3��}��}�x�;��~��e^y���w���zH`!E+lm��^� �[����9�a��hh�aJȜU���E��R+���Z@7�$��1��{C��=#MK�[�����@��IlQ��xPAoXGh����}�|�1U]X3�,7��<]^����)G+x9\���᪫�3��S{��L�+��:�{��9��eP�h�8`���,�����XH�T�0ֈ��"K�|�|�0���z��i ڍ��9�y���l�
WI;��E�ˏ�TXe��U�*��Q�Ճ{R{T�o6��"�I��:PpRd�v��:�Jk� �����j��FǨ��o��Z�!�wa91��?8��>!�U8=���ɛ��܅t� ���q�����즇�SG.D�A�	1������MJ��:�ഛܠ&���S�����(��'T�E��1�l.��^�����A�z�������!�1�-Ь��mS�+9�Um#}���?E�g�6�;+O'8��j���1^���	';�/ǋ���r��!S�w]ߋ1�n���+\�|�i[IWА�Z��@����ȩ`�h&?�JҎ�>��aʈ|p03%҉��G�{�kJj`5��^�{��:���<����R�`����"<�k��]�6At�wR#[� ��Ιy7������@}[�)��uN����k�)����#'*(qk�S��@-��A���0"a*]�IU��Ӂ:%%��F'΋�"�}���Mx>CJ��V��0 ;Ow�X\^�ۡ��i�d����D�ͱ̓������a�'�*9q>�]���ݫ��b.���&�YW�e�韝�_	�NrU7���o/�϶o���a��,}f���6.G�D�Ƹʅ�}Ru���+�I뇍Q����Ɛ��x�Ql������'��Fr����}h��mA�v��2�&�OND��(��h��^�.f/M؆ٙdQx�b��I�"�6���V�Z�6Ox�WM��~����N�7�����tE`��.�Y����� �D`(\�V�vP��9�m��焛��뱡L5u�6��_觨�X9��&J���P�Tߣ+��z�y�8zX<��k'�)-(s��C�4g-��qy��u����u�lӖ���h��lbLL'Rn�˽����Wy[��JR3e���^���k�a��� �"6�(ەJY�(��Z�]�Ei;��Д���A��通��W4)����u�k���=@�������Tgf�fr����_��r��@�;�Y��Q�d�(z ����'������b��6�t^���=^�1��~;���%/4�^�"\B6�5@�t�}d�:��h��R�_S-$�O ��A Z�7b�����Ƣ�jL.۵���s�`AIU�8r���'��k�L���:9����bs
�"��2ѻL�b/�J4X7.!]ٕo��'~��*l���2D�G��g�K۴/*n'�k�B=�	``H��q xKi"��z��&SJd�0r��&ƀδ��"���{5]������f;�VJؓ5v@SE��-��|Dh-����]�+�m7� *�R���L���aq��{��I�販�Q,�wm?]�N�'��*HQPO���,�Gp��ąjٯ��
����O���g�@��_��Q�d�&qԑ+S�d�eBإ�6�V_v^��qg������n��|��l�X%�WjZ�:��ۄC�;	�S�!������JR����z�患,S���Gw$�/��AsuCY�Je��A��|;�Y�gps3�q��ɵ�F��Df��-�zƹt���\|i��Ҋ��!u�`T��t$.�9����+�f��umy�"6�O��{�̿m[���67�C�Nv��s�� Y�+{3~QV3�ĸf��מ!%�"�`e�͗
�lx�a�T}E�\���O���àj�%U[�VZ���w:��qKy���Fh��w��� �m�\J��-���K �q+�H{cE����T	���,���)d���@�����,�|14uvrG��	$��U9.7^b�{���&yoX�OY���'n���B�Y�����I��?*΋0`�9Hjt��v�<�������_���_����Unǯ�FW\�D��G��ī�Y�����yn�DF2~��/O��\O�9Ȏ4�;P��z���&��kr�=���w	a(���;����nh ������ǪI�hi� %�U��M�k�
��恃n��li'*���'��X&&gr�:t>N����pR��Dc�Ѵ����,=����Hv����[��#{&�8�Fp��GA����0�V}B&ƅ;�
���y�r����<�"ǆ�9tՀ�4S7���D�����U(�I���_#�A��u���%�fh7!�H�l<G���dv.����t�Ώ7����{k��|�5��h����#i3�`5����JA�31�xV�]����t�q�j�V
u��Q�:�tc���Y�e�⻵/cp�=r��4x Z�r-��M��*��VI����*�]�̉�pv�Y�AQ,H:�5�S6�+�A2W�F�hh��/�8Z��T��'D�d�ݼ��*�E�sR�&_��@���b'�M���H�&��.r|�I�KO����-�`�}[i|��t�&����у�P��)�7+d�2Pho���bԋ�8}�I����Sa�G�wn�G$Q�g��7��B"�^+UO��#*��c�;��M��囲o��]�FQ��b�&A��&�R�u��ix�Z���dk�]�N,�C(�U��%�jbĿc*�J��ċk$G��'ȴ�:�����)�Ir��I�h�#^x"C��j�[դ�Բ�!�,Ԣ��b4���&�n/���� �Z]}���}-�_7@#�d�@ųv����9����q�`�!���H��/FՖ�H$�Ц����4!��)��p� <{�`��Y4��-�����Qt����(4Ur��Շ��83�G)fkA�����+�hN^�xcO�٨�$��)�#t;4��m�!╼��tR�Lo �ڑ�n��܁�z��?���g�x�k�:~hɬ-	 ��?+qze��Ώi��=���[T`�
%��]vS��gv��I��<���#_�l	PhA��Eq��}F@��Q�N��V;&�{[y+�Kl��:��8|�1������B�[Y�3f]7J$�;��Mw�:�٪�����T���¾���J�m�.�$jn��XEu܇�j�Q`V���n�qg]K��/ST7��+�<�,��U��
y�S�k��X�P����d_��w_g��Y+.DQ�ꔿW�@�6�J\|���;���s��`�Fl���C� e܂��B�S���`���&_��� H�6i��F��0XH�L�5#�L��,�y�,��X'�)���Z^`��h s������mչ�@�8��"x��H�e�B��r<ľi���E�M��n5$���{={/�r�QT�|'� d��U#r)b-v����B���͘VVSm�t�x�_��o���7c�Y�l�g�y}֝�)&ª�
�@�B�w��-C�������O�f�����#V�8�!~q���=^�8�"���̵;	�rԴ��-WRVp��[ڰ��Z�-��a��E|~�w$�בvsZ�1W��d�+M��ȶ�ܔi�;�:R��a5��|E���k�˵a��*�Cҭ�RH��Ǝc���Ԓ]���@CgӢ3�|X��p��A�U��9,*x��t�&���Xx�� @�t�������K��a�>=�4i��h�\�_�#�m×�@�'��F:���z�sU�I�ϛ�lJo/���d�mp��?���Z<;<�� }���ȷLs��ds�����r����w��|_�����P`�q{����(��9�`>iI�?S�q_���v�:�Äm!�`v��4	�"r��/���N�Bn�aP0����j�Ӏ���*-	اc.i�Ք�� 9�T����@k��V��7�0���jM���h{���{\"��*��ZQȢ�Aяl� |O�-S�Q�ȍi}�N�馇R�2MdC�N���k�-�ºnGF�f�P ���h���!���{D��=ݠ2+6C�PZ��ay4�"�'A|��F�G�_�"�9k;�9?�]`�N�vTҗ����A��G�Q��aK,����9�,��SV#�z����M0�ԀA1�!|�y!�k^���ڄ;BȄ�-k�9m9w,�V�o�:�W�X���|&�����Y;��Kw SZTa"(��G0\@X�%)�J�mA����;}/�V��/ߔX�}�gA��O	W^�����%�v�,f��GC脊�4n�g���~u�T4��UT�p�t;���j��{f}Y ��=;�]��6)]R���[u	��?��R&.�aK��4�96�qv�������GS��򡫂��&�%[3��~�����¨���k�V��]��>����D��$#��ž�\#�f��J]��k��rWG�Z)��� Q G�;
x�O��4�vH��+Jb�JL�×�]�NpeW�h<(�%f;<lC�EE�"��x�(u�z�+U�g�������̘ه_;�?P�sT%�#����k�CG�\a�N��^�m��@.?(VO��vj�(�FTsx���k�R�8����Ҷ�j6bu�d4��+�k�0�Y�Djl�}V��^��%��QN1<���Xye��7�,��B������F~��ɒ�H:a*]�\[8�)%>62��{�0�:*@�j���w����p%fu�W�*E�p�	�8u?T�FH����KS8���d�6�C:kc��6<�C00i��c�ԩ����Ib$�$�鯶��'��;"����r{���K�%=X�-@b#�3zٴAp&p����}k�K�K�[��Oq&�>�������\��]����6,}������f� ���mü)`(�������S��c�C�V���VL܍�ݪGVӤ��.���ʘ�jE���i��Hf)t.n�?F��h�Ff2�^�yk��+��xI�N?t���y�6�(Ɓ&�����s��/���W�
4�R�_�s1�wmֱUX����y�OP��M`�9
s4���ۼ���!�o?G���m�����C�V+�~ol�8�o���ݼ�����g��,�&���2B�����7w��rt�sK�W⫏w��Zv>?X��L�v��,&�����n7C*�#su�'��-1�#s<{?�,}6\$䮛+:z����ـh=�<�D�ff�y(+��q�؍ö��X|���K�2�Z� ���䷦���:�'���Dw����{E�0��$�T�F���8�I����vKv 6���o�?���͙�]+�U�B6��M�*��^�6�F�����:��u������X������lkR�iR�퀾�A(2,���k�N���]!�}"ń�=|~�O��ؿ�g�`S^�\��^��1��<��uL(!�'���ț���G�te4G��+�^ū�^�:��@��*fs�eq��0`�� �}+W}��Y;C՚C���t.��� hQ�a��'<��0�UBy�]��p[�� %���Mڒ�zFx+��4j������h��R-ݶ��mY�Y*b�iP�N?�4�'E���|���P/�BG��gS%��ϛi��Y�$�qmL�h�
`t�����{�Gb�����
Un�5ڇ��\d�>�\��cOX��P�:������S����d��1��7Oui�����MA0��Ѧ .l_`���.0r)���0'�V���k����14���<�i3
��׳ױ�$_�+'���Oz��F�ڀ��d����Fލ#[��(h�� LѲ�cY�"�s��Hz���NT�uQ��tj(�0�s�!d��T|m�3�����P��Za��tq@�/�������y���`/_���T�*����L`6�m����!��lX%��!�FU�p|h�~����~TD��c�a�����(��B>wlE�W��c�@˔,�������0�~��K���ZA.��׽%߉�km��?������%������L�諠*�!W������z	BN=��/�(E�۸6j�A�C��qZ�:Ų�c���3�_֘4�a�gI��%�ܠ����"���Cw��;
�٘��
�l5�A_�g�������~���g0�I�<:0��|����<D�	���#�w������=*0���RE
���o6Յ���1����bI�kR�:u�����ld��,R�v��6�Wl��S��w͑�� ����x/�M�JH��M�*�F騁�o��H� �:���̞���[v��SG���?PT��+���)�ס{@�E�X��qK[s��Q�<R��o�"�.3_dc�0b�z��.+�
�ƹ~�@d��[
�ϡ)���o�/eҰ! �W!l�����|~}kR?��H}�}�)H�y�{�80��˝r=���V;۞1�x�.���E�w��S�L��Rn}�����Kfa i�GC���<����%�n i���%ڒ�R��ɼ�'��FбGJCA�R�n�� ��]P3��l�X�쪓��AY��;f:�k,w�A��/��jk� �.8������%�`; �D��|;q�'� s�A ��V#�
���?����hW��=g�7K�9Sg�K&��O4����%@}�v�/3�RdƂ_�la���H�(0��\�"?�O�k)���he�R��C��5?=�G�No�	��ę� �;�:�P�9F_q�ז�Iz�8z>�(�6�n�ŌEb����ۿ�j��S܃8��!F9��E�(�ZTan�H=<q��V�P�U�Q�֌��Wޯ~�-�܇x�0�|`E�b�"p��*������)Ǿ�8mu�\bI^����(+���x&�t����d�I��;�٦�rs��b�Q�>��_��kU��"3�w�ޖ<	�l���fWv��Zgy'�;n���XD���<Mջ�
������Nqr�E9�>�0{�q�M����7��k7��f�G���Jи^O�G;�����#�i�'��f�ܮ�P�`�$�M�N�V��	��{Q�Ҳ������ˇK�o1bn�iĂpC�h:��u͜ۉE�48y6�	�L�	�c����z5z�Dj-��u�O��E���H}�c46}K�N2,#e�b�ǣ����̆�:��?m�j�l���C�E?3���f����^�BbN�!�T����V ��J�iL5q0~r��At�k�7�*���MT�F��L�/�ԛ�F����^��n��$
�`" �0N�OJ�0��=��{N�"0��i�#�<w���D͋]���#�!�Hc7@�rXے�Cg�_؏����T.��c�G�Ūj9(9��N)���HXg�����ZR��y�����}��a ��&�R��� ^�&ŷ�.L~rӘ��+�j�S."���2K]7kjp���$�_�
wTq,_h��L�;XGK(�?Fń���Z��X��� �V�&ȭ,����L��&<����mO�z`�5�&^�4�qm氵@||;N�ǼQ��/�4@MzZ��Tϧ���]^q�Kۼ�d����U�r>+�Dx�W�K�v���~���*U��<���{��/�\�<��ئ:��������M`��$�?[g��ڙ��Y(/}�I("�$GL������=,��4L\��m�B��	�}gi�\"�%8PPVJ��>#�r��T~j�_����6L�W�'�(���Y.s���f��u��Y(t�gBDu� ��;V$,�8���_�yej7�|���dm�Գ��/t�i�/��;�r�.�~�X��mL˔j� *�Pwo`}�G�t�?f�KU��)v0�I=�Q蒽%��J�_���j�nѱ�AI��r�~�R�x<��f��%��t�O2���l�4#��H��B�׹�'Om�v+�#/&�jH�@�Z�8��C�C�J�7��fz�j��E�D:��n����$A�<Ӯ$C.�1����>\������C
/�+5'_�#%4���ej% �����B���(rњ��]�N�x��=��6H�!�Ⱥ��Ȅ�)����Q)��8�h��N�Q��hV��?NM���*@'!2
K@��`匐ࠒO���(����|#=�}^����n�v�����1�n���VVD��kc
r[%�Q!�6�iF�� ��.pō�U��be;�ʭ����Q,�ݣ�w�}��%�tl�X����n%��>	I�x6/̙����#3mu�սTXDa�Xm��<P���Ntt���m���x**��!�&k�N#�	���p��K_
�E�,���	[������bC(�{<�Ȳ���9�(��e�*��B�]����H��
�ur$��J>Pzj�g��������r7�����j@�N��)��?.}�x輎E/53��1�%[V�[+�r��%��\%R�Y���Tt!�$�s�n�͗�+sc3ު��3�t6�D�2�H���ç��,�yM�<>��s��#��o!9^S|U@H�������p߆�K7b������ע�MvZ��AJq,݋E�n���*
�����L}D$V@���KA�rr���\|jX�p�L�*�E_����2|��i
t
�h�p���/���� :܇K]�� ��;����%�T^�V:�y��o>q)�>圫��D_qo�>vq���=`a}	h�j�
����T��鲕p�]�һ�9��
5�C�8f�&��� 3X��y��'���A�{�V�Wpl�� 9H�tC�kbc�E�P�{�;��[�l3�yD�O)��ڌ���	~6�i�+147�e���ϔ5;������	�3�?a;|%�_�B��W[��臾�@��5mcm��]���Gn��F��H�MK����;�`���]�B-��Nd��|��<y�OPW�|@�G�3�ʿg�>���:�%Z���a�ɰM~��mW�%w��3��)VA|V|/k�މJ#�}L� ��,ju�Ļ���XJ���+��aڅ��'�q5.
�`/��P��V���{1�����K���T	���W>N���6�3�#m]nmf_tJ
�\�����Л��-WLV��;��JU�����'"����V�fE�'�/˿�&e|�'G9�p�=�p�Ŀ��}/M��]e@|�/����U��[b�G�ڿ)$苞6��`����:O|S�����Z�YG��t�&a��8�OH�v��t�H�K� �Ê٣�̴�tǓNo��/i�4'�&�Hi��"�!N
����&����>�1���"�!��W��M�QQ��ec�'_����d���X�GYt�D���:��( �jN�D?��G8�;��ju�������= ��ǜW$vF�M9l+��pT��ONE�+�����CVe<C��1K�Iw����k5>��L��o��r�p���R>s�Hsm'�%lIvv+�[dh���e̍��[���݀���� $_�2�qz�C�J��ٽꄣ�L\ >�v'I��hE�����_&���Z��4kQ<m��,��3��TRu��^�/�&�e�A;Hᚠ)���1�'��A"�$lk��
���>8�	Ap|��xp!�ʉ��nŏc+@�Ӗzև3���*�4�����p
�w���FPDi�RO�R��f���%n��b�2v�q��TZk�ښG<����(h�\��`��<2���5�sHڲ{��on��7��z�LT��hj��ɝ�s�b��g��SYRq�s%�x���Y[F��?��S��?qv�W�1%��G[=��Wt�L�e�r��j��L1]T����UUt4v��ӌ�ZRh%��D��?�g�Q�����5K�-q[�Gh�`��y���y����&���맫v���^��h��� I�3�6��'Z�h
 L���i7��Ww���#�@��)�?��>��S����L�[�$<��*U)t�e)���o�6��=1�:/�Z�yB"E�I��K�N�'I�d>;��=P����q"���vL�ě]�<����۲6B����Q(��"
�J�=�:*�C���3Z�^��2ҧ����%�&� ������?����	i�qQ� �!^D�ٝ*�v�H��� a�L������-y�'5_���_����~D:�����S9h�&�(kDWEvb �����
k�{nCz�V`Bt�����e��� ��)*��[e�F��D
��v�'-�C�-njݻf�6eM�E}���S�N���S�,�v^Ą>.4���2��@j:�g�A˛��F�qq..�� 8��O�vJ�FN���!Mq���O2�ܘ��b2�8
��V��g����Z7�m��=C��G[�����=٤�P�EE�>�o� ��镬��������텹A�{�=]��7��!�ݗ�ok��.b��A�rY0�[q'��mhv�eYY�����,j���L�{t�����9V	��)��Ԏ���\J�=wķ���gE�s���s]�v�����:�f�m�)5�8��B�-O;m�.<9B-�x�_m��J���oFK/�������Uk~�K�x�!e0pM<M�EtZ�j� �N�V^B�_�n�n�#�܁����f�n��q�v�<�1�͙x��T�T����8��N�m��%�i@#*.�?��j]�E�eJg�qd�AGف/+�u��u�i�����Z4������+j(�3�.�}*��_���E������%��x��|�����r��.�)ʓ��pX�z�嵇����dեp��cM�"��L���]�!~�Y��|�c����J;�迴��3��+���Q̒H|�Q�^�ֺ4�)����:#e����!��_$�¥�=�K�}o&X�Yd�Y �/�3v��	�"�g�5��,).M��ɿIm'�8~�`v���Ȯ�<8Ǉ�A��E;�9�jY`!;wl%?�Z g�	r�����.��f�1b�F�-u��>�(�"���*�\��=�v�*��k��qWЊ����8]Ҹ��Rh�q�D������x�U Z��%����u*�#r���	�lP��C�xl9�pZ��>��3]��Ԡ�J:C�A��^�9��ED�\)>;ʶ5��\��o&v5�s��m(U�֯��Y��]�<�E�Y���ng|X�LWLXվ��Nu�
F����o������G`w�@v�N�Pz�g�}��@O@qt
E�~��qE۸S��Im�-�Q�*t��SkDhO���9{�Z��C?D |�3k0?����NS��b��a�}��� *ii��a�F���AA�yN��c�R7�Qz�cĂ �c}�o
�t[gn� >�Q��#�<H��P�"�:4J%�O8�yܭ���]R�~�I[�'V7

vd��'9�Jg~g�rC��w�(��2�������-�Gu��2�c���irڔ�P�ќ}���ÿj)x�5�H��6���Ϧ�z)5�$���X?�
���^���g����K�
�%RM8���zx�TR�9�����s�+�ɧ���6!�?��$���w{�����l�g@��Q����`��A�[����+yҋ��&#í�����1���T[Dq�&"�j�q��_*:&�h�<�;��G����#;ﾻ1d�'�"�bߪ0�^� b���%r(t���<"d�� ��g4�±�x�a��~�t��Ze1�}VO\
���h���'����!��?0,D�Q�e�����K��܅���s�	��=a�AK��m�fy�!��M�.
�E|[�����'��m�!;��=��������T^~�F�m&��(��SLl��{�Ȯ��:�lYX=��z"M_)�n0I�����ϼ�z=h���|� �\a_���v�͛�+ӹL+�%�Tf
@�,�m��U��)�~��3�V���48x7$�\�G��8"Ϝd��˓�G���a����D�5J#ԏ�y�Ċ8�a���$���@�ze ��Ή�v�	q�c�3�c:�]05_��$��d^�9A.����Zhkux8�ܟ%���8W�F�Gw�x����M��'�Z�Ip���&"!�r�-���}����(���XǫdS�����gԷ�������9A�Q�S1
�^�Cy�R�7b8�P�T0x 05�V�g�s�A�(��<��y�m;�t�=��G����*�R89�1��-3�X�r�+�@�AOAc���9��YS��O���/�P�!ҰnA�c�H��FUa�E_��=;\5�o[֑��*���D|]�]�Yb��9�JӀaP��ٹ�5��4L�|O�{dR��3��+M���o[�;>oO�Gm1��B4K#G�$������h0�&���=9�ޤ͇F�!%t�'�-=���r�t�zx�wWV�
8�j�M.��<�� ��=ij)��KO�9~$h���B'ή7�ݍF����=��X'0QT^W�=	uL��$TG�Ҫ��mh��P�yo7u)'�"����Zd��ﺎ�8�^*��߸�1;�4GRӭhz�a���vm:�(��k��r����C%a��
���돮�x4L*�o5�?����m�]	��aQ!?�� ca�̉y9��҄/�f��Qj{�vNn� Vh�k�8uH�E;8�q��(P�c�P����O	qP�U�(SE��㆒�h׹�p��L��x�F@�Xy�}��;#�>a��s���F�mG�46W�ث�}kX��������$�a�_�H.,�|�;���$u��"�����S� �T�d�և#0ԯ��H�q�;�[���zǞ��|p�VA-l#�6��r���Ga�X��.�{�qt��cф}�xx3 �3� &���y��Ȍ?I'?�k��v
#�ŵ)��(�g�]cSa�/ro��_��.W:������ҙ��;�����6�dA�N�k���ؠ_^�?xbS�Ni��H�Q�e�w�T��l��\=pᨉ�{w�~���E;��ݘ<F�Oa.S�����O� ��l��H�}�d�������6SRD!V��-={p����Gq ��~Cf}���'R�s���cλ����\�s��=�gtj�^�bx��82r��	�⦪ ~�Nn.g��'M*��@�w{s�J����JZ5�n��{�����Rz��ظ�9 �)%	���鈄J�(��Ef�	g�x�����?��׀���2��d.��ƗLG�N���_��u'̛]vlBR |Q<�� /��������R=L�;@q`kG��+"��9�3q�7X�C~��.���D�^v@�˵��~d�w>���r%B[�~J�5(1>ta�+t��{��mgx����_�=v0G�-��/��٤�VF��q �x�0���"� W����i�[#������[�>�`�4��~�́���v��R��Up��G.�L�u�@J]�������m��^�	�mK�f���}��Ҥ0���ua���\A��Dkq��
��$�p��4��
���@�p��ķ�7ǌ*�yj�����v�����H.�-�od�����{����2�ɥ���8�Y�]oC/���"��t��0������,����NP�Ů���ͬQ(��n��ۦS��Mi�{Yr�������J�_�8p�YTE@O�����Y�7���b���v}�>)��w�� �*����D��䏏�3r�'���Q���L<��� Q�} �!�7	���T�N���w����]j~{�l�B�<��2C�nI*pB��\�Ne|�+�lz�[!X�%�d��T^d�/���$��H���]5YM�8ڵ^D����"�	��Oy$i��p�Z�/�� n��Q�xr��)?����\���#�3�9xL��^�����"��(���K�q���1���D���x뢋�h���CR�?�҉;(~�l��c�s7�����qc�L��'�ܠR��(�����%��Ļ[�������;Q�q���c�����}�Dqr@��_K�	�*}��T� jI�!c����z��;�%]A�-�>*�1��HL��rZ��R���J�E)k	:J*��bs؊��zi�PK��{�I�q�`��Fn��0�pC�;�������~A���BOh�uŸ�m��viz���bzk|3�L��`�c���� ��C}6�H��7�������]�dg�g T}�I�xv*X�/�z�;(������a17�Ѱ�l�^��z�pq�F,�(H��l3R�<l���cY�>�13����k��&��N59*n�c5���|�f!�8��2�,5'���!�5�$�P�y_�Ƃ�_t\,�*���f��t���j=�.�υu#�!ɍ[��M�wI�t�
�������S��}�>��ؿCSs\��4�H�kh6��Z(�ySn:v���s�*7���y�`�_!�1�զ�Q�Zrj!lfI�>��3��s���d9�����������@���� 2>d�x�+���IK@��Av�����>�;�HÍH!7�
���y�MI�Rw�t��݅�8k]IɄ�58Q��AKK�����犥��q%!�������K�Ѯ��f-v��[��¢K�
A7��:����{X�H��/�L4�:�s�4�HGZ��������XY4i��ү8��݇�1����D��:'(����YÂOK���w���W٬���V�2�ο�~�%�V���]��9[���u�qy1��-�s�%��jt(?�E��j����F������N�b�{���m�C��c�&|��Q�����}�td`mL�s����Gt�զ�~	\���Μ�.|l�Ӄ�o⏈,���̯Y �N���:�y�<��n
�"�CM@�i������U���ǅ
��7��e��A��ߞFƖZ�cl~��C&��t\!䗌��纛���U.�Y�eͨ�gnH?{�"����s���E6�'��]�W�'Z���a�M1t��)�q�����)m�z?��k|���@1�3߀l�B�1������Op �?��A/%��kְI�¾����)�.NU{�;����C�%[M��y��L+;GYX"q~:;�W�7*��g�ъ�m+��"�9wj3��=0r�!���ɪ�����$������b6�[
�%>�UM�>W�%5^�;�����g�U�*�n����oz�<j�Ӵ����P �_?�zMӵ�d:V"�ݕ+x����,�E�Z]�'2�^�,%�hE]�oRH��%5��L%m7��$߫ng��r� �V8���,�r�*X��5
	v�Y����ۂ�I6BPVHs'�0�x��,4���H�:���O�_JE?�o(����T?`�2�R�۹�����̸���1
��5�zl���?���M�c��j�)Qhh���ta�����S��M?�=Bj!�x�S�'�m�����h��ΚH�y���p:��E/����C}��2�z�N���m��fS4RU��ؽ�b���qVg�l��ף�ǎ�7q��Һ�3��V�H}��{JD̛z�� }�,�%�kܡA���ͯ)�5|�ϧ��X.s2��O2�LI\v�xK|m�D�k���[<Ŝ���.M����"��/�Wn^C�Q�T�&x5[�B�X��p���24��K��T��9��e�,	Kt~{_�{(�9-�r����fKĿX���Mms���KA�����J�a�%�Z�G
T�����j�ia�(�d��H�s�Ѳ�ݚ���Lkv4��|ӎ��#:���CBME=P�"�m1�@U]���*/����ИL�\����#�߆���D�._�v�F��87�Z+v`�8�@`F�%W�U��F8&��M+l��C /N_U���W؏|r��;����LBf�є��t;ؙ�I��d����[P)� ����~��	y9yA��xh�H&U��5��2�:��XtTކ�HKm����U�~�F���y�M��4���s�>˹k�Xχ�F�Z�Y ����^��2��q��Qw�6��3��
��8��(5��_��Tx�D�1}�Pt�g6P�7� o
�p�=ja@.��7_�h)��򓠏�������C�}�c[�GwaP�Ls��/oTn�Q���_b�ŖTz��C�Y�&�d�����q�C�����%�\��a�B^c���GV3�USvؙ���eR'{#���@#��)�Q����{��������H��-�7�#7�s��(u���ᄉ>���b��� ���by�֣��Aȋ�RU�xP/{0c\�)w�!��+N �c8�yP��=�����Dz��D�/�s�|�
,mϱ���\�.�ɿ�=S�"B(��&�\��n��1˲�Ǯ���������j��Ж���*�GS)�2$A��;89�V]�0Il�:�d"h�k�TJ���tcx�BHt���4J�"�%����ț����=b��\���u�ITwԋ����9�x}s��3�z_�;�Sv�'Ed��&�`,����6��\re{�t��0�lٽ��i��_�-�|�"��z@�7�Ҹ�G���RPNU�cA��Tg�fD�V: S�2�0�O�gx���+Z��i�ן��B��Sٱq{a����|9^�^
�SO�Sw��Z�� ��ӟq*�E�Y&/��u�f�A>�qw��]�׈�U�c�,�ahjc�h����0�p�2����F@P]R��5�P���~A�$/�^��brA�5
�bǰ!ە񄵶.��w�{��s�'b�vg�"	Fk�6x_V0GS`f"�nhԗ���E�HL�RVjT�����l����\�n��`6�F��#��`�S��(��*���2 Qb��(4�%��-(���魴i#�$��Ȭ7�F��|� ��S��J�![�GY���(�����DQ^؇���bU���c���_����������eDii��D��f��XKE�
T�j�Z�x�KZ��� ��)���{�;i�9LQ[nI&���e$�x�U\-��;)�⢝a[������������?���Gv?��X��)�t4�ES?S�[>�HS�[����]V�\.�yr]�B��{]�C%U���
�1lBq����Ig��m`���:v�t��2�!=�\�]��3Y��.��p�]�hd�8
3�]�O���`K��@"�]j`u��flc�ӿ�+�����v{:�C�,�Y �orl1�{��?�6�'�uh���B
(o^ϓGw���v�T�Qmg�Y��s�����b��EQ1Co3:��7��H��nR�������Gk �����?�~PH 5����	�VnNr�;����r��s�ae�k�GH��]�:����r����h1��m=ݺ)��
�[+�:	H�
I�6�<gI'��1��l���N�^$ɾH���^#�XhܚB%�f,�ռ�x0��q�U�c���Z��Y� Ի/�X�^�q������&����$��uj|Og�z��/���JA���%�ث�"5D�,V)}]����������q��#J���{����n����d��1��흳��	�}�.f��a��*�^��w�CA?m �8�P�U�&�L��?D�w���{U�6��������G�ܲ�1���o_R�o�NH�4,���Y��Y�x<�a�� v�O ��Kp��!G1��U_=+�Z�G��=�ߒo�M=�2�A#� ��շS ZqY`��u'YR��dU0�<�b#nS�@���&G��۠O_=WLX���:	�� [[$L�Ie}�����wXg�\j�W�Ikc!@UHv^�G��8�˩��BW�^E��ܐn�H���zy��*�p�ޫeSj���5܏3i��z���W��cn;}��ӊR��Z�p�@�*h1���gkժ�i��Qc�q.Q:d�:9�#�~/K�^�q�jh&6�ۜp�db�r?�j�j�i�D�T�Cǿ��OQ�����0�� v���RUu�%��L�K��\\.{̏�+�]��$��!�S����C�	tkgxR�<)��aE����H�B}�+�|0�R{8�{=�
a&K�X}�8Y_��%�ۘrTnֲn�6J~�� S>_՛°�����T���/z����j�қv�;pOd�
c�׳\�ZYPA~�$q�qj7��\�E�XC*X^�U���^�w�s����l=�b;�f��͉���)g�_rj��Y�F<�B�^��NZhA�^���4�������%�蕝,q�:7�f�z�~$��o4�xq�Z�NH������AK���ȏ�3hX�#C[�),,g@�ĂnVm3�=��hy�Jm�q)�������#����d�(UZE�K٘/.ŃN�#�z /Gt�i�\#=�SY~��K�k�ɀ!Vá"�:ݒ��&��L�<h���ݯ^B��G��r�W/Qu���"�|�ro���W������#�@t��Yx����Ov'��[u�qyݪ���?3l��i�l�GA��y��1g��z�qFm�ϸ�;���B�1;���T��}[̾ږ�;�;Y2IL��p�W^� (u/���j���h���5��jr�,�X�>T���Fg`R2J8&d>�4�״���n&� �����PC�I�nE0��H�J�Z8��>w�^���H��C�G��\�wty��a�hzU���I����]H+�ASU-j�̡��@>��EfU��DͿ��`����?��6W۸sž���È��Z�q�W ~@V(x�矑v"� �]�%�>�&;�t�����\Pޅ��e���
�}�Q�|䒧 ���,y�D���>ہ��'�`:�(������)~�b�=�����YØ�^����P���bw���~�����E�ٔ��ks���?׏2.c0{��GZm8����w�c+���-: �vԇf��p�0=�|Za4X����'�J!�?�p�51�����8�p"=ju�C��Twu֥�FV�n���j��i]v���_j�&�}Q�:}����(.OƩu`H�i��a^�:E5�(4�d遥ED6��:��&��
w;K�m~�� �����U�)<<�ڻD�p�\acV)��s 5�a�,P��8�S�R���K��wP٠�\�G?R	�� ,��,=#�.Ί� ���3J}i/[�u��B�e���}
,��-���u���ڿa2��0�+��}�̉�}'g�ok|�g�H5�-�����Ct�t{r��`����Dh�6^3���X�p����S�,���oY�R	t��ɡZ���k����_��F�wp�+a��tdj
��Ó'��#0���|	C���7����N&Κ~H�gk��{Z��*_Om�#����j�xh��XH���'m2�q��oi��Q�<�.��"gQ�v��y�L�6X�F�A&���L@Oʫ��φJ���ٻ/z`́yPC����Xsc��\��ууcK��f�b	'�gn���2��WJ�=2dKN���T���Q�&�8:`�,Ŵ�5y�L{�������{���֣� �֍����_�9	�K�@�����7,e�@8�bɁ�t���35=�������JB~�����t��{�D��.5�~Y�s�#�Z#L����ω͐�3,l��ɤ���� ��n9F����J�5����c�{����Yq@�U�]�}�5N�㦲����ϩ���pnv�,���y�iQ��覞�1!���Rǅe#�D�
�p@�FX��&#�
�W��d�(Jbj̘��[�!I��1�0�Sd�!��4�B�Th�'j��(J�X
7	�{��N�-�0��QZ:����X�\����m��]iO���zQ�s���V��j���C�h��UО1=pJ}�e��j��\�Dp��G�!�2�j��T3����9��bP`�$,bB�ZyL̯�'ǠI6���(B�����$@�p�{$'�����u�K�M��H|�(oҙ
ё6����g0[ȫ�+<�x�Q��&\���G4/2�
��4�~}�;RSz�9'PU�L��N�h ��] ��������[m��s�A#&LAC�M#�πmWO֕^�{hQ�d���dι{���]�[7u磨�,A&���h�P�?�x_ڃ1�]���qh��XQ��<�s�*�]&r�?�϶�l��&4�2���^9�U̕aJARdp�dZB�pp�E��6亸�&�z�K�����>$����Z�:8C��$�&%�?R?J���6uE��z%0v2���dO���� �U� ��.���=��yV��k�7?1:�c*���.���[v�h��>��
�)گş��-�$�D�&/��k!T�߰RP�ͷC���n�u�f���-MYm�����~F���Ke�8K3�M���������f��d	`�aV̷?��uA@X����Щ/�X,��4�n�.P��������N�i���$ �!-���{��3���y8ۮHɖv���2}�Y�OH�{����6��M���lC�bK���"���;���	���|�v��vfx�d&�P�X�DOe�\UQ͗�-�����yKh��-V���sZ��_��+芜� �c/{݅/��=�
��gn�$�f��`�����s�	��fw�J.��^Ҿ�!c�����~����S�A��o�3�׋�;�.���]H ˩��jmx7�6�~#��tMP�2���tf�05^Tw�AFJ����;��տ������3�6`Oxđ�����o;��&�$3+�I-�|_ r)�y'tveb(�P�9���������VΙ7�����x�s �=�jsr��I��Z�D�wY?}	�c�	�p%�B���Yé�"����|���>��4�r�[���lu�?��� J8:���7o2�0�T؁xC����\ԧ�x~�4k�7�O����&q��Jog��ؙ'�$Gb�>����Tz�f^篃aU���4����*��[�t�F��AB��!��t���H�,��bˣV��p�]G�C�ؘsw��s�ֶť�η�9�#uͭ
���
H�@�
{�'�%���T~���9���%|ebƿ~�_���C)�N� v�ao��{����}0o����df!�pV�b/��I����"�90�<Q�eח�h�2)te:憁�?)j�؋8��*>����2�4SHC����l,�J}�³�mi�Xx[�Ms����I�%=�ރ��6_��$i��%m>�u��=�����&�;�sw�m���$���E�Y�~'H��w�:3���Sw�Z����ν4ݹ%��9_R9���;,2˹*-L+���o/���<�1�4[W!�
Q����y����,5�0d5Y����b�(潁5�a"������J�W���Y�wm��l#���b!�t�\�sT"׻�d�: �;y��[�崧�C���\fyV#}'�?�^#��Q'���H����:}�Eu��1h��5��K��2@r8�j-*��j��^�2�9X�^��j��0E�F:��`��C����n���RqS:�M��BrxaG�����>���R�,!�T�w�����[���	5ˡ�=D���n���(Ϸʴga��(a6�_�����&D��)� �OƶA�u`�Y����a���� _Ɏfڱ�0�Xs�d���u]0���$9�1ĥ-M8�J�h�}��~~)Q�����R֯nI�o��h3�SE^�o�l�ڔ ,	�ࢍ�W͛T܉���r�L%?�l;������f���{2�z��~��d�@ER��0�G9��Uē:(�R@流 A����\Jz� i^����b��v�rP�&��^xP���-��vY�."	����ܿ���Վ'^�yZNp��R�D��\�<�u
b�[�_���t�a�B:�rV6D��p��9
9�2���n(��pw�rF��L��,Ŗ���? 5�Lp�[t�F�{���/2��R�	�1�b�U�EBIٵz����b6��Ma�ԣ񥭋;��I�S�Bm�=H�x�{��4ա��5�)��!h��D<���M����Wa��\�GGE���y�$�#44�����/�f�P%���d#(D{y��?�@Eh�S�HI..���Ƚȇ�-5v�w]L-�����\Q�s\�X�[!kX�_��-� �밈�*�'�p�5��)��x9�?Y�|������������$�DJ�'��0�}���Ԓ���vަHs��V��j���y�,�S�o��V)оE�šK��
9%^�w�;9�9�Z��Q�,&�زO$�	󮕈�Y7H�m{Ȟ)L���pL��ޤX94�7�y��Q�F��cJ�Ig� {E��O �.&��V��9"\����\ANȣk�@\�Bl'����Urz�I����FK)rF����k�I����f9ș��2ZƑa+�n[�8[.^b������L!����ҿĩ6dI$�d>�����s�?�!��
����JO#^�ӹծ� ���pN����%��Y7�/��ysT�@o�ɇd��ћ���A�����0�$�_Ҙ�gh�E�"z)(�M���&I1�F��ajB����)�L�p?%�9Y5����KF���q�8?,�\r�tx�B���Ql�_m�B��p�)�bgX���>l��V�PQ����%���э�x�\����Κ�c�	Q���{$N�q�!̼��
�v�כ�l&3Bi�s�Bwi��ݲۡ����8��vO�$q��U{��e>2��3�j�A���{��D{޶%�<��;>O���Ę���L�_�
����)	�u�S���O�5��{�����}�u+��w=�cD�o��Z�c;+1p\_��g��ͳ���o���I�t<��:S������uX�%7�E����d����ǝ��@'�K��� ��]����ю{�2�jj��d��^���.�&��w|��;��z�|̩��.��/�K��tȥ�{�v��ө�ef՜~*����GU=�¡�J�'+�_!�Wp���0L�LNu� 6��|���wG�X�r9C�&�F �/
2� �P��e�fdG������$�@�6�v�թ��ҭx�a�����ǹ�W���z;�Yx=W�{@"t
.YfIlg�V�q �9zp0�F��La�5�ξԉ�ʀ�=L���S��\�03l�\{��'P�<�Ai x+�j�u�2ų�N�<��l���bI����)�Fy�Uwǆ��Ʋ$^���QC�1c����q`��CZ���u}��z�#t�8�&���F�/��D=�g���lS�0R�����R$6�+�Z�:���n��e�ay}^�T�#=s��G�����G�>���[�rW�@�^23`o���H���U%�g��1E�T��bq���̏�`]�E���]����L��L��I͈�_n���@_2�J�6L�F�q����A��f�L��7Fz��������c�75�O�*����K�T�fk�H�w�(�a�w�G0mє��t�m���6�WTf�;[���hG��?Ϛ �O��]A����1,r��J��5���q�#�!o��o�`4�LZ��Q<Ԯ��X��8�6�Q�5�]�qi>&���c�ߣ��u@��W#hx?����%/�7�����j=J���?��r&iz�!��GYf��"~v�	h�.�W����<_m�k��;�3����c�.�)n镑�e!sW.8�m��X��N4|�gɽ6;��haݐ �K2����*�qJ�d�Ӕo���|���QY�����g"E�������d'�]1�+mf}�ڥψ�	-'|�mH����ƚ]7�N��aI��[��%��]uT'��i<��ڼu�/��0��X$�@�W[|ƼDm���&�x�����8"b�&n+	�l.X��9�Ym�S�B�K��h�2��·�ı��s�=�O��!��o�Z	4Y6��i;��5�`$(Ƽ���<��<`R�9W������ơU�A�J�6���S�an�e�M��q�����z�+���	��艹���0ř�b;�B�A���c���t����[F�����<S�(�����z�yw�:���D�H6�>����]���J����	5r��e]-h����8о3�y=0C���-��k՝f���ߑ�wg��V�A.���S[	����0AX3��
�	P�pL�Wii�hpէ!�΃t:Sh>Z�$�~P�K3n�d�]L�lJ�r���dSt�l���);(�:���µjY�d��9!Y��0�����\s����.�?�`���r���;���w#֛����`��j����k�E�|Z~�w�� ��H�N��F�F�������ж�1X�J4�b�aMJ���Sű�v&��=W��������!l�@�iFN���,0������Fk��o�C~�P�NPU��U�ӑ�]�)�ǹd?�J���
�'��,�Q�.�=BZ�@�6�xE�hh�_O�ʹtA ��]?]p��w��
�@��T�I�X?=�x��g�X�3B�I�{`��ƛo��ܸ�!l�(�\�oB7ap�3��f��i�f�0}�E3l�n��Z�
<Xϕk��0���3�&_L�1m��E�|:��,G�`ϼ)�큹��^��C.�U0�Z<S����F�]0�X��l)r��4fA���&` `ˢe
^��S���K>�f��yE���]�~~�+`�'��?��ͫ���R�v�r����;�b��g
&w^&;�lN���5�\P��0��]ÛIx��?�xVa�f��w}�������I��"�5LM�ϤNG�X�(��6>G����ʋ.��U�ú%�ƾ��c抭�K(�?��FwsxAbF���a�|[i�ݑ��H��M��A%�(��|9J�$\)(�������C��ݴ[&�i����I	�R�~tf��c���A����_T�ڧ^��1��8��rud�D�:EYi;I�iô�#�F)�q��h�Hf�L��ss�Fy��U\t~|j(m]6Zx��fa���c�;}��<<{nP���s�J\�����ҥ	ٸ�H'}�FY���s���3%�ps�_��0�1�'y����Y�cU���2}B�W �1mg�� �7Dp��d��b�X��_������h�g����e�cIPzz�DN%5[�<��v
	�I���������c�8x��VK������j'R�Kz��v�M�#�!�*�����
XZh	�%C�������c����g��qOOW�/����A41+h�>���/�[޺.�ۑɘnd������R�)߳G��>�%�t6~ǐkӧ*�1?��b�ȇnB��a�@�N���aU���^�˸��v=�~m�t1�a|7����z�ڱ���t� y����SH	�ʯ��kcW�mt)��&�θ�C �*�@R����k&�i2�g�,���_~]Hی�����,1M����ڑja�Ϭ8�M/���!��J���#��{<~4��c1|�*WY�@1-�P�^���eY���g���I�Ah��O�J���	r��z&#dB�TR������YX�T�"�w(�ܾ3r��ة[�������޷�)�v&Ꮏ��h��L�G�2pu�]vy�/lAs�!'Z�+�j���J�/F?̤�0��l��G^TV� r�6Z.,�ຩ-�I֣�W�(g�ۣ4�2h�W��˩Go��5�� ���l�e�F}J�3���#˚��8��o���3�n��]����`&d�y�Z;�	�������\�Δ*	��=<>��$�~o8�p~�¬3��P��⎚v�ݑ:E�H@����2�Ԣ�|}h������ ��$��r*��|o�p("�zF��f_�qFq��1��!M�Df��LC�r9������j�eb���
]1T*Aq���}j�Ћ�^5���A �h�Hx�60Zo���lע�0>�T��=i��F2��`���d)p6�s��~q�e}�Ϻ���T�-�a8V�d*㑼���n���&�92�hj�-�8�P�[��oV�/�^��oY�VH>)<�x��7fu�&u�OT���fAvz�z(���Y�O�^���W��8�3V85�v�����8�>_�\��F����6�fi��Xֶ�+P&h쯺\ �W��%�O��mt]��#��JT5`B��_�4��3V�*U��+.œJ�0�;yq b�;���Ҳ$6o���KD!L��EUמ��$�Z�8$���9N�A��i�Վj�_����bv{����!�,�g����9d�׉%Fc�/�;���C������k����a]9�r���Y����ݪt��X�C\����;���k��.�I�gKT�ӛFY�ي��pl�V�[,F����H��1^�������9Q�뮕ԥ�X+�?J��]3�W+�xO,%�w������{lT"����ō�|�|��1I�X 	kt&u��׍��̗w���_�ո�Ԗ�OD�F��X��H��]t[9��r8%�ڴ*nr���|IO+�z���Ж��3�{���C�U_�.����є[o���q�.C<A�b�a,��ە��y]���;��5ߑt+	��fݿd����:�<>�������J=l��Е5��{P��z��68u�3��<_�G����%C�r���u�1��]���Q0����h�����7a�I�/L�-ػ����&�"6��k,=n � � �L��m,�-�{����p����J�u◝%��w�GH_f 1�ܭ�&f�������$����ZZ��&H�RGj+w1�Ю�]�焙<	���u�g���q�F�j d�	�ӫ��J�#y�^+|�LtNr�
2W97ny��qn==��I�i��CQb| +j�R��������ǄG�3u�AtG��W21�z����/��Iu:4�ԅ(4�)��X�����_��]qO7�ŏЛ�Ø�y� ��KL0�n?���z}٧t4E¿���Ε��ǁmmq��xs~�ɦO�:C�	.�ĶZ�F����X}n��DMy������,�1�2�[u�f�x����f��}�WU,1���4��O���ro��e8	x���Yf��K12�w<7� ��ա��L�v�������	-�m��x��������~!3Ǝ�5_�aL�4z�OWT.>׽VFڵ�<A����?����F�1\�X�4K�N����X6ω�'_��> �d�p����<�d�K�^�_�)a�5����򨒷��d��z�����5���.h���7�wc�B��%n| �5�@�)=`�ؘ^ e"ƝrT���<�}~S�����oy�t\����L3��y�`l��ا-��說ھÑ�ln�B;�.�r�@Ϲ�z��� !���<M��DK��bZ��#���~�
4ZZ�$ȝ]����4b:]j�Ć���t�Q�9��}�B�qC��olI|�,��DI�SG��A�4�u��T�W1��"���e��ir&�Y�0D$�7z<9��±��5=0�p� �"8�2nIV����96tUp���$�O�A^���r�Ee瑖�׫��*9���z���?�$��*�Q�*r���'@�{�wiK���P8��[�i��QDC�	�&~��40�n4QJ�f�vۂg�Mu�b4���w;[���! �@��Pa�-G��<�&�p���m5�đ�p|�[���j�!%��wv��{�V�l�{'S���a|u�>y	��*��NF�2�O&`� g�kք'�No೐����羌0�N��J6�� q鎗8��=V���@`$�P8�s�)��8��>m�١� <x�%�:0�[�@% V�h521���ڿ��廟�g�\�!m���?=o�@̉�VQR-�6Z�� �e4�߈~��aZ��#t����U��*��JB�Ū��s�zg8{�肗7$/�=���T���ĸ�k�n�G*s5�HW ��б���n�%d��
�M�`3s4B�J�`�<�ܐ���B3z�u0��y���G8x��D���L��G�H��:��ȗxMB��u&��s2oB��ͼ�+K�AY3h[��͓=k�Ȉ����[n>k`*�Hc�.fr�]Ӽ#��:y�7��]PR�����ͥ�*���@�1F�4;�Fz���R׋F�+Wv$�t2Yha;@���9n�9�A�^O�����$�����q����O�d9J��u9�l�D$�$��$���ʱ��G&5�gp���D�>�eh���WۣჅ�H��a�Ө��ʁ��A�K��0���9_'�2����$��4x�g�;�Į���6A��$9�I�F�nT�H���h���,Ga�a��}�� �KA�T8l؉�؏��H���n��,p�3�$I�7��-��͐GGO�;R�ߦ�$LT��u|o����+*ֳ�7"�W9�޹�oo��vj�myw�B[>�y��0"gn���}(�qȃ��v����#BQ=���4d�/��i^�et^bD(����b忬)?Ս���^
.��z�;��I����_��&m�E���G���F�1@1��m_=�M���Mw�f�Vˋ%ý��o�H˷���:, 'm9`"2�[U�j?���8�_w=�X��(��Ð9;�r��m5&���
	plZ�F�O������JW������� Rˈ�]�����Q�&�'@d/�dS��$5����8����K�-6��C[�)���D(��(�-�G��7'�y6f���3�
a�`�3�qh-g���=��k[�K-]кF�����h0B���w�@���$W�ۙ뀅���`�r6���Km�����H�`�Y&����ث���1�~2��#u��L���!B-�������%�8��#"KXI8v��.,����.�^bq�����.t祖��p��g�iDu[��q�1�Q���s��Y��j�`��:p�g�U�-<��6�1*/�.Ț��2U4�o�����'�����U�i�T[$��p��L���U�k���L=�^�X*���H&!��/�ڋ=�\�+f��(J��ꑨ�+"Y-�d�p]�  "m୚Ԣbl ���t_�����31�WG��ù���USd��Q�e�N�5O��/����3 �68��g�@@Û���@�/p���-�sc�:�2����^���O�n#"1�,��.���*�k��)���ba	���*'r���kޑ4铘�Ň���&FȰ����$V�*�=q��{����>)0�RD�ЍJp�q����sWS�C5�~lFb%�z��K��e��=e��/��&�����)��@WZ��*A�#Vz9��:��RgS�)jKi"ԒF�h�?ǔƛ�,�[��]���ތ�i�\n \<�M���w%���.�'�o�,y��u$fw�%>�ǈ"��0���/����m�ug�n[��&��}�Ͳ/��#��n_�1í�?��{��r��W�>/���X8`��c����sC�`�=��o��ֳ� �6�x0��O�6����؏�-Xu<���3hr$K~�j�	�($�m¤�l�;�	۵�*T�,���ed�o���wD����T��ը�	��5�K�C�Sد���m���Ha��#�u�S�щqo�PK4�Yׂo���7_n��,��a���P"�#H�6#L.��E�L��xu.T7�0>���S"�qH�#OK1���0��s&��c�䈵�x)m������������Z�,�	l�a?6�Yj��]����Ȝ\Iډ��6?��+���;��'�L�: G*���f�-<4@��6Mn������s{��� �7�#zZ;v���L`��!���� Հ�-f6h�X���)�Ʌ�n��
�ݖyjł�rCý���lPg=�������z����ڳY���2���L��3oT~n�8�$H�B�bI�d[\9=�|�Q;��������������"`LUYwTvL��3�4�� B�iX�d��`\A�&�d�,��6θwN��EޡPȟ�~�~��CU�؉�{��vs`,��������~������<PTfOUn3���n���oHݱYm�،�uoH1ͮ��I�,[(�����"m�caHZ��j�-B]�O7mC�黮��	�w��~%B,��f�q[�1�/���dm��f6vPv������LGg��N�f$Sc��0���yh�<|�u; -Vp�@1[ԥ�@i9��`��Aڙc^���G��;��m�0$�H���
�J$��
o��s����_v�m�X���l���c�^z����&�Sp�!0?g��F���$RP{�s��'8�;�1F�'���okY%����N�S����fX/�2u F�0�G�q��)=��_�߸�E'I~ �LY��3��������CFeG��6�ؘ4w�,;����������wk���EF"꼥kVW�m+ҙ�쀬��3�e'���17��ݱK#�8�b ���>؃� �2"]�� ����.��ȱ�A�G�����tꊞ��kb@]���"*��)�{B�͸����#>u�����R9��X!iCD��5r|��Wt�Y;��$4�`���FV��Қ�������8�a_���\߳���ܠg����f���h_ς_��W�Z�=�i�r9]N�y�Z����+�	$�Kl!�J��ib����[R��>�'M\�$���K�8�O`�M5�`Pf9�0�C婑����7�m��`,à����`UҒ����6�kh��]��N=^�Z���]�$R�_;�V=�AQ�d�޿��Q8_� t�����j�}�S���T��,?d��v8�tA�
����c<t�kW*��t�%�R&��vm��D�k�g}�R5�Rc@{��Y�	B��x�m�5�ߠvm�!�=�wQ��]����R�Y�����1���q���.~#c��r��f�wC��k�yT���T�lo��Z�D̃@6����/�z�=�����L�.����k�Qڻ"W�A��|(��=��<�ˢ~�4��9˗Ey����=�!a�\z�:G"o�hź����/sqe��q�~���o31ޟ{�ՍQ~Q�a�K43���M����_o��ac*�ڷ�������a�(z�.��5NQ���$��� �i1���9[��R9U�X��:M��o��Ma�S�8Z������ϯ��c��_�qI-�������lŖ-���Đҝ?�Q��:z]E0���c�63��Y��F��fV=hޮ�H/�Q��@w�^���-�V���#��N���	�l��0�&������ŤWT����=GkK�T����:������r?3r����d9h�|�D�R/���ZR����$$x�I"<Ć�=`I�8Px���9�ۤ��!�0��R�ɢs�Q3~S�t++�\��|�faI$����izSE
�U����a?�b�\$*�#{��Ɖb�S/O�&�$7|�#>A��՘C����E? ��>�C�Պ��̻]'�s�%�I�]�j{�����N��-��F#�f�|T���4D4]$)�� ��_�b�ceZ/SN�9��W�Cl������aW���^��]u�i��i��޹���TV%>0������]�?2�\�|/iK�џL�����T�C���R��3������r��#J�+���)��]�b4˒��_���/H�>�C�έƠ>TH�N_��H�SWh�@%H����Ů���q���q�To�ֶd2�[�As��nU�s�eK����>ᯙR,
l'
�um���Ai�vv��l�g�@7�'� �IMX��BH7q�X���pa)�hxdj�y��j��j�[M���ŷ*	΅���t��}�#��m��^���@x$�sljoa��%B|(q疹4�ago�J�f��h^���TŖ 2�(��b�)��\���Uw�l��*��O���%�y��*�U�g�mj��g���T������܊=|_��q��)�J�y1Q��}�M1G{��cFU�/'�U�a����xЮ�c5�1wh�X�ލx>�w )�=��uv��Çn������{�G~�QĦ�^8�F�	FEŧ�X�4Fdt��B���˯1�n����k6�Tδ�@�T>35nda�6P��J��M}Dُ?
FJt`K�-IZr\�`ie����"�� �ud�}���r�҅?#V.(야�:���6��ߝ��U�?�鄢E�g� ��.nR�m�ǖ��'U �qk�p �"�W�q k㱞)NעjF�)a���I4>��``�g�ou��A�>G��-�R������%zˤ�r��F�[�m�=����p�\�[m�ϩF�5@.�K����&���'D�o�t�ф4����J�3��D�Z��Zvz����+V�H�`�r�� -V7���S��oi;�k��~���������HGOn���01�⷟�h: �r%A�]P?$��h34�m�D�L/�)l���l� ȫJ�*uT��/9X:� �.�%��+�X�]x:��jP}�4<e�&?�op�i��g��5�"(�F�p7[��LY�j�]���P�����}@{���8X�\S��T��%�}r�ZV>'k�w_#*pg(tD�%�%��>y�IM�}}��!<��<fR�n���J�x�N������h�ٰ+��:������I��n7�^�o}��a� 
���"��I�68��ˏ��Is�<\�W2̳�S.�"ML�V'03��
��+�~f׳y���C���}��*��!@�/4T���]��m�GA��[����h�)��_FC���W���<$'�ҽWTR�29�'�\���O���'Kd�vfQ�鶩u�&".�i��}K~=.%�2}�Q��G�w�i���E��M��Q)7��/��v�S(�Snzc��d���RFW"��f}��,�!�#�^����'��"7�V��f<�G�!"_���P�T�����J�:Q^�*��.(��~�F�H��d�r�����H�Ԑ��* �t��:<iW�L��,H��	�Ơr'��ʘ�1~���C���-��h�O
�4nMa���Ŗoє�
�%����r��xo�
����W�PӪR���5�2�),7���"���� y�Xd�1���2��I�"D�1�3W�kv����z���`���V������D1g�~4:��o� �m��s���I�Aּ�?=��(W;�$�x����7=n�ޔ�@�W�v�}�s��x�<���>~���K]�gMQ�����9�`�2jJ$s�ɸ���t9��9�l�,��&�,@�:j��V)8y�$��Tװ?݋&���	�TG�X�*-E�X3���|0l!%�^�obU��2����7g9�h&x$?(ھT��8��e�<S�Z-d�U�l�^��\p�,l�MQ�aجE0!_ƈw��tF�O+�l4r��=Ű0J�3�D��}L�߹m����܃HC���L�I1����wУ�SH�Z3�/����\z���li[p�]?r�L�[
475o�Ŀ��m��K�m����$�fC8ǌ��(��0�X����:�Y�U�p��˥�I���$�#R-�����Y��U��wx]���.8�q���Q�/�2��� �1��\������!E���x����FѰ�jE~35⏸#�#Us˨��H��a��d���R_^I^ޣ��"eOw�='�s��Y��L�����j�]�82B�tx��oV��7T߁��~�*��f���c�E��{����;��9��Q���*X�.:X�b>���c�`,��us3zx�i'h�&l&�v��� T�B걗�ʳ��Y���V��Yo!ѓl�|M����?�.O��S[yN	��Uc� h�����7R�'`̇�t1�WZǫp��F��fJ-oo*�
E����� n	�9Y�(PN��-�P�(9�AW�]�y;�"SxEB�!����/���	,;!�7s'w�$#��v���:��S���X>J�q��7�7�v����3C�[�e_#���Ը������\�5�}h��[d��y�_�����1U#�Nk�laqY��t�^|���,�y��^e������ʹ�rU�"ڃzM��h@�N���~?Ү(�H���'��^�X1i���l����|�Ŀ�cS��ۈ϶�����A�gM�u�x9������`���6�=��E�d+�T���=l�N��n_�5Hw7��e8� ���:�l茖U� oh����p��~�{A��>�t>�R:5�~�2m1�o�)�����G��3O�Z�N��VE�
(��%�]��Aw-j'l��X�R-�`��$�[�=��
�m<�f�N4E�ǌN�D����z�h ?)^����U�����)���~��3��Mg��cf���p-&z"�N)�z�リ���
������;J�p�+#����A
7���)3𿡶TC�x'^@(�uOe��Rڱi-����<��o!,Υz��e���aۚ�j�n\��f�(�ٷ8ۦP�s�tz�\)�����Nq9�Q�rT�7�lO�ށ
����bCE����w�}�`L� s�X	*�"~'�U���'�$*���]�s��҈ت�4I��`���q���*�� 2��^ګƮ�)�TOQE����׶Hܷ�ISSnZ��&*7��1ґ��5���j���\��' �k����fԸ$��zP�aB<���kW��Z'X�d=*H[�ȵ�*�J��<�^n��4��P�?��t4��}���~*������Q���$Rn�( F5�S��s	�n0:��F�knY��F$��ށE��mҦ�s:y�y�����w�?M	!�p2dߎ�u�����C�eXt%g�P��;��JwX�^�'P���Lz!��y�Ɗ ]6�g�N��4��8���Y��؍�|v�"d�}�+k�Aa�Э0�4�5�Z�wl'gҗ[��s K�����Ж�#��L���%��b)�؏ɜ��������(�oI�s����O>�!��_��xIU���R�Y��CuS^݁��k-k`�3��?Zޅ�W+������y���U�E3��hk�^�������^

���᥅���v�FK�*z�T֮W��(�.&2v�VA����􊌔�;nyQ��Z��Un�Q���/H~?;u�\�;��ڀ�@ߢ��g��*K����ܿT�N�_-P"Ke:Lm�����<�I�
Z�Dx ����j�ͨBe��� ����Z��1j�߄������@,m�� �c���f,���4{��ҧvYUf��!%?J�lQ��ť�'�k�����K�B&�,e6�X��^j��b5�=��P���C\��r���+F���[	��qꇰ�pX[;'��]�(�kd�}F�'+U2^/  bSӝ�t���D���������8��>4����W�O#?��Ȗ�!�7yFO��?�)��FoaV��n�|�J��8q'E0��v��Ǉ�G���~>ڞ1��2[Ii%&���٨8�Zv36���(
�ô�i�C�|^3J+��n'�`}i�i|���X0F�L~�g��W�Y�cB�Q/ ���9y���Č\3� z��d�	z�
�.^�/��$���)��;!��o�E<�oW�r�EsüU����r���u�&�4����F0 ���J�� ��U�ˢ�(H5�7�G��]��Z2X,m�����4�w�a�&�����H��	��0����u�R�ɔ��zQ [}5��Z�B��
 ���K�I9��N�-�@�j��~O���9���M|�q��xU�����.H��L�y��Ņi��Ϩ��%�z�*�Z�홃ޛ0�ۺaY�bS��18:G/V�Ѽ��������3˼aׄ��F�:A�w�O���E�a+ڃ��9�������[?��/	B�����2���?�3Fo��M����bNN^)J���k����� :m�>?�2>!�v�f�&@�gQ(��g�[N��9��N�.3Vz�hˊ"õ�jZ�.�	����C���T\��	Y/#��$��q�p�G���Ԩ�d4��x�,����� �$R)UA���Ϭ,�e�_�����[�hֲX������� ' cCxۤi̳���,�@q�7[ŧ)y$���U���"���F'�3?��M�jh9}�R�$���U�����p���l��>�ؓQI!����\�jE� +49��g'��O}^���$�����I�����e �u(Xaj	��*Ņě8{LĀ^^W������b}l�)�ӰY�@?縵�0Y�eȓ�/�b��0��P^��N�w<k�Ul�2˨z��5	��a�������1lt;Nӯn[7�蚌����cH��V#p�'!>5��9�9l�@⃨Mޫ)�����q���qai$e����o�/�ߘLdzp����nX �t�����UP��SF8�j9+�"8ʽ��N!Qa�ߴ$C���)�n��ȃ^�_�\3!�"�=���sd@?G�'H������Q��F�ݺ�h[�����(2:0��Va���٥#�5��w:IO�B_j�w��6,RU����(�HX[ǐ\�z�����s�62��CMi�[�Y`%���J�6_�y�vS!^����_`����,�S�I��6'�ŧ�z�X,P')�U�b�Kъ��`.�9�D�+y��K���JEr׾|�� 8��v�w�FIf�3spN�u�Z�{{GB����鏋�N�t����g��S�K#<��\�W��"4��l>�o��&�Y|��M��.i�R�|���'��奎�	�Pe¸T���(G���ӳ��O�Q�5�$2�����"����1ǐGT����W��-����Cb7\µ��#r��ïU_5���/���-�a@=�G']{H���ڐ�8+���=��/���J=��˹�����b�Փ珏�zs��1'�`p"�H��k��Du!�MƝz��.�����aZu�M�g+�����1[�	�Y����k�BͶ�8�B|U��5���N��#�s�ј�k4Z��e��?��md<��1��b��"SL����1���KʱF�r
Z�[��*r���g�d���\
��,j�B�Y�J"�3��w�7�Zgx��;�灭/r���a���D�����:�T\�
|�q7?dlO���[�z�r����Bt�x�������[ǯ�D+��|�����j�%N÷�tl��]<(4���+%�
>ac� ��ԈW�Ը�CP��cicW�4���)^nYؘc��D��~V���KŜ��äTl�{�(>p1�+�5�ɚ���K5��o�2��YN�%~����9	�si��@?j�bn��K�Dؤ�FA�Eᦆ�cK���\��51' oq����wv�p"V�f*��jf����kV�C���(���@ j[��6k�d�t�7�0��Ǎo6vs�	E\G������[b'$,��Λ}�׮~L,&YU5�A�E�}:��&r�~ մXV
�(~l6��t����6r�T��"�?�! ԋ~�DJ�o���%i>*vAd�E����vm9Oj��%�/�a�e�.r�r67j^���a�I���x���g�0Ԡ����H*��7�;G0�����-ފ�"SJ��u���	�J����F�6N҉5z�TN6������?��8�ڡDt�J��4�#Z��Yν��\���N����0�z��20y���+���͆:&��O��	H��@$��'T�i�aZ?JO��B���º��H��A�W��>%]=NI_���&j6���� c=��\�[-׎�1���(�q��/��sX�d�I#܈�4Mᆻ_%�x�L6z��m�_#ɰ[�W{�ԟ�7�����~*����b�}�^�ܬ7
G���������R�P�D;Q�,�xbs`$?�_:%z��yET�������[q�������@.y�`�B��y��5������OD�g,�H��M	.�\��NH��eCx���誊>�����ȥ��u���pI��t��28����g젆����)�/�G���ԥVc�p��#݁J�f�Y!��c¡fp �3Ӫ�`!��a������,�� b��>R�g�.ѱ��k�	W��7G[[t���v���}S�T�o�m|�]?�G��w�Y����NJ�4�9p��ףiZ������ %A�%d�j�G
��у�]{�p�8?n>1�iM�Ǖ*ON'�Љ �;�����2bh��0#{��\1����E���}ǁ�Њ�i�̯y�4�"yO�����sY�E�;�� ��]I^Mz��٥�jKž,�Y2���z��ۧ����������C}K<��}��M���f;N�v�s���D/�G�wƝS��_Cͮ���d�Rќ0z�Ym�څ,\ �y�(�ly���>?0����e��@UL�"U"]��|t9��t�f��e:�\�Еȸ1
��۪(��U�ܕ+�?ٍEc��:I���1>��a��K������lO��FR�~d���Nn^����GA�	սI����,��pW��DBbkTD�H�tIc��!�}G�K�$\�ϔ�N_�lL�����cF���r8.�)������~t�3Ŵ;�Ʃ�
w�Pmx^�^�`����8 o�Ʉ��5q��u5��+�Qb���&͑��W��k�蜽ql��#T��c��x^����]�qk��xV�]���S_mk# "-�'�����y����x���S�!i�t@aA��젍��&���0���2��2g"��M�6��n`����B��  �v�YOZ@+�t���_~���g@�z����|~����mRy�-z�)^";�1��`vI�m�f�HG�����-��Lxs�$��3e$���DV�A_� 7�ڏ��zk¡�b`:��e�W��0�$8z�o���m,?7c��9�R��l�C�.���	]�0��'@`��.�V[�m���8�/dV/,�U�g��)[!�=&pB�S?�F�_Y�\]ǹ=�m_e�\�5�J*��"6��ì�4E�d� �,:J�-�I�̮24������	�6�ҧ��B{�/En�I�Y��.�u�[����c���\J��o�U�=����!�x�z��F4"�-}��o�^W�Y�H��-�Xm�K3�Y&���B�Q��8����:�]�4"�O�b�D�8�X�g��<�Ű <lP�r\��T�A^���I`�+�7����jH��:����E7������-g���G �"Ĵ�8F]+1���R���zM��_>O!^����ǿ`Do�d��	 |mp|֡؍Q/��r!E�d�h\��q6+�K���	ߞ~��]T|��D`}@M�`[�#^�[�[�3�Ѫ�Nڧ3V���#xpn6<A����d�Ve0��� ����ݵ�����=��J@{|'N���-)�ͣ=*�����{�r`��W�~ÎI�z�h��R�I��?�Q���Y������Kj����0�돱�(��������ۂ�)���%g����@�ZN8)#���^;�`WS,VΤ\�3���ZO�TC�Äh���đ1&;*�qPGȘ?��QS����H�<@nY!�V(����c_�O^M����74p��VB@�~Y8�X�ډ<Б����1+6�f>��.y͌�,��4Z}�N��x������w��6� Ǻ�E�8� �!g�Uu"
-yEj��"]��d��n��tf���]�w�:ԏq��9��(THth$�0��
&�(.D�7�^�����i,�*I
*��mň��&@�A��[��+���$��Qk֜�~lmt�>����1��ژ��įA[�.{�ᳯ1�cU�m˲q��y�Y����bk Ƒ�2��0��/��9��Q�5�1�����P�7_���z�e�J�\�\�p�D:<�>
�RQ��ʙݱ��y`�(gG2�wy�ɼl�Y��&`�����yA"�#/�9�	t�+�@�$,pG�i�pY[=��{Zs�9�ƨ=�>�~�[��FC�(��j��l�C���(>'*�T�Yp��#��3u�;2�����N\%D_h��K$�8J�l85~����z��$�,�vX;,$,J	L����f��aI��a��!��i'*ODr����2�f��[��>�ߒʏ�m}YmfI�W�
�gu��p;��ݻ�A��|N��߰W"��4���$9,��j���r�U�����b^G�E�Ɇ�|��2��֧�5̑��'�u�������}A�e�q�xim�z�����z����HU���:�H��Ĭ��X?�Hn�o�W���w��������0���2l�d 햤z�O�4!7������;Z��ˍ�V�"�گw�G)���䡾��=�b���R��Xj���q7���ό�6��):�:�	������DDZr���3��4�H�y��ҙ�{xMρT��*��t�7�'V$���B�3�]���z�8�);���԰�繳�h,�)�U������H%H7GRf�{H,=]�S`�1��gR�K
��W��w�J	[e��[H8��[��.ldR�$����υp�OR�+?a�M�g�D'�A(�o��lܙ� �~����@�w� R �v%�;9�7��D��&�`�n4c�h��s�<�O�䔤-�`t��%ՊmTpqnq�Sd�|������ɬ����cG˲�4�d=ܑ�����Fnj�#�`�lj�8�1X�Mr���@I�WR��FB�/ҿ��_,��[��,өPkH�����!�ift��<��<�º*)����))� ��������C;�O�Yqع�Ҙ�:<ɤUC��7@+C�]I�����Y���nCr;��
��ڮRJʹ��d},��%	S��ϩ��v(c��$�y�5.�3#b�W��~�ϴ�Wd`f-�lg�<�I�|��D��~�x�SH�������*�qC��W[#���`i��'����F�yQa�Y���~�!���DZ��-��b��^"]5?V�(��kU�ihݞ�2���c��n}��K�͊}3���Ҋ�o�b��:j�$��Md|��o\+u�'����8׋�O������"ݤ�CJN���$q�Q6��y�y���$�M�#�d���Z*����#�~M�(:�E�Ϛ����Q'�����}��Ɖ��=�7Ut�_-�ʹ����p#�$�D'�)N�)K�Wm��+y�z�e��ł��|�>�>X�ϧ�c�����g;����{<*�1n#>j��D����J?�f
Л|�E��wC�$�Q�t(ۣH�Z�gᴌ�����MقP:��3�tN5����TM\pdo��O�W���*!<��[��*%ݹݝ��5��(Lϊn�#~W�G���6��z�1'�܋Ssg̎G�����T�x�a�ï{p\�E�>�x�\>�R���IO�P��9��x�D��!�G�@�D���:^{I��IK��|^���4H�G܊h��T	���Y�`:�צ�����M.YB> k��G1+q ��������2Y��f�$�J�)����*���G�����}��Zۚ��&��-����)��~�6�"e�l��nԳ����ӹ�w�l�G���i�a�ݬ�K`x����c��}��	>P,�2�I�c�^L���_���"*�'���NO+�1uM�޻�%��������w�1~���))��V'䦥P�sB=9��iݫl��J7���A���u1,D-���#AP݌�� �q�3%8�r����'�΁(:����W�	��z �v��$���]&u�v#na�iz�V
�l'/=㊱���N����D���>��`�c���Ct)������0.�5e/�T�0��ۨe���{=.���i����c�t���P���_���շV�ʤ���BϔkZ�hD<1(?�4�KײSZ�pٗպ1�ʘC���:9Ÿq����2Qv}�F�oc'ȱ�4S���T��~=�P7n��EjA�O��G�nbKk�1h�6��}�0�X�R���%�X$mIWBvL����Q��S[1�s����uw��V�d6
�d0o�X�cA�%���	�����؛��N8 +�xn|�Jmg,5���-�H��=�� �n0��;�Z i%|�̨�G�M�ڤ��������H�Kԡv���=O���rX�=�{���spq��ᐺt��lM�����@ݯr}�<O�+��8(���cb��w��3��4�ލ��p3G��� ��řg镗�Г`b��d=�0g�v=�DΨp�yc���s���x��"س�lUy$�7��`OX8�u�7�l�X�D�\�0�cn�ހm<�z����%��ӷ���`������;z�|��}Ne�p���t,|�+Ia��L!�&�����{8�+�Ð`(�#)�%�-� �_#�R���~��O�Px�;�X�$�8�� ����W�J��3fnbm%�:��h�NN���3KM�I�L^Q���AU88�t���#�c�zoh_�W�y��SJ�Y1�v��%���	Ǎ7�H�����ߜ"v�����;����|h�q 3`̧i�}�C�U���<N.I�Wf��x,b�VѠ�iR�V�f!3�W�5<�^�������jr�=�Է"�k�G)��HϜ��=,����` a�P%zW���Tl���?�Z^���s���x�E�L�!9����3�M��ߥ �O��}�=Ta�X���l�h���=H���G%�g��DH 4�R�'f(�=������|c��3��y�n",�狓��W��}U]J�E\�0��/v���'��(34���#��7)�M&�E�	7B4�|7�J�%��=���d��hV
�� �N��^�v���[z��SU�F������0�����hٗ���KpG.;Iw�K9s_�0�?=86������l���+o���8�co�|R�N
�?�X�\xI0���)f�n��~�ϗq�!<��I`��� A��l�wŲ��o@�� �=*�0����E�ۂk�D�j��lsb)�'��;m-�G)uqleJ[8E��[��q�*�.�Z�]�j��<��\r�x����H�s�����ߑ��mb��EkOH�c؍< �AIp�~!)� ��-%���m�I����Ce��K�C�X��7zo��	ᘩ�:۞[\س+�Dx4�tf=�������xo�Y2���ͨn��{q�b�n��1���D�k���	
�(Z��ؠ�hOB8�^ݢ�EI(~ed�}t�(6o��Eƍ���*�$zyoE]�:����^C�!�Y�=X�{X�[�
D���K��=�<U�c8���1�IAӮQqՁ$��C�ߙ�D�P�Ιx�j�99������a��{t�c��`�Mt���L�,�+ux�ϒ�i���%�M�{�� ,���U�� ����)�Te'yU�4;npCFNB��;ZU�i\"?H�شjm]M������\���%"!I5 �`ф@�
��.~�X;,)�3)6�,X�=e����㛻�ӹ�a;��O����V��b�1Ē�q�b���^����@�]�t�w���_����Y�p(���=h����]����w�`�����,�X���b(�
��DLF`�j�2�e'�X��\jA�sm��G�[�`�~��z8$Fg��g�o5B�*)��pW��?���d��M	���tF����4�P���r)��߷������"��kx{Mj�(�9�d��Z6
e��lY� ���� ,��ņ��1G0L?�՞�IZVD�ve��
���^fhgS'�4����:�?���&iŎH�"��Ě�(��.�_�x�t�N�+��(�O���7*��Q�N��|OH4�\^�@
�=/�ଣ&���#�Y�jpP����fi<������+��z���xo�K�����<��U�q�PM�JRp��q��`�e��V�J�Lw��i\K}aN������蹱x��|��k��i�K@J��~#[��=!�ӱ�P�O���wӾ�%��Ny5cN�?>��6s�}w�{v)�{������=� �,&w�.����&>����'[�X<G�0BE*�}��_V��j?�i����4L�:�h�8��3F�dC��!�/'��`d��,��6�?!e~�߷�u�ĒaZ�c��Ç�TPD����x,ڲQTըyQ**i�կ�ӳ�4E-����իmV���ÙQ��FlۛG�F1�.���lХiEYSr$�D0�+r��õWk�Gw��,'�s_�po����D)\�j_T`fՀ������c��V����H�h�MC��!�c;<��{I 8��v�}�f}>󚴃���^�s����Rhp��� <4F�bxy? sŘEi�B�h��"-�����Iv�ex�7�����Y�w��R�J[�o���Τ�S��-��0�_�T�{]�E��3n��qn`С���l5�qsû���������/��T��t�$ª[�Q����׏���E-]���
�����W6�&G�o�U� ��f�pN�jl�j��:�F<>k�z�)�;;��~��÷_���_��B�X�z�-Ez�ZZ��ǋ�Ti�M�:����� �E1�2��^����]�l&�twq���S3�O&�.��@���F�w;d���v��˭	ە9*���C�R9 jU��e��gy��ڌ��%!�x�F~xb���B�� �M��}4r�dQ��ף�1?��U����P0��~�̱j6�PC5*2Y(��L�-�KY �{��ǉ�>Q���Ҏ����<F���ڡ@�L������Ú�QQ�>X����	�h�.�5���i�@��Ƨ��[�+h_S�eh=�[��@�B]>������^t�1!8C�'���U�q�V~{��84i�a֕��n0��}Cz�� �4D����vJ�ڟцλ��S:V�~�H��󤚨I�_�_Q#�0�p�b�+HE���3�R�I���#�{���>�	��SS.����(S�7�ׂ Lj������4GD���~���$��>���<@�r��(7����o�c�ڞ���a�v~�h6�M��s�L��
Sp��ܿ���T=.XY:$��[�I3_����v$X���R�g>�
}�ű��t��O���n��vġs?2ȒK�����
߳�D]+�P�RK��/Ԉm8'feQԯ�w�%��v;@�*��_�YdS=4��lp���'r��r�幷,h��:ya��T@7/Y7��6>�ύگ=�4e�|:i������j��lb�!�z�K��X�_v��,l0��Y��X>D��%D��D�_�W�� ��N���k�籥 ��?�s���֡���7Mf{��v��,�_�x�(^x�
ro�u�s��P,2K��q(�@lFM�ß�o)�xu��@�-�􇦻Dpmm֜ꙡ��M&�*��Q�@"��bS}�,��\��;CX���^a"����	��C$d!��Ka�6�~�ȀN�n(�?�W�/�����)-1�J�t	u�{�A� �0M���u��e1�%S.�O��C`I]��r ���6p;�@��kh�l|ۄ���v�����B5�Vn�
0
���|��w�� وI�@FC���b&S�s��o�Zl���?)����j�K��$�e$4���aX��]��bxۚ�KdtB�=��@��5v�c�M�a�7���#�򘺦�Jm�ب�OfX�5�k�Db��|d缥����9��q`!-�[��AP���	�{�$��k���8�!�1�k�ɣ�F�xV�W��6�C`��2"���.s�E{j}�0)��@�^���?��MMn���Y~�-�Za���8��˩���%����N�A���I����^b:�z:I���YB�!��d|>�z
��cZ�a�c��j��/�� ��ًa�L�ڪo$�3,�4=�U���u#��>m��h\��o�Hf� Y�a 4K�jC`֨���"��Mc�%��s��b'J$��$c����alU�|� +�%o4�.�=�ŝ~�φ"5!}F�����q�ͮ�OI���s�!��J���?-��1g
�Pr ��-Dk�[a:��S�z��Q��Z߾E:��02��hz��ݒOܫd ̭ɛ�[
@�� �
�cv�^z�t�ֵ�yI�څ��|����ô�&�b̸��24����*���)E�|� �P`W�
�d 7,z��e���?r�V#�{W,��MU#XH���&<�[�a2A̬B������G���h
pXg�t0�a%mV�����d��~&�,�/�X�.j��4W����O����y]m���x~�����/,\)�B����F�1��R�h��8U2-��\9Zě�|&�R�Rս�>���D�'�]�1ԇ&����<@yR����/}#M{�[��{�@<�)2Ԇ~x���xD�����z>1ϰ �<��e������v��U�*�%R�!-��G�Q�^��ibw����h��%��ev,b��9|�r��'z�7�V���;n����Y���;+���׮Q�E�V��8��{��9�q1�b|qHESՌxēi2ѨJ�l��DZ��ޞ�:)�C�H��:����n��m�2�\1�-���A�NO�w��N�^�F�x�f����ܾ�/4�nd�j�S�>����G�&�}���#ѵ5�՘�<.iW[�P�:��
�{��9�vv5�L�C��X|b��4��H�Lr�|+q��R77�դ���!��M	�	~�������i��Y��&`=��Gnƶ����8C��\�r�����q�����)D��J����.<R.�_=�%��˿�N$!��S��R�(y&�В9��
HR#�x@tQU�s,��4g=��oP0x 3g��!����_yM�po�+�@6 � ����]�b1t��\���`�gOM�6{�D�b"��0gG@z�~��&�88,
B��}�y}x�xF!��ou�f�.|d L�(�DAJ%Cz0u����Fw��K�Ɨ/���$@*����Pd
�.�A�IA���Xp ~PX!NC��N98V~������Z,�û'@�#��t/�����?��N�S5ۮ�܏����H;�����
���A�z��fG�=���c��X�H��|k������y%�7Db����:�)�@e��r�R��q"2�>�:l(`9�D�i(�>c�����H��:�J�ŐYmT���5Y��(r��� ���2S�Q������>KGƤ�!e^h�s��h�� �*�@�O��H��Jǽ�0%��+�|�/���w/�̨�/tލA���X��oճEw��Km�a�e�Z���~��FFw����8sB���B�Z�:>B��U���Ŏ�D�)��������ui+��*3��*�Q�t���[�Fc�ı���s�IZ!��4����~D��{�V:�����k��SwT&�t��T�?�C*�ʆ��K��sȪ^JShw�K"k�_o疉��r+����Qy,N�G�aī:b�$6'fZҘ؇��IgO�={j(Ir���ex� ,/������w��7A��wMn�VUw��ݦ&�hy�M�� ����W�2V�����&{�;YGF���Z��g��-����L����J����N�+R �	,5=�*kg�cX��ǣ��zh�pk}�v6Gv�L�#l�5���4T41P͞���A�����h�@,�y������LDƺ�"&�W���f���iB��gù���9���q�ؾ�4����l�����e�{��(��l5HT��+%Ma��e����j>�Vǔ�:w�����ai�I�v�{�i�vՁ��7���QEG�@�����1�IN�B^�R�+"|\uU���e���ZT!�j���� `�wzV*ҫ�ñ���J�U�j�'$�^�0�����|x������g�	(�ds%�gם�Vg�yD��j=$/�1�+X+d�_a��/�S.��<�~R/SQ�UQ�GU��e �L�{ƴmZUzg� ��!uh�ַ�}�YE�0��7�M��F��)��c�J�y.��b��Ss�����崦<%i78}�[W"�9��V�y�fs��M�3�"X|�1����GE�����<<��ji6w~V�2A�,j�QNͪ��V�	���8�����y}ܿTMZ�p�0�ҐM�RA!x}�W���W�<�Ā;#��#�r�c�s�q�����ފq�ͦ]oP�pQU��@�4�b�o���GН�b��s����i��'��E,xQ�/�y���)h$-j97	�w(hwS�f\W���M�P������[	8�+[Α���6�=��CTս����J�r�v�~U�R��h��֘|O���`!�{5��oK��W�y*�+�g��� `�⤝e�ѵb���p�U(�^��f��+m{�i�<�� ,L���������Aw�����A+/횋���qA�x���E�C�+�i�-E'��N!KȮG,^��d��+�M��u��>l�{�7�5��d�	�略�Zv�%�F&�G���d0�Wȵd�"]���3��h�)|/�y�*uˣ�-�ף�����h�q	��6z6����J������y��I��ʡ���d9���}P�����l�	м���	�0?lܔ3%#��96�Q(�3��fX$���4IiS@e�	�B�mAb�V�c#V4лo��.;�~[�����s�Vm�U7���~��e&�_��������ZQ$�����H�ˋ23��H^,hS9�!ӿ���K:W,¹{�Z�Rf���U��G�+�.�p
|a(�X��\�����9a�H1b'p3�l��e�b��F�6�9sS���mC�օ���[�@ �om���C��\�m��+�z��S����#��޳V_x*+�����]"��"����>����̤ns�B<�*,w�N�Kh�m���v�V�{iw�#�� �z�)������H�,�tk2d^�� 	��sc\���zȲ����p恨-x�JQ�Q!j��sx�;�צ �A�_�[�^7����U}#�����<��C�v �6�~[��XP�w�"�S�j�q��|UcGz̓�m�ew���.5UZ��u�������%��"L�ʨ���6�c�ϡ�UWۀ�A �]I��N��L�ֿ{�2%���
��#W����q"���W��m#�bg���������8@oY���E��q�/��e�\����d�]��ȍ����*�z/��O5qb���E�i8v��;������JS��&F�����("U� E�!�B�u��NO�ռ8���\��(�����~��5zXd��g
�Fb;���ݗ� Q�Cи�bT�mw�8jpb��&�'t�����
-�iuW�_vknH�{�O0�_0GXO��PCA]�W����kñ�C7�$1145����Rn�=�h)���O���(C��C�m��R�k@� :78��Mǜ7�I3s�>���_8��Һ7���x�)V8�F��YM��9�n7�<��ɏ{�al�^�K�Η��D_vҐKFq�J��ʈ�ؾ�,��GP ���%���F@�����]2�o��}�=��澋�( T��G��c*��r�Ϟ(:�g<��S�{`�BF�;ٚ�& �%.π���al��ծ�k|e�T�:�s'��	ey���1��\��t��É,�$�>'�M�Ioځ�Bj����Y��!�E ����՜����������$k��O�ɓm>�]�"� cn��[��
:��y5l
v!�!� �7`G��8Y��(���0���
e������4�.ZU���rI��/�R���f���?䯻Fٔaec�O��x�Pސ�U���u��|�������3JG�k!�g��# ��*v���s�{��+"��Ø��L�;�.�αS�*��l�B��N�:U=:Yg~�p"��+���x�e,��c)͂�Sw
X���t��4Ja�%�a+��?����� J�+�=KqQ�2��[7�kKD�O�8]��-@�8/H���EQ���(�\�L	7(`�b���H�G1Ƚyl�gU��I��bz|=s�>�5�t00J�z��
R���5!��
�k[���F܊�WY����f.�/iQ-�l�}�+-^iD	��� -��^%ޝ��ԅ4�U �7���gN��<<Y
�'��h�I�'�[9�C�ڠ��6x�2�YC#�<��4%����U����ZLi�!�F��`)k��6��p�+$��P��"����A�~�Z�yH��z�4!3/,�C�o��8<0�M
��F`��{������(��5�-�<�t]�ߓ�ϸ�_��Ni}��0���K|o�����9��7�����3���ճhm���KH;g�{���q�$�Ŝ��:1�,�����+|?9:��
�,�W` � �(Ww�,���D�:CR��P��?�ÛTl��	�%��R�⍂<��"|a��S�ÏL��ъeF�;6@N[�Y��X
�﹔���\���	�u��f�Љ�R��t�����Î�����م�V$ú���)��d?�,H�z���`n8b���4!oL��V��=D���=1�ލ6��u�e��G�I�_����e.�4�w������k�!�a�q_:�����co��(�'�Vg���fl���>�#ĀCr�΀�
���=#I��q�,��ma�5Ȩp����+7�6+0l���}tL�M_E�^�������!o`�	����l�ⷕ�LP�;5>p{���uV1�L�q�UN�$���o�\�ʮmEO��k�"�c�xY���F�r<�Uh�ٯQ`�}8S�K��C�(8�k����[V�%��A�4}�c����
2�����*�����Idm0�浕]��Dt�xoM��=F���"��$�r�.����h*R#
�����.^�����V<�S�F�E&k;/w����{Z�]FP��K�TXH"b�u˕8Q��T�UM�!�A+��e�cր���L;Q��}X8�0�i�/�@x|T�>�l�]`��kE���n~�)U3zN��#{uRy8�⁹�Ky�2��AH�y��i-��BވS �����ű@J~6�j�te`qw���3b
�/2������Զ��	[���7Og�ζ6,�C��=2������#�� �yJ�����N�TS:���:H��c��\�2���*��BB5E�K� F�n�E��<A���<r�8wě�r!��P�6 �`�,�>���F�%q��ż��v���	������������>���k	�"��ƻ���������6���w��{%��:?�zM'3����vԛ���AD����|����S��}|��Zs\w��՗���'�\k�$���㶱��恴���e��5�F���t0��_!�ej�*h���	�\2�m@S�w%��ʪ�S�2y���9 E+�����³J��N��rwϠ"�c���t�\�	��a����Z ��c�%UZ��m��6)��V%%yT�,	����;<�mɆ�v��ʗp
��6��@u��a$K�<;��r�@��4���3�k�VB�߾j������\@G@{�TZ�9'薂W_6'�>��D�a֗~}S��|Q�����7:�W.k�o�,���?�ԗ����0`�ʤȠ�'�L�}�3LQ%��X��Ge��k��{�$���8�D?8g�4��`ϵ?T#w�<��^"��7ߎ�?^L(Ql{�)ncdDB�Fh�b`�  �j0솱~�c^ӭH�:Q\Hc���8����'=i�P���>R@�"��J,����-��&��������Ng#�-�O�|I.�JiZ!�/[��N<@�3a��)zԪ-ی�?uq0����N�%]��da5��=�U�_ZAv�z�T�x
-�g=R�ڞ�)�������P�^ԥDE�Z�w�Q����T������-��Lz��o��"�K:+6
^n���V$�&��i�7v�5p[1��b����q���7��F�T�N1g�E1���&��5�Ң8aä��GP��0)�)d���Yy�=?@=��1k�馒e��.�3�|E���Z���/D�lq ��;�쥸]ܯ\������ w>�w���;0��>=�� HՍ���ȹ)�	"�?��z=�Ϩ�nI��:�{P}Ȼ"�a~O�DetfD����=�Y���(�]+N���U0FT&o�����ⱚ0�e���L��Ly|?0�g�CG�sX����Ӕ�i3���av&5��@��P��uzD�Ufx�LeK�K?6��v���zV,>L��oK?�Y�w��m�z�NM]��;�Cf�ְv!�6ؚ\ی�3�'��-��Y�lb�������_�!�r=��ˇ?W ,���P�f���� 6�9W®�i�`b4[t�	5�vB����br��&g�:t�Y�;�V�n�"�����H�V�S��UߩΟ���r)�<����<����zEg��$���˱Y�\�P����t;	w`.z���ʸ�O�$0';��̀}�R��H�	
{����i����l`ᓎ�R}b�I"�~���Pع�GBo�l�e�ޑ��A�L�ރㄿ�ډ��k{j� ���%I���	?>fA�t1�I��Ү����H;�?HRޜVR݂G� \6�6���zsi��� v���t ����K#0$~D�C����L3C�&o� 瑦W-.�d�,��ou�_�v*�a��Y�]оb}pIJ
����;�F����m��$�:5D&a�>W?�$�w{Cc��n��&�ϊ���;�pL
F� ^���#��P\���B?�Kuˏ�ϣ������@�ߒ��m�u���Q%��'�w�����S3��+��ᆀn�<~���˛'V@܈�Kn����1QP�\I��}`��������g?Yx9��>�]���Gu��URĮ+d�D��}�׉Nxb!	9�<Ή͏�Ӭ�i�Aou7�쓊n�t}&�ܸL���⹊yr�Ç%(����7#�P'��BGSzظ)�Ԧu����?����:W	�Q��#[��C�O�Ҭ}�`s�@ĝ��
a"�:�Ԁ�_�{��H�a!p���_�$T�C^��� �0l���p��x�=|�gL�������J-h=��`�5�-k)�C�K� }<�����a��Ăap����_
Ggz"�]9����\ʦV����ҟ���~���A�hD�U
�*�ruC��N�V�T ��e�Y��;q��;tn�O�"�Iv|�:��K���f~
�i8��ޠK����sy�'�����@�����p�Q����sx�P��}s6���(�0��tL@���Wo�/��\Bik���.[�������{�:͑)��$�S���T�];���_ME85�v�v�4�0�A;�J;��Xj��^L:��lĬ�>�E�_0e �7NВq`�6����sm���_8�G�N�=ή��U��y9cݍ<	"dZ�%�ٜ�h�C����>A=�>�dԪ���U��D$�{�V1����(���j�oD6ʃ����Ǣm�1�]�H��'2���N�h�Ctj�46��b"3(��0p�GX��ZwSJ��3rq��{u
FF9�)2a���;�AY���1n�!SH�{bG!��^����8����Ӎ�.�@X%q���(��T�BJ�S��``вbGwb�Ĭ�z�
N8�y����덍��oD�z�_�IS�U���Ûm_c��\��b|�{g>���nk�����*Kg�u������V����u�Q%�%�mЀ��]�h�h�^����:M�(Ln�dUZu��Yo<U�>\ƛ�dM�K�e>S����D5���Va&cw�=n�?jjB��xUv9���N������L����k��t$���;��+�%_����X��M!�B	#T�E��h�/���Sμ������X1&��+k��h�N�F]�G�u�AȘ��șh��k\�K���s�B���C�˕>(퍊N��[:�Kw��e)��1��cuq	3�I���S�r��@�_�iWXZ�Y;�Z��sG�mc���b�f��K_�a�>�=�����T��L�ۍ��+��� �ќ�J��,Y��m*e���tsȈ/9�%��;{5R��ut�A�E��0��	�"սx��g�N*%���B�6d��2��(Mz�	�H<+1�A��Mjd�ۤ~��k�	5^y�^U�3�Z<��9 �9�vV*����b�?@2�6�}�O��%����9��T� ��n��z:�=�!~-�4�+zPK�XQRG����S}4JΌ���Y����}�^���0��}��b�1C�v�mi��(B�SO'<�b�*��6���[ʇ���^��&p�o�,C�(�\B*!���F��XbIE#���2����2��]h���#�ߝ��V%�������/�ȑ��2�\��u?�=]������zw��'W�چY�=���{K��#n*H�(�Ԛ ����֕�����l��{��yY�z�)�����<zM��j�V�h��\�T�ě嚳._����ך!�y�$<�U1�h��T����3u�?#��ϖ%dǟk���f��=@L�^Gd��E�����:|�X>冕�� ��e�B�:���(�O�ƺ���a>�{F�W�#P�/V�_�L+D��u6�J�5sM0�_'"$`��W�6fٙ�Ր
���6G�S�pb�G�~ws�p���/�Y���Z45�{����[ν������&�>b�?��>�K��:�[u�#��+$a�q����ӷ�
R����OE΢Sa�~'�Y�/Ox�X{�P���\��쿥�"Ua�W��f��A�� !���4xW�0��S�1�'Ts����r�a�	H
�H��8_lNy���w�SnJJ�F:"-�wș�xn�uim�<ôghӚ�O	��p���e�m�վ��]e�h�+K(��3D�:��)'ZW�}xy��&NPj�H�����ͯm�4r���ɕ��#���PUL��&k~��H������օ��z ��zh9:�#��"썳��gu���,������ Dkv�?p4�*���B��A1�5n��L��T!���4&�VZ7�U[�0�		�f�,�<��؝���*�����z=]��5�hQ\�8�Qu�������{��q��DL<T��U~1���Փ�6�<�q�){��߯➽��y>�!�#��܀�BRW����l�]����aDEU�n>�0SXn)�F
�.���Wߌ{`c�+,{�3� �wT#�^��F��:wk0s��l��˽��]��λ8\�� Qޥ���d��_�*�~�?c�*�n���%��>�<*�Os'���gC�_͚��C1�%�d΀y9�Fr'fG�B��n����G
,��:7ܟ�#�������-�D�r3&�������C���v��*��l�F��+Lڭ��;����֋�e�A�E\Ђd�R��r?tKGy��y)���edF�
�[�¦�1������«�\��O k�f��b��֐�^���Tǅ��;��݃��[���x���c���I��7��-S���4��ċ_ѿ�H=���TWk*�{�#SA`�u�MD�Yv2�P�C?&v��7��~
/z��9�Y��0����\,���QMbq�u�Z1��eW@!`R�O*ʹ�L��B�+X��&j���<-��z���!BF����8�Br�g�ۤ�&�rH�pp���z3�5����*��?9�kY��E��e�)������,����4��ef�h���Z�L�b$���:�g9��畅����j0 ��~�[��� c��e-�zK�bQ�	�R~>�
m�SW�����\ �C��<5>��(	�~���󌺷�I<�O��2Q�)Q��l`�hҶ/ e4�H�U�� )�(v�]E��[��(��y���x�3��3�A\b������]�������M��MA�|�g������X�-6�&�Z�a��Jᔫ�����R�E�t�U(d#��<��M8�0��"�I xN�玀����J�擆(�f�;���1�Q�
0�+�y��,��4!���E.-~�(Uݳ.�=Xy��=�����r��U�Q؟4x'(�dn&|��:�;D�2`<��-�1PI�ـ~~��)��	7��P왥>��:T�R�=&��/���*U��c�'z3�1H��/��*Jo�H��Wפ�P�Ϲ�k	/��^N��p��ҥoɢ���2e�����JE*gt����eYI��b�j�kձ��KK�9`��'��=(��
�r����T�٘�l$=�S��|D'5��Fq���!���(�����|]�ևm�Y��3a��!/�<jp������Q��!n���H[']��F���j�h��<������9��	��W���q�v'�4�J�Z�b��w!w}��\
d\��E��ؕ�;��!#�>=����|�E,;��o�z7٤�$��x��f��_5^��M ��:�l����QTͿ_ٚͅ�;�T+A���qG=����*�:8�d��8��bR2zr�*�}G>{G3�� �hK�1l�c`,�ض�`����_��9���
q�#��a�c7�P�	UYw�����{EߘmB̄><V�_�f�uC�A�]�i��T�y ��:`����b9�	�V���8;�q�W2LQ��:⑞�6�^rN�1lD�.�r�y�Ԅ��yQy!S􆭇B�70�����L\m�
[�(� D̓7�[r�\���N��}&�@��>�9m��9�j�c��	S$���$f4�����w\+�-�����ժ-���{�o�&M�}��8�QA�XY�����p��EX�G�«�;��|���u[d��/>�aߧ��:��U-t� ��R�ܗP"{r���-l6229=�p����ی����z>�f7�l�2�D���&���c�����C�]�c�Qcs�(���z�:���'Kw�ر'J,�"@+�LJ'���7���6��M���$;� �MR��y�;8��L��4JA����;#��-���x�������D���Kq3w�ǉ $�N���B;=��)�3�v�/5���r7�2/C���~h�t(vW���Ͼ63�c�&6���� w�"cU���k.���ÿh���v�i!�A~6�zF�]W���N�Y'e�ܔf`�gxK`���g��C��{��G�E����׼G�J��|�B����ؒ=�a$��z�%���\܈����y��x�	�IF���g��LSQ�W�zH��	n���%��I�l.�(Yi�5.���Ƅ-�����|:aS���Ya���4|g��nGɱ��4�I�Nu�ƤI[�6�!P 5�3R�
���Xs�(�qz]_�t~g��I��j��]�Ú�B=؉�0ܻ�)����B�{��m�7�T�2��C4�%�ח/
�����@�=�]��w��O�R"A��d�k�l�n�=oح+��5��8��{��Z����$®����$��vQ�Á �q�j�=j������̊�-�8�@M�x�Y�'�vew=�K8��:����o����T�n�E��	{�Y�ؤs��\9�?�aU娦�]
����D�T�	?80��\�Z��hH� jj��?�?��C����9uglM�u��$>ڽҼ �S6�-��٬P�E �(a�����[?�ch�y)�=h�tu$��I�H6Z���kV�(�_MEHİdUo���D7	�2����$��b�^�^�����R>}�-Z	����;���{P�i�>a=�>R��3�0F������Ê:7�$#�dUd
�?D�y�H�/��w�L̈́�<~��0�.Q'�c��H)v&�X�[Kb)��O�<��p��ZfKN� UPT��
X�;�}s�qs#�`q�-(FB�~.1�<� \4c-��x�̉�@G���{|�3u�`�W��<V�Qq��^a\+(=2��D��Cz3�hh �b1I^��$?�̐�!o�I�԰��	���O��&���ds$_�f�`ϣ�L�D��J�!���Ĵݭ}_K����|Ȳ0�(���F���9m ��8��{���EA���譝I��GN7.
SׇN�9�*���3J�8���e`6����%C���]�ؖV�d550�c2Kv#ե#�(ۏ�t�Rpb:�o;�{ˠ��,������AM�?�}�Cc��A��4y�ͮM��y�!z���-�(�vч����W�T�V-l��N�\��qόąsA��pN7�.<��6��v�,����c�G���BSƌh[�"Ƙ�f��r����d��v���K����O�a(,X�T�Ջ�Q�iî�3���'-k��6ف�T���SkFK�H1�5����R됈�X˞٢�����"�����A��D�s75 �7�ڳ��!Upj��zB4���"���$��Nl��$k#>���)�{E|,����Dl�%��u�SP=�3�0������/u�D��@�/w���g �}e��o}w�o��8d��]eB񷚸�w����[c�H+�y>���`[�����]��M�wt���Ӣ5;w���us�%�b�B����,��Nh��<A�i#Fp
Tӷ)wI�^�R)zM�l?����b��s�Hy�u垠.���<HPA����cWКf�M�v�^��V	X��{������@�f���n�1b��~N��GYU�
� �9-�Ĵ�~�&c|�ø��R�붴�bE+�f��,Ri)�C2��	�����3�������i�����K�>��\����ӯ
�nu?�"J����h�zL���s��8��dQ�;g@��hx_Q�Mkl1C�s�Ir%�Cqb��B7K��za6�B�����:��?S�Ѹ�BH���=�g�gRm�Ya������oxgRlJ��r`��?�'��!Ќ6L*!����.���Z�]��\av���H�;��h��XPO�6�PO�)w�Ԝ�(�#U�@"=p�j����K����~�;gD�a�N��OJ���?\�U$�Hz��,��YyS�?m�eA�T�������(�S���6B'20'}m1�z˸�>�ƹN�(�2�	Ҿ�,�i:��d�~����	�o$� �\[�V/tk���	�P�(۫}t3XO�Ww������g�%��랏����R o�����O+���|@��V�ս�f�����X�N^d0��b:Ox�k%��,�����6M�P�]ʼÈ�Ts5����D���B�<�C�KѢ�e�P����/�W`t}鈖�4����X�9�i�#p�>���O�����$����1��I�z;�$�a�cX����|ѷI)���N	X�4i�#��0Z�x@Mx���l��o��[�@�t��ir��{G��b�TN��T�X��tY�P�e�}�y���k��/��RE�w<��c��Mt�c.ԧ|h^S�c�ޒ�[�`k���/��-2NVU�Ȭb����!��l���7���_�|�y,/��&)E��T�{�ُ�]����ǡ���s��V�m4D%lI�B�����6��g���!���E#v��׶;�{��m�+ָ��1��r9+?b���YJ���B�[#�J��.�^���4� �Df�n���I����˰�R׫�Z`�d�Gm��7m��h?�Z
!��W���׋��d;�x�\s��0T�W�K������z�o�4�����8�e�p�ͥ�����/���:,3�d��l�4�k����ҵwsqv?���殞F(
o��e{���Y6�2���zx�	�£z;�8n�֩9E��o��!;�wF���j��l�P`�g�-8��ϑ�Ӏ*WT'�5F����Mg���y}(��d�ѐZ�b���Xy&�s�SO�"8�����C2U��Q�8�=����_?�%؇+(��*x�z<<�8�K+��F�d�AzF'ahy)��tbin����M�'�fbM �C�} ��P��ԵbӓGx�DGc�~�2H�V.����t�.�
L�1���p�m���NW�j��'Yo�>Bӵ�� �*)gK9�����������������yP�1��� �����j�e���E�^���l�i>k�z�J8B̘ۛ��W7i�׉Lg�+������n��C�������_����TD8����}/�!J<�����R�:��#y,�E�%��E����/�G �:(7CO,��������"�zr��G,��TL!�k��1^�L:�����@0Xt��0�e��h,�X�)��gI QZ�"e��u�v�`���5A��|{%^�_p�����oe�0f�T9v�F᪭���<�5���X�!%=m.!��y�Sx��LE���_�ބ���ϣ\��,�h�H�x���ZL���2�����}��i�V��.�R�x
a,L�Ǘ�F�ly���'���&v��B�O?�Ƒ�eT��?k�)G�Җ{�$�8;
(6g��.c�^l-�+��DQ��
��o�o�pcH�:3�}��c�S���|-��E����բ7q�)��Ǚ[��ӰDg7���4�`�L���J��j<���` �..��
�/*r̅���m�z�GA-�Ҧۖ��a!v5�4�r����������9ԅ�#���b�� `�PU��J^-��C�|�|�2�m�3|w	h( ژuRM�$0��s~�/|�I4�i ;5|�([�����EtBSN1�;ݨ*���G��[w�����YA����������KP���Ob��i���sk`����qV�<?�cr㠇�*S������w4L �g=��6�#1���C���	vH-�
�ui�(�0	W�6(j�䏌��A�I�gK��M��LB6v�u�_��}�<mV��~�?���f�޹/:��|ฯ`���w� �G�E�/w���q���-���a���T�.r*t���A"�E��[���}�}q$�q��&�\���;�!�Ҹ3�aW�Fy���q&~��Wȥ�lg��Ψ)�+�Z�V!����os�>��6�|�������"�%�i��*=G��?�4~f������\C�\Ƒ��]T�������Ԝ�E^��]��R�fil��̰�>Xr�|"M�ð4�ܭaqE�~8�'X%����֪�Q�ww�~ŕ4��t��R���*ojo4�Kt���A.�3�Ֆ���~�fI����c���
������5m�)B�wrJi7��
��~?���c�x��:�������i��Ф:���J�l����B�}}6�%�s�NSW����ѡ���㜃���1S�%�^���)�>)��6��p��x�8����"iǐp�"������K�,��_��֋	��19�u��H���8@���K׆hn�:��`����@����6�u�9��֢9�6��#��VyV�c��Y�{����o=12j�� I d��!��w�f�)M���ea����u�sUr�2?�?�1Z5g$g��	�4�aೆfl�R48�<�]�CL���@9a���~H����}��m��-�>X3ЃV�ia}N�$/ɲ��)��z���������E���F�o�qS�pf�r�l�� 3fsBdE�ފ����(�k��{���F��b��{9��k�b����
`J��bx��Dӷ��s����Q�:�O����Q3`���>�<#ޞ��܉&O�J�\��"tl��&Xy��������9��8�5���n��'��`��)��䴀P���8��SJQ���vI����d�z��Bp��B¾�"Bm%fZ����M��g��JI֝ٯo)i�[�}4?v�P�T����A�b\ M�������*<ݮ���V���/�n6����.ña�����*�I�����ȋm�s�'I�ϤL�l'phG�\p�}��uf���_|�C�i�6w:"�gUdh�����e�gg�v��x�dY���u*��<r+p(�<ɞd�m�TG~��;.�B�Q��A}O�1��X*H?���Դ6�Pr�Q�V��z��n�L����v��sǄ@5]�G���F�2��D�������Y�?-�J)�n�M��M?q�=;Gh�=^]8w_���\S��|�\7_����<�l`)�v��ŉ'���A��n%[��QDgz/�e�ʀ�Ė2��3���Ս�C��P	��'ؔ�s���
Oȳ�c`��Ll�n\ea�Ü@�;���[�c�C��
��t0{��j�S����̇[����.��!��ztl�%�d��3D8�p a��Ab�N{**��b|�$S}Un^�$���W<g�1�CG�t�m��,*��JO�ߐu�0�`���EltB��:l�O�j�0�gt��yV� ����̸�)pW4I�[�J�c$�?��(����n`Zc����b2�8I�K'�xCU7-�D��F}k�����`M`�6��gb�{`�W^`q�[%�14�* �~�Kʔ�B�(��3A��	U�d;���UFxp�W�mTo�_#�d���=�Z�D�G�l�s ����c��ݫn�Lﰑ���y�{Qc��I���~B�1�zRI��Q.N�QUIB����,�|��gHYnP�ys��| I*��A�ka����3N����*ލ���ڦ����`�����O�e��|��C�f���j����r��Ӻ�&,��X~O['V:pѯ<�u
�0��+'��?�!�)�x<��@�
6�mZ���B�J"�a���
N�b�4��WR��#f0����5s��UA�͵MiI�%�c�b�$X���i��lU�r	0p�βC�(XP9��#7ȨL��5�	��¼��eɕ~:7���� ǁ�&�7�<SL5@z��Ȕ	��+g*8B��3�	��� ����������1��;nRt��nIy:qB�9�m޿��W�e�R�=��{��B�֚_7�+�õf��n,�z'~%u6y"m^!C��%��^�<�A���Z8;22:��Ao�XL�a/-|�3GT	kK7L\_g�����ѻ�<�CĀ���
w�v�}�[«�Q^">�pE_���LdU!_^���ae���h�oꗗ���N=�-�<��c�ZG�G(%�m>S�E�˭*9![K����Ċt�3g�2���	cK�FY� �����/�/{���_bF�t��A�����u��#hK�k�ںx�7��Jan��m�qc3�!`�N�M�XK>��n�߁!ND�ZW㴺��D�����*j�Ʋ�/�uA*4�~�\U0��c�"�&��[v��]f��B@�;����@BZ�~ck2�^�Y\�z�usDV���6��#�Yw�!\`��Y��$���]G���(s�I�WI�Ţ03F,��d@
�ש]�@ 
 ї���2����y:�i6�ϕܢ֎)D����i���������Q�o�/-{����(fA\�D���۞hR(��$����Y�w5<�K� r{1���������!��
XD8�G�9� ��<=�c�&F�L�ƹ��y�7�BZ��2F�pR����K���v�c�#;�BAzӲ4�Qӝ8B�;�Hc��M���?v+�����%�_O�!�����3���&��9hf]F׶r���`Y|���p��P8�Bð�!4>��%#E���C�a{2����whP��Mm[M�2S�ٖX��`�C㌺�^=&QkF�u �����#�w���2{D�'�(�9+�Ïa�Uu�Bl�y�M��@�d�1X��\�7YX�#��t._�9_�=~H�=:�0���<�=�kEc��כh@�'�M�'�&��	�+u �tȄ3-�ɒ*]��QK�'?.��|�-i�D�x� ��$'dr"� ��[�>3-W����x���vO�g�˫YLD��E�Z�45t�e�d�N�Ű0�f��HKJ�T��l���A�Ԡ�:d�F��X��d����e7q�w#Jy�:L�<[���O��a�,�Q�'�i��cB�Al�!a��/A��.��d�ԩ=G=��^24�T��:�N��Z�qy��K�'��(첿T�:�C'��!5a:����H�a���p�s��q�
��d�܎�P#�Q�~s��& ��bcrɤ��]��G����O��)I/`���L9{@�]Ek��:%ji1З�5l$g�)�C� �O;���d|��:�t�N8�I�\�e��s�p&����!~�� >xg��*M
���䔐�X��/�%xK���F�"mU~<�M��qx�ɚ�.W��z�,�${�nP����t��a�5�,�%����'�:���H�t��6M"Lt%���c�vO;�p �#G(V�<�F��Q��[ٍ�rE�"'$�+cj�y������� P�<Gy��*;lƮ���L�4I@�<���̱�{��S���ae{Kv&)FueZ �K��g��B�wz����E�˴�����}\:)Y�~���v ���`BT5_��9��L�^*#V+�/�HI
w"I:;ڟ�`�(4Ǣm�V�`L/�^1�U�Ka��W�zOw����7�9��C�_�D���+�����P����`�;��AO�{NxN�+ٗ{�z-n}������P�D~����^ �x��QA�衇(�Z�D�U��uiko|�P@�:O�挢.��ڢ��oJ�ӂ$�<���JL���6���fu���}����ЭMi���v�[^��[��|�y�C�^w���Ss#�#��k�]pOtm���q�$��@��WA!	�~ʛ�Y($�Y[L��2��"�84�b"�]�|N��uy�e)x��)S8�<�v���g����-`�|����*t*9øu���ab�@Z���)��^�у�'�UO� ��.)�2�/�n`,!�${9K:��4!2-`:翬��&�!��P̨P8#	�G��3
������n��-�P	��oUsaa~|�K>_Zʟ}塛�Q�~9��8�Za�z�9���C��kb[��K�e�G��`p�(��h�uң�*1J{�C(��]9A�
RIQ�~W�y��֪�D ,~Ȧ�XIs0ޕ��z��0��(�^�7�{A��j������m��g�p���s1��݇����O��ɠ��w�2ӼJd� �=C����9I��[��}��ƌ�ݣ����0J��?T�`�������O��GL�����B����S��p�=�ۀ�	�ׅ�3p��j�æ���+�4��KŞ�c�����NK4�V���I��l���}֚>�������LS&�b��;�z���6�7MaT��O�Ճ���6���;��V/e��TV�P��<���� џ�1g�U��S�䘷V@+�C�'O�I�6:�r\���Y���������Ʒ��q�@���l���3�s� �OȠe�i��I��?I��Zm������8�
��/9\��j�����xY�����5³ꁞ��ݑX�+J}����{�gޢFx.���+�DG<zr��Ozv	#ү�"�Y8�+Y_�����|��C�� ��ߑt��i���-~�3yJ[�k�b����k�k6�������O�(��<9`r�1~�њ�Q��ҏ /.�?^�؄)�`6� Q3Gd#(�6��ׂ k�҃�
��{�>��܎�;	Z�I�v��6Ň]ٝex�vM)����w���*#ɵ~�~ .�t�e��J�*��I�xu]V;���o��vAt�!��|���q�b��ƒ��i7fe`�Ug};,uU�3�v��!͇�@
�zM`z�"�ʪQ��F�~���Ê#�� �Wiy�G��(F�a]�l�`4NG�J�l�oQnr(փ�H�~���I�<��"B�}��Z)m�@���V�W���R���v�lA����K�Ō�7�Dt�1�Va������@h��莡�(|�89E>�KT��Q�g�Hk𫏬�3p�
��G�|q���}����WIޞ>4N��H��4u��7�_MO��5���ղ:a0���T��UJ�V�.�Q���Ь�^����ˮ=n�;�[/Ex]u�I�?�k�WK�}Yk��$DoK�����&nA	�C�q[H���g3�* !g-@��"���yloM���P��k�,�)�h�p��B��Li�%��(=8�)�֋GB����?��լ���G�Qa`x��c��>e�,�ɔ��>��$��,�}J���A�U9��(�1Z���4���4G�|:?�$�/p}`/3�]}�S�ױƞ� �¡��XꗇV��B��9jA�d铵��V���A$qcn5:��l���~�Wt�rӱ�bt�6M����K[�,�zT0�;7���I䧽=d��T�[�\�nF?C'	Ez�8��g��#���Ob�U��4���W��|P&�Z�{a�x |�'�Zt�?,�|ޝv4d��῾!�ت�[�Ƶ�cI㎋!����;��H�!vew��<:ZW�`�/-�2V÷�s�R������P"w��~�z�C�~
�$�te��:��|���T���f?�`�\AZ���% ^���#���𾬆{�R�T4i��ʜ�$�'}j!~l}rfgr�;�}D�ׅ?0B����M�{�v67#Ub��S
�,����|�@��(뽄��]pQ�M��-	�mo���n�������t�ֈa2т��Kn=G��X������F.X�,眛���s�*gT��i�� 0�U�J�t'�>���'�:� .R/Xvа{�!t�ʷ��dj��G'�5������.���a�W����ּ�ew����C>`va�gg�+�y���r���4�}Ƈ��cs�U���Ah�{(d�j�#��l�s����rB�_��!���'A�A�R��^uI圜���M�����R�6G��&��-����}R%#�\�$�{��ͧq���$	&=߱���/`'�V	'=�f��@R���r���@g"�{�K&_b���B��=���I��:Y�bJ�S{c��qRP��q��YF��+�r���ӖF����x�Q7��>w��W���jJv�j��gC(%�lBy�X�W[>�A�U�`/�#�Y�����0W���6������}����`�_B��G!��n7��~%L��Hȫ��ht�g��6�C�7�<�B������6h�'GP��,�&9��n�S� ���PY�?Tn��%�l,�3z�V�;M��CJ2��T*X�����Q������Ա�D;��(���j�d��Ĳw��zik���I*J��W����䟮{5?��o�n6�L�q=`/kEe,�1�N:���v�xP�$Gn:�x�?�#����l�@��ݞ�Q6�{��RUs^i��x�Rd�y�=HUr����ђO��/	�>X��+��@�6_%?ر�gp�Ч��R��w�}v�D�s��ȰPܒ��3-S������p7����賓]����[�vWh�r�!�y"T��͗��2��T��4��匪G�mq;w̡����{Z�_�f�%S�ZQ"JnbB�L�I]H)ˏ_
0�X��T�[H��8v�zz3�^'�E���P�^�c��?����u[h��j��H������2�G��n�O�sOWJиr�7���GZ��D&ozL�wׯ�U-��7�v�v1�q��QS:>�j����-� �2�.�Ћ����<��r��tj�l�!��wx֭;N�~i6�kH��Q�,�܋9�zn98^��\��� ���._�s���hm���eu~ݓ�Ӹ~� _0 5d�.�����(C�u��}�c���ӻ!�F�itN����6SU�w�%?��Y+밴��g���B"�?"���S�I�g���3��d�r�̱�^�zq H=e�&������s��-_�3e�ʇ��)V�o����\׸���ߓT��� �9�ԇA୲�1o�8E����k'�'޶1#d�5.�<��
˺��T�� ��#:z+���fzE������T
Ey��6���,�l��?�0�����A2���㿺�R]�j����6�v����u�u'局��XT��i��D�G�S!��S I*ߤ�N $څ���BS*xW����9C� ea7�%E���5d[:�]�/g�JV�c�=~v�0YNW����5r�4*�E�;��}�X"L��{���U���{e� �V�r��#p2��*�E��x-� v#�N�'DDE���������Ռ���>sF��b���Z!�=�~ɨ�9B��!���5�GrGì�/��m�}�,�	ύ�e�����v��|�oI7�6�������>���O;,'sq	$��_� 䞎���%�X��B]ЇS?��0R��}w��$�pf9`K��EH��11��x�$yS��`{~��a��cMU"e�U6�>��eN; y�h�t��L��k�����YG��	���K����#�L�x⼘E.j��wT�eӛ��5]x�,y�^����?�B��mz�)��?����=ED"��W�^��}=�r��A��9�I8�J� ~B��-��c�,D*�Z��w��V�T� [܇H>�5:P��
�gH+�e��<�c�p2Mesom\ J=?��8�58m B����z�j2�0��l��D��!����k�կ�L��3(()e��=�k�/��}@Z�j�l�CVW�X�Uh%�I��+?������� ���f!��e�	]E�{J2���L&�	Z�$�����e����ߖz�������w�\�s��������˚�K[�3��A�E8� ?�jr����}�� �/{w���s_wR: ��X�����0�f|k2S�����:����7g���ʈ�!��m�U�*���T�:�'%�i�gX��'�m ��+.�"ʝ#�P�w=&o~�L䝰`�[�Wg �"�B��1�A�PsF�#�pb���&.H�٫Vj�R�a�S6M�	�Ry�� ���I���bC�,*1έ�2�P�'Bl	�Ƹ!�|)j^A�ʲh�BM���L��y����6���J=��T�f�W�Z1VMF��2��;�����aʳ��qȚ�	��Р藙T\�x��efGOٳP��M��.�����S#_���_a�.����d�����M9J�N!�{.�ǸZ�Z��v�t��$�e��y)�8�6X�Bz���!���k"m��/~�S͍��-�l9ͱ��� �τ�C@h�[��ŏ
��J�GP��o����z��vZ��@����F�^��Z�I��|���ؑe�uB��*�CK`���)���S��f�P������*�ѯ��݋<���n����1��Z���f�	�b����ąD'�� ���bj�&�Kh$�7&�kX+[�P�C���)^�KC�=���>�lB����[��/D/����f�BO�kx���Oo*�G~T��Z����J݌�߿:-N.o�-�R��}����4(W1}�y8�!��Cg�&���%�}�'�AS�n��n:� *�uoW�3S��Hʮ&q��u)'�����w/(DkԪ�^@���+3m����51sGjZ�[x42����t�}▗^��֍-L:���L��9��w{!A�:����ҫA*����|���(?~� tz�$.�!��,�je��Y��2��窰�6�6���6��	-�k�U��
'T��N�0o޶zK�0.�=�8ql�k���߶�9\���֩�8�Y��)a9�aq�|�����>I�{��)H��.�t�|�>����˃�c�]-��A%Q*��Tg���챰ԠKo��fJ��.�2�e;2o��N�F3,ܣ4����UQ1Nk-u~U��^��l��c-qi��=�����/��yL��kӁ)��:F�m��:%!%�9�+؏��K.cG�Q���_�]�WU�s ���8�C�l�t�	��=���]�#��U+x��t���Ѻl��|�]�W������,��8��8`f���͑>EČ���M�t��q����dO���4�f�g\�_��\;dN��z�j/U0�fyUڹ	Ј0KƦ�_gX�{r6��q[�rb��?b��ݕJ���5���^��#˂��^.j
|?in�i��`�����֬=zdr7�!JF�ÔP	�H���׭���[�A>�3�ʞFB?�%�? ��]��QV�3��h]�����	�4f��l'A�]�̵��7_Zw.��������d֟'���;���$@'��/�f�Q�`I��Nx�0�"�6������d��3+3�<�^��e�#�ݺ�����#�7b{H�w VlX'����YԬ�p�F��c�R(�Hs���&�r�²�����I�����~UV�tST讀�M���s,K�4��j���B���(B#��q@�'�����K�d�ef,��B�9sF�iv��|���r����U��!y��8��O5!
�I���"g��t'��̦7��|�
X�����B^�S���!�`�➸���)Y�����Ș���q�Ag<{~�v3�q�}mF���D�j_9��ݵԤ ��#�W��R^� �Y����|��V�J R� �L4SI�j�\9�Y����3�j�lx����{	�p�d4��-�쀍!U'<I-N�{祙E�ߗ��fg�JQ��&C>�b�W���^<yqV�׌o,24hL��pRAy����q�qn�f0�X�c|���aj�4{jq��6Z�9@]<�S�"e�D�W�~D7pmFAVn�#e#���A�6�.䠾�PmG�b�N���b#�5!!���YqUZ����5Bj��ԉ4?)��ܦ-�6P""�U��ګ-&�-Re���t0I� &�S��&)�VE�wyd��e�_R_<��}�f("���_q͠��^8G��ܞ�Z����`��膝�d�'�6��A0�[B��d-%N����М�����Φ�������-Gm�����c�Hፚ��~��+�,bKGw�>�ǌ�-�+�J�({C������2���!���"�[�7�ᤏ�g�����s��Y�G�ⷈ��
��k����nU�0���/ֽ�%\JF��yl��L( ���;A����A����.)����߀��AobVt@�2M�C1�Ӹ:b\�_�Mva,ʖcD�XĞ�5�ˮ01#�>/��h��$-���6qKu�af�oH����������$M9��+��qQ�
.�����::�uifS2�fUԪ�����V������Fb��� ���3��V,��}��"Fs��H�W�j�(nb�K��5�O2<fZ�����Jz��<��X$��p
Lf��������g�:���GàHvW/��=K��8#z��۷T��Cɐ�:�$�7q�*V��S?�C��ޔ8�"I���΂Ό$�}�0ў�d����S�'���N�P ,7<--��fp~�erҷ��ؒ�ȼ��9Nq�|+6�����LzR+����G&�6ـ�h��4_h*��de˓E}=/�qjcx'���"�~��,f�@;�!k��V$�ܟ���@�����o��^��[\h�ޅ�Uj�E]w�g�\A�̡N��/0DZx�r�5��N:)<"���8�A:�O���0֔"d����	 �N0^[�j�b��j�'���z�T��lt�s����l�A1G"�C0ie�'�&��p����{��m�J�[����
�������EԖ��I!/������m�7W���M��$��V�S�Ο�Yk;��Д ��%��g��e#y�`�x�J�ke�� ��襥�|�Q�!�d��ll'�.YX�[z���u������o	�/��D���o�
��3=��4U����2xp��5��='~D#�%�����+�����3��95M�IH�Um�Z2��8��3���SIE{�rH��,6���4�*1ԛ�|I��;[ҚȖ�i�r�c���P�1�f1~�P��?|Ƥ�g�gl�����l���׹��TA��ytN)b&���0k!��y�PMSj�4��i����h�0jcFH����4������E��G�\��v�Ȕ#�a�����t�Q�� �F�����0
sX��6R����!�5�*��:U�B�SĄP*��},7)��{��ce9I���I8ϰ����%�̴�H�4���o#�4�ԷHw�Jlg��~5F+8��k7���s^�Pa����*�=��ٕ�DSD	���jF�'��.��J�S�B���t�J����3����d&�-���#e�?��ʒn�V��E�ZѡT���?~�˂��~T��-���}�d{��ԷH~�{���n)q����w4v+�?5
�A���SU���:����UͨEv8�����Đ�k�x�@�Z�sq-�F��Y��h��=�g�#8�#Y$��<�zp�+vw�mGj%U��<��}�0"��~!I�ф"���fbuGی
'�3nQ�����-��>�q
�S�<�y<��&�Qӝ}Y�&���܉�LY����+�`>ts����U�Bҕ�	�&�r'�tja� �����ZA��a��>"�^�D�7rB�Ð."�-�#�Lv��o	���Ȱ�̳2�1�V���_����(�U43��	����{�i����@.�S�O����A�Pwڃ1Wb���Jm�#�?ir� ����,�/?@hg�8;����_�<x��ln��Te#���|QqD��r7�^_���6��(��t�5�f���[|��,��z&+C숮�``a��������h@�N�G�D����K؊�����?8�X�o-�tb�	U�C�]��av��M��@	7x��Ѫ�Y(���95���΄R����2DQl ZM*p��Tyd/�)�吟 ��#�r;e�V$l&�'�`�k�~�I�忕�,��9*)���� �����k��	8Mc�#�?E��'��Ǹpf[(��Vx �S�`��1�R�ݗ�:�v�Z_�0�  GGL�*��t�e��&Wa���&+�I�N�ҡ�&�a�B`6h�.��D�����Z���	T��I�Y2,�kb��K_ͣז�8��漊�^u0G�Q�[	��%�i����f _'�<��ՍK�����Zs@婄RA� X@��)pS�3��Aw��$g��ܩi�RDSuf���"C�՟L�E��"̵��W��V�:.A�C����nUb�yr\C@�x�@�	-��&}�%<�u]&h�'e
U��Y�]��hJ\(����1��)��s,�}�:�.�����-f�w�'ۧ�U��l}֖�	��bO��������ګ�	U/��Ga����D�.�k6	��Ht����+��ڵ��7(|�����5�����5���K�'q�\��=��JW���+�^ݒ3N ����P��	�M���t�=@����[[deP�h~�0]�3�d>Ngm^�᲻ס�%4��e�j�ՁU%���#��L�6�o�c0|�LY�*�8qqĤ����>��������z�C;6�ToͼDj�VL�+�����B �b!9�A�bQ����;�'��}aSdڃ�KL����/��7K��ؗS�BH�q�LQ��t���}��5n���i�M��^W%�H���L7KU����O+)u׃'��?�B�Tv� k��a���T�{2����G��.�Ŏ��]�*�$c:�1�U$���p���1���zK>�&�<핎j�qWěU�F쳐;g8��s8T�2�ϐ��c�hD����b TZ{2Z��sK�jy
���H���8u!���
�Ė)�;�j���-(�rSoΦ'z�ѯ"? �>z���q�=�@i����J�3rg|���7g��p찖��������t��"����;.�,����[��FE ��~�j𭉜���¨X �@7�d~bq�!@g�*��?b����Z;5b�,�Cݗ���Ti�o篧h¸.��&�Ƥe!+��j�W�������qɱbG�b�g!R��@$t����ŏ��`d���3���H-�*o��PE(�d�gW�;t	�7�rP����F�lF��hV���"mĎM?�H˫��1+g?D�?��*��m�+�_��J���Q<檙1y�-o6�]6P��T8����E����v�?wb���{54Lw�Z����HI2�h��l%E=�>.���>�V���+�KnWo�d�����l�@�o����$�&ܻ�1�T��R�I�]�cǇU�<~��^�@8���k����5�ǳ���|%�>O��J ����y��HM�h���"N3��[���s/�ViW�tW�e���;��F@QNi}C�	V��jI�c��U<����#�"�t��>2h�Plj��9�vǞ�mڲ�R$mZU#�.���A,�L��n�֯<���5̓���.�Ցv�H�f��Cbkj=�&b�<$�{Շ��.71�������Nz�-j��9�FXYJ[��nip-h� �v�xO�R"p�������ȚH4��Y��n�9��u�`��g�1 ��L����#�Zr>���o�Ɨ�M���R>
,D{K��@]e��{މ���^[6�sFo�NbCP��(��u��M�~xc�Y�C�A2��;�0�O���F�I�5]�����1���>0�#UG�AQ+��ӇLA	B@bӿ��f��5<�U������P,z�bkz���&�緕�Isp$�9w�3�_G4W&�ң��h��(kbz�yϸ��g�W�5q�'ú�}�P�s�dZ�C[Ł}�U0s��mM��"&z�����HA�ʸuV$��㪡m��NvŦ�]٦vJo�����wqh�b���k���)q�Ђ��eK��l�q�̳ L�(�=]��.�h� 䡝�h�z��x���o��u�Z*��fv������e��Y�����6}�.��AᘲԔ ܏U�
����]#�>b}E|���1o��kI`��� {>����;�����T�{�:�-{ЄPӑq�������MzO���k�q|�
�XS�;	R�DJ��'A�`�	Y��m ��@SvF#���P �o`h��>,-K,1����b�R6ay�2�;Z����v�
�O`0��1���n��5Y��s�:��wj��7�N)CO,��G#N�n�؞LI��o�#�����қ�޽���E�Y���IM���l$�`d��X�&��g�VbQo��$^;y&�]Ը��:�.M DG`%U��OD-����!��ԙ�R8�[[�����Q�~����^M��`���I������־4�%�ս�7��i��߽$zT��h��%	(F����qW��ہ��"�8�d��^�^�ѽo]Sv���XQ���q0�L�S���i�ӭ>���H��CFD�-x�]�@�����~�D�Q�Tt_�A�*�s�;U��B�B�����\��7�>���.jŋ�f@M�Nk܅ ����F�( ������e�y�����g����J/�$�.2rMb�z4���yY���e�hǮ�]WiSG�Y��ě�j�Ø���}�HGwgz��.��1��dZ7���sA'�$t��{_��8xV�TG�g�l��z	�1���`�*pY0��9�a�V�D�8�k �(װ������[�#Sn*wo�1Ӧ�]fTT�rv�O�����?�&D���t�Tcxr\���Gg�� �ΏwU1�d�	^�u_Q!yj�~�����U�R���ڽ����f����rd���?�{���	)ί�CC-UZRj�5::�L��#������YL+&�фk}=���ͿG�F�m�T�����������5N����/��5i�ٟ%b������v����4�9�w_�]�4xim�(<¢�4�̇��K�v[]0Ш]H�����d/�˸]�0.@�D%�\��R7����:Ν��)�kÿ�����n�S4���D8�su�E�G��ð����xjݛ�hOR�D����i�a~���zwxy��u^J22�T#�Pַ�fǰ� "��� L��+xy\�	IBd��^���h-c�:��F�R���w!�P'���ud�:+��uQ"K��)�i�Uei�	B�����D�Y�{�GZ���h��������e�n߶(��t��f$���7@�Z��W�ן���z4B��[�	IW��~��/�&�n:
4��pKX8i����?�����F��=���� �_�ԏ�>�>~�[�GeR��{�[�#@5����+��8*M-kX��B�8���z#�?�������#^�8f�.�p����}�$� ���\�hyPNd&΍���2<4,�^g�%���U�b����B��R�{7Qd�c���/�lβ�!#he����">�7�ۡK�5EY	���L4��nF�qVF��Y���a@W�Y5�Ib&O�Z@�~� ��N�[�����hK���egN�#���������]��,4|M��a٣^��"U8�4xx]��^���s�O[t9��բb��2�<1�H.|����1l���#����>���M%RYɉ�T����:�l@� �?����Y�RF8��]�oД�;��x�wX�6�8������E'��z{�]�%j�:�1󓋠R"|z�Ǻ��y	����8��P)�t�/���,Är�#a��pN��2r�ow|9�HD�ڦs-ܿ2P��vC���G���D��lW�z-�IW\ֆğ���C������KH1���gp���O �.�vx�t�A��̐̈�ՍK��s���z8���r�8+4�ˢ�a�D�~���^;�b"ƍ��D�U~���t.G#�;��[�>��Ѥ#��\�$�t�ₘ���~��<7��� ��k_���X�#�{�qf ������䪍i)2���|�qA6@����	����!t�~�q|X�6�o$x���{��|�/&_��3�d�^k~Z����	��4�	��O+�>��H������D���d�Ѿ�r��P�o��5E�-�.,؄	�N���B�^��*����k��|��D���ÍX�y�:�.��0�@����P���2�ׂU�kS5�Gf��H��C�o�@7N���T��k�0�����-r�sH� ��o����Ti���.��}(�gr�gզ�������=�����;\j��X�J�8z.)�`���	EZ�/�) W8	�u��$el7���S%>�����۫)ў���}6��U��O��>�6�f�5T��G��0V�B�t0i����r/Wh)8�Fg��%�f\�~~�P)�n/ڧ�R�┄]�jZrn	�"�Q���!����Yg�,mU��hK��P�5�j}%����|��,O���촏iN�N��p�?Q'K�W�,8�*C���&j␄/�Pq��j���BU��I�)����/=d�Ƿ
	U�b�\�N����̢"f�H�Nc5N%yf�y<@r��辰�ݸ'b�@�k�y-U�Jj�\�f�퟿��-�(^���S����w�候��츐���W�������=��*A'V��ٳDM̌`��T����"͝!�[d!�9���4�����|�^ �u����x�Q�:.�5�k�\��%�-���MP��?��"��_8�)5�����q�A����A�hV��̗傗߂]l��ϖ.D�N.�n]}�GE���5�n�ئ���>���/��iYB����L}���N!�@L�N��@�/KZi��{�e��J��c�hW��-��K_�=�׽$ԟ|HӠq*�t�6O�Y��b`��!1�4%��$J	�)*��v����6�"~���-w݈]�yfq�.��`3�K�����4"�����,�VXd���i��5��2G[�\P�󱕅�yK�o����c6!g�z��m��J��A��> ��xʔ�9�Ԍ���O��N�iÈ�q�ǥ��B�|)I7�p�y��X���ps~S�ی�����a�(E��T]��#m��?I�+#_�G�
��0�MJՄ��إg�m�l��A�PB9����z�p/�������Xz�u����D��)/�l������%6�9����]Cǎd�B?�+f�:�������V�� �)4\BP3!���õcaۙbi� �<�I�r}_6^�]��H�4��}����M�\6��X��f���<8�@@�"�$3��[��7��y�m�ʕF��-Y��)�������l9�v�S��Ӝ-l�G�l���@�ސ�|T�,����AhN�!��)��R��oI:�D���UՉ�p����W�v�W,�3�IRr�Ό� %��'n��I2�G�?*�]'j����Ȑ8�[x~1�X��;���x�ד�v�NI�V�[�$5����j��@t�n�Pţ���q~Aix ͺ}N��ZKc�W/\7�����tM:̿�)<g3�UF�E�;�q���+H�˔&��F:UL䇗�zO'���:Z�����%�O�8����0�b��JkH������cW�8#`ϴL��2q��m��~IA�l�9���J8�G���PGX�J�4 K��Ӟ�4q�Y7�8j+!��8ѯ[HR�:39\<z�9蕂k�Dϴ���I������L�#�m	�B,��8��ϟ�Qm��v b���C��s���#ü5v���&��i��l�2=Oo���H��6����G��M|��hT�	@�4Z���� �[��=�?�L�'/��5���<S�[�=���!܍K]C���B��4*K��G='�r^�U��]Qӓ��p���mk�v|��K���gu�@��Mu<�فV��q� �U5\ɻ|��sr/�"�hգ:����	ݑ��%�B�N�����'wb����5�1�����dd$�	�9�ct���O%Y��s u�T}$��/ޫ����(�f�������GX%,�̐���K����_������;؍!Y��Y��l��]�ŧ��.y�&�Aw��n��V|�ۏ��diS�|S��tG��,
������&�ad��H2K�ӓ���SYH�[�i��D9>+��z�V�8��恌1?v+ ZWeԁ�ƈ��bvS���W4.�s�B�25�-���CS�gJ����������O~�� ��h������*4�>����P�߁�P	�O�(������܍��T������I܊vɵ�{i3�?���eOC�4�k"?���
6J�`�Y�����w_�t��?4�wt�b���%����N�.��vC�6K }/���](�)4@�#Ey���$�-�b�;�g��:-ڧƧF@
�f�$�@��'�ؙ��Ү�"^��t঩��إ���o��PptC�5��Z~wO�ɬ�;K����i��<(W��N���������-�,$��%�������������i~�Ϲ.wԌ�a���ޫ 0O�i��>g�"�'^�3�7z͝�,��tS��Z���(�~�A�Vv�XbwXv^�8"'a�m��9�R5�m��B����%s���?�Z��V�)����'��:��5Xo ��#�]#�`��[Z��2�^��VҖ��*�v���0y�f�jK8�!L�͇x/k��*C��N�>���"ڋ�P��D
�/'�laOzM�1F���h�}�D��g�q�����=�/����bl)S�S;�(�\\t�Z�NdKi��N��]����B�;��^���V�z��W�w	B���V�L��f4}hM`7}�i����p��C�!R�Dv{k�����X�	W���7�BRi#�O�@y	x��4�$
�G��l^��c�P�V���0a,
�����N���B6���J3��_�"q(=Do��<;��$�c#�+�_�Tu��_�I��d"`{%��r���7HGb��J�@��Uivц�9� Ԅ�jK�f|='��ǵ���f=PƬ)��:{n�:�
qU�9���,���x���j�\-����3�ц�>��#u�u�Xh=QǨ��3�K�ab*�v3�RF�b��v</#c�pY��:{1ȩ��-�$���Dٲr�z�>��d.�LH^�kNŹ�9�a�|�q����N�G��b_m���Y�?�os��GՍy�[t����/"���PdHA_ڬ�_լq�E���hM����r/��w�n�-ӱ8��v6oA�朔��p�� �<�Y��ω�k��?psn���3p竤hґg����U�1LuD
�����k�꽝��LR�?�DG�Y��c`�u�$��J{��v^8��ȵK��h�61���[���M����}!"��$��ގ�b��,��ҵSRG#8�%K��jp+	�qH�S%���Q��B�w6��y�{���<m���oI({�����p�6�|^�y���(r�w��ӓ�Q�������s�?r��,00|��H0�*]^Z�*���h���,z|�)�C��y6�HƗgm���z�����܇�d���J?���겅��g㨛��y��]-YZ��ᘘ�<^+��B��j��_��z\�&�PKm��2*�f���RO� <l��e�
Q�X�o�)�8��������Vl�D�;�nU�k�Zja_�-ѥZ��]�������߽��AN萸pp����e^�������^��rEwc�U�<�/vF�1ճq�zh�>*�U��	Ps�,��'dwC��^��4"�I�Os{oK�[,���^Ƹ��yb��=� ƛ@B�2��#\R�U��ʂ��w2�6�(޹���ק�幞�����شC�L~j=���n�," �a~?m4�+0�M�L���Ȋ�L�r���R,�a�0oo�Q4�A�=}I��m�?�2�I������� ���Ū��$�q��l�=\�k���/|�0��{�;�S��翼7��Ow���^����$�+�S�vim.Rq�~|At��W�$���4Ԁ�lQ�x-��۽�����~d�2X���oa���jQ�����!�̤?6���O�S�6�p�kذNj�i�S�hH��ϑ��BY��P���������v�W���X�N�;��#f��Ή��]�0���V�&R`�J%7��fA�k�[�Y~Hm�_	�o�(̠�r�%mzr��z0.�OSuoS^����]�R���h��+ �H5m�jD4'h}+�7�NC�:,Sv+��׻	�7K���d4I_9h�|��CD&mǗ?�����`�إ��~�f�i�4��/CX巐���tB��e�T�AK�c���L�~(j����r/����N1�Fm Q9a	�Zg�y�rB�ꤩ[?C�>��Rp��c�ŏ(3U/���f��sdW���fǝ��8N1
��%��$g�Fa2�3��<����Ď+�fO�5��YGi@��ѷGҪr)��>��vԛ�pK�5_t;X���_��C��ւ�����*�+���[Z32���i��j��L�"�d2���Y�X{�F��Q�ӧ2��+H�V>��M؋=��a�}�Z�\���*qD_4>�[/�d�5��@�Gv�gBq.�-�����W��X�������*���ƚ�-��w�߅*R���֣0z6v���f�2*�>>�d�m��Ϸ�!Y��Y��_s�qty�F�6���v�����G�O��T���K︡�^�޳3��q&�kX��V;�Iԗ������Œ�tR�,j��^n��HZT��s�4Qlv!����lz늬<{;����2�Ɇyq�Mh���t�T�Μr-��\���9��c�����$�9uq�����XW��J�������L��Ť�m'�ޥ�سEU�R
� ���,+\�$�3*W��5`.J��b.K�#�yK�I�R���.ò���B�U�y�Q�*6�o�?� ��3	����L�����i^dTC��)�bW�\+a�\�,��ɫ�a�-�=§�}��\�Eʰ/�H1q��s�yHu��U���#�.3B#X�����E^E IA�u�t���ݎ*�w�`����C����R\�������� vH�Gǂ:g䩂�<����M,�:>ڕ|��ϸ����G����m��9D�9=�����C8�O���<�$
	kDC2t:�2��VCd��\)�o��d�K'��G���{vf}H۫4�gad#�h�Z���m�]f	�9�_��qH��E/�h�!���Fu��H��
��������הX��0�DA�G��N)�=ⵊ��O�2��Ũ�������p�
}�D�>v/����]1~�����+h�c�*���g���i�/�;�^F�܎2�jg��Z��3(��}ر ��Ӈ��9h��T5-T��v�[E��t��0��;[_�+���91�NO|��b�Wn��,i�&c�q��coP��5e���� ,u�XX�㠂 #�%�J0���V(�ͳ�[��^do*x\�����3Wk1*�:��ڌ���R.T�� �'��J������>_٬�>��my�a��-=������FV|���ʢs�Y�m����E)�0��X�w�l�<�菻���gO�F���l"3,���տ1�V�D�`K=���g���W#fl���'�.9Xd���Ý�f��Wi�/�u�$�H�)QW%4�P�!_��Eǯ�dY������Ì�Q�����$�N<�������%[#�6�P`��s3d-3���"��3�l�t,���pNt�.�n�ț'ٌy���=RM����L�P��܏��;�T�]W��yH��`K�����Z�q���Er��vU��G��GB������q7(�>u(��{�"L!��9 ��,��p�����z>Ե��%f�����)V�����eT��+ͤ0��#49c��-�"��Y���!�\�E��4��Ы�:5��G/ͮ�H8��9�F~#���0�l�d�_ �|��j]�+�A(�q����˟���m����?�AV) �Rx�j�E�(��w_ǋ�#W!"Qz��\�u~G\�}�Q���7�࠙��S��q��EQ��^xyeZB��ԝ���ǂ��B�����y�2~��p_mb�W�EnVۚ����ᶢS`�|ڛ��Q�]����'�Fnp[�Y�{"teG%�8th�~�Z�vԛp`�LLW-@�=��
�A���5�5�P���a֮��_#��� +��P��{�<��225���V7!���1�]D����o�Ml���9�%'HRN��{�K쇖]NK��8�uڦw�8{[��+֬H��W�Es4�c`h,<���Ǘ��'T�
�y�BWH�g��e����e�J	�=�dXh�L󅖹���%��=.snI��,�a ����)���&�%m�Y4g�#�"n��Ȭ6����g&��a[���b,��j��{�೏=��_㝧,�q��	�(`�ؑ�W:H@�f]<�y��!uߌ{�S8�N�-Nh���~�9��9�$P�o�_����67I�����q9�5�+���������0o�������1��3<�}��m:s�|9{mT�l,�V���T��s���u������-�ĳ��@�]P5%�iU�l�0�p1����$�`e�߂o
}��Ч�٤�^ZQ�O��8eE��_3�J,�!��$^Y*�����?�
áF�@�I�r\��c�20Z�������U��f3����3�i7��|Ms�p��u��`�i[��n����r��iƀQ'��<V�v&���y~Ƭv-)S�i�Ox�﬊�3Ie�1j�~�[��(|�&S,aY=N�)-��qxGk���|��*ِ.z�"�s�"i~~ԡ$w35V[� ��	��싦�{��k�W`=W�5�6�J@��9�mæ���*����둦�Į��u�f� �Pŉ�3��\k���vR@v�E����й��s�Y�g	�X����K;�v�k)���x�S �)*��e�b	���6�!�݄t��iLd70�7��ʹt��������e7�(v?� ڄ�%)��1&vK&��rt��+Ƶd϶.�W�/!^��/�R/�lߺ�ݫ}�lu��2(M��61�"
0��h�2���>�-����n&��,_��uo���爪9j�Єl	���ݝ���-��z�9�3[�J�!�Y�n��*)se ��0�C.N�Z��,�C����~��V��[ש+@p�w��<`�؂�r�A�rc��4g�I��:x����'6@Y�'2$��
*���# W��b2�B�[�3҈I�Ǚ�h��\Z9IU�:�&^��ݥ���?��G��/����,�v�^B�<M�ޜWWw�O��h7|X,�h�Ǹ��G���LXh?�ߐ��$��3/߫ct�~V"�#����:Ǘm�"�u4y^ib}�R�X����0��7�'X=t��W�jý=�w��k5F��"<�/l���^&2a��gP��HqnW=���t�z��������QCko�|y����(]?��)��WW���#Ԅ�V�&��C#�C�T���L����� ��m^{Mq��ͧq�#%qb�N�	��0�Ca!�_�����@`-OySob���ļ#ħ��Hi�gq���H�SFx��8R/jq��F�}�m|B�!����?)�+<��bH�8����5�Ɠ=#�{��h;��}a����Q���
%?z
�삥%����A0��>��u:�>���-&�oE*+����o>W�ʗ��:M=�u�X��%I}]|T�K�i�:�PN�.�^�4������=�����J���7݇���c��E�ތ�zH?/E�bĻU.k��:=�6l���dLoF�hv��H�3��{�����[QԲ˿�}C�L�ݥ�����
{��&#@�»��;0���c�0�O���'�.]�V1�i��OC�d\��b�a���n�{�#�	>��o�0��e����-4#�h�ΊY<i��	v�ƕ�G��1�\��Nh�PV����������u�jA�PR�����+�f���dM�6N�m�1��F�$;��}�G�t�$�v�*c���s�\�}�R�P3%��iQh��3b]F�����O�H���F`��u��s�#a�WL�	�3�X�T,��&-�T��6
̢c�����ʢ���؄B�5W�b	���q�B�m-S?�wC;����[D�>�1�:��PLW�o=b�s����s7/��ʔ$7�?�:mq�Y�i�A��f�|8�L�TMB)D���`�}=5�ZS��|R��V�7O*�g������ʳ_���N@�f)�n[h���j%�ehɩ�ݾj����MaX*b�5�U�C�c04[f�e�Z.Ps�ۖWC\&%�ߍ<̎�xT�Q=�	#J�hCn�R��kH��Gk�4�)�f�mWv�l����[�����(5�����)��T6�����l�}�~p��8&�(��5hE��H��Th���@��ѲT�f���� ��Ê�@A����!����[o�9�t�E�_�H��&߭3j�d%��k�֟���S�(��a�r
nfS-��]K
�V/3�]��LI.UWj�9)�|���/J����)|j�3����Qܿ4�d���� H�q1�Sˋ�� QA���=�H ��<=�;��*��Y��s3)1h^�e��Qzqm�y�Ͱ�Ώ�ˉ�bB��D�IzQ�fI���x��ƟS��W���w����Nw����&��!�?$ 䫇������-��=���<�>tUZD���(��p�����ê�h�R���}�J��Ҽb�8#5D���/La$@FOy�����J�Ļ��爈*˂$��(���G�87�ѻ�e�#W��Dؼ$x�+�d����z�4&�����49>��.|���!���)��o\�?Ɖ8*��{�$t�́�"�Zق�&�O%/���a8TH�~bo�
El٭���Ww�u�[@[�H��~��V��md}tY֝�AYcu�v&E����~�ӭD�:����\]7h���Zߠ�D�D=�r�	��?<ϐj���f>ndK�����z����T��+�
�c���<=����.�e
qiQ��H��
�;�P�G����2~��d�v@`$섥�߳����y��v07����"��݈�"�Q�~ɼJ�g#��H�4(a�N�z�]����HA����%oh"�/�(lS?pr��/yu��_5	�I�Q��E��^vP�������{�(͑r3�����+ٔI��|�$�
�/Ѧ F���fL˙�if�T)|I�P��FS�*s���M�^�]v6I澡x	�"ݽ�zA�>[��4����x#<y�&�U��T��JV�X�3%F�TƹGv��� 
gMR�۶c���i� �-ž?���n�G~]������:,��N��/��]mdaWtb���m͋M��[�?"nU^�	Btt����Xg䂒��˥^_IOl
�l��Q醅�ʧ�[ܵuI�r�~.�05D2����7����u2����*MC���*^��6#�|����oo�fz'}��Bk��3G��m������bV8#��d.��f^�:�P��Z���E����M�ܳ��k�=R�S$�%��n���,
u4�-:��Sz�q��?���H;��FL
n?m�.R�MV`�>�iqda~0���?����_�n,0�eB����hPx_@G유�g�XW$��%x���j���hW��r̈s���j4���#;e����,-��7�Ts�C�ʐ�;�%"��B�c��{c��^��!�r{�so �� �E��D����:R��B�c�:��\�d6wk4����w6E�Gf�tY;H;8�	�K��ŏ��=�Z#È]����,�	A��n4/�@����#R�� �Q�ȟ���U%�;��r4� �6�-��������_�<r�!�S]m�q4"ΒV-��ř�Y 6���g=�����V�³f��GJ��ʐ��V� �;��D����Cr%����^LJH������V���CRǈC���D�����(�Ё9G�p�߰l���������!aC5���O��P�0_=Uյ]3�_���� �>ë���k��:�Nu���r�ͱ�����쥱�b5n=8�[Y�Y�T��B/���>�Jq�V� �qz<::�.��$���ȴW�C4vz��R�MU�RE���E�"�Վ��s��r�<�@a ���+�r>�5u
K�9�s�$����Ʒ°}B�v���C������ݤ$����kH:�@ �Yt�=ZI� ^���D���;���0�5��j$�b�zfR�Q&��h�ɒM3�����J��;�>�T���S#e�F>���Ӳ�gt��g�`�X!_�]�M��w�Sx[���M�̀��{NWXJ s��T�XVn:g��h[Rh�y�Tj�(�=�wGHZ���b}�d[ZS<��r ��q�$�A��$���i͒��ȴS�#�܆���m�RJs�����ݴ<)JxK�sn�����F�z�����rf�w7'�ԓt�5�t�5�Eq�1��zR�L�q)\hqU���ܿS����ښVr��
fA�,C 6�B�f삅q*�oE+�<��*U�ꌋ3�i�Vm`�,mu;n����"�l�uuy����r
E��	���k�-�J��y_��8�Ϸ���F������++o[ʤ�Y���e�wx3������\v�͠�<�Hf��� �5�4�w��B��*@����<Nf�r1�;xq�ݏG�:�_�ą��^읲8&�C	�76.f��y�Sh�57��M��}Ol��T]~��֜>Փ ǁCe�t��_��	�n���	Ȑ�u������lF.�ҩt�Dm�R`����]�+�Y��ұ4�ZOVDw���Mz��ku�������%LL�Y�xբ>�A������C�b�~�'W��-v1�t�Ӧ�3���L��w���W���
	���*�"=�. OL�lDۆhI'�C�~C*��Qy�������,���*���(�=���K 4�^[��}�BH�qrK-�٨����|f���A�.d�@(�_��'`;_�.N �>h!����}�Y��1s��UR/�.�3���ҊrV-�mco���Hq#�R��dy�[��v/���z?�B{��fg���R�	Q>vt	���֬�B��Y�jg!ыD���ܸ��|�Y�`��s`�s��Ϳ��j�䕎�c�J���-� -����D�Gc��μ)�W�WA)�Ta{�Gs�7�z@����v4��a$�\��b�N���������.1�^k�׸N�9	l����ě�t��%��&3c?6��ܒ�w�|M>�
�wݑW� п�����t�
lq����l;+���IP��j"�� �6Hk��,Y�m�v��G��x���*�V�c��z-_3B
I��ykY����U��d*�R�.i�Ò�f#LXp����:?��e|9��|&p�(f:W)����P��m�A�ς�E��.i��	<dDB���V�z����f�V��v����'4I � �e�<�̰���.N��� g���P���|��6��<�m���&�{ c��B n*�����s�~U�}�7f�86��e!�m�ٯ6�1��9y�Ǡ�l��EQ�\��ZOL(7�d.��P�l]f����In'�Vj�RsTO[��p�&�������FG�'�N֦�<Oi�g����H��d�tW�?M�`z�%�9!����V���D����4���䟐�
;��
���}����X�� �~n�Ϻ�;�r�}J����=��ٞ�>y�4J=�{~甭5k���`�:A�dt�:3=��qM�y2����,Y{���8ۢ�+��3aoU+� u��{��!<��C(ټO1N�(V��aF����c�P*X������GkQ�!�L�����I������
V��8�����Ġ��m�9n�~1k{"�!l��>���(�?-C�����~�^�8�0e�xR����������V7��!�xlP`�c��ήz�T����;��{N&�_;�E�j�#�+��w���@m@@Þ�=߽�b�._Va�qv�8:����*�u�bK ��C��z$���E�3ar�C�8��V������e�*�K	�Z�8�[�A��
����?&�z�ġ>z�'�1�*�SbI��>6n���)^�|#g�i�o� ���U��ai�;��U����(�]�]5�Q�!e�j�N��E_�q�g���w�K��Q�6�{����[�v-�0�Ϛ@@D*�!\�C�c ��I�=o�X���'�o��>�_�PJ��'�dh�?/\T�f�Ѡ�ϕ�T$�ݽç��	2�`��b"I��dnʻ�U̤�U�ZTpeo���"3�D�����슾�~��}���2� 23���v��-�^X�+\z/?���FNfq36?�+Y������"U1=hSr��i�|�l�G��@�>�˰/�/F��%�҉?yJx���Vʿ~�˨P�J�_s�7�Q�GGE�s�7 M��C�,�A��6т������xg�/E�h%��I"�N��g���oȵ/�'*g�#�|�l��&�;~��3�LaL�g��B,~�5=GG\fpn&;ߣ|6z��2Ѷ���5ݏ,X��˯c�ˮ�AO�H��� �/���0 6P��.����J%�?���2����_w�`�9Ω��e�\�.ؖЄ�2��S����0��I��u�QԲ����m���"�I�SRK �>(/���f�b�
ǩc����rCG�)G�A� {ȭ}#k�4^~����D:�J>�Nl/�N�G�D!����@�+��7%lwW��Z��4�	O0�/F����l�yE"�
'�{�f�D��������h�¤�����O�O$�G!=:`�4���nZ�ÀG��	��'L1�����`ؘ�G�KA��(�+�u6�i	P���o��qo��b^A[ �y �����cy���ܛX�Ve)+I�K�/�	��o��c��U������u�}K4X��?:����P �[~c;a�7�?HF������4�P�gAY���.�"���1�j.����n�'��;:���[�*Yܖ���Ԧ��R�83�6�}��-�:_�͒��	�m���7&p��;�D�����6��~���R_p*�U�\�_B���!�CLU�����ɡ�jL�oW�`F���;s��52d�$K �p�}e��0��U�B�[V�3��ɬ������Ś(R��H�LA��Y�#2Y����V����� o��ҺE/�S5,׷ hqyt���T2K_;d�>�K��z�3T_�3�Fj�IV�-�2�|!Y�"��ޙ��V9�B����͞_�@������m�.X�S,(Fj�'�j?vL�)Sm|�&�m�7�7��v>!�P�Z� �W��:�"T֗M6�	�B���,�5<Pȏ��#U� �[i��y�T~��xM��F�t>b� ��R4��o/Ї0^��=�"qEC�����S����u�QF��_��7]��Z�H���4i:I�iH�at�� �L��e��x�s,�D������#v6�p�.�t�P���~�<t�Y��L2e�-�Zg����y�#�|��-��lW+X1�M�8�P�OZG���Q��L F�T�T8��>��+��Y���I��u!�|�F�J{�����z�?>C�x�I1�a��68�>6�f���Y-�B�-�`�g�	�i���T�Sȝ7��sW���Ř��R���T��H�k7#��ŘA|f���"���J]���V?@��>H-���y�&�D(l�O���oaR�%�a"V����W���ӭ��
~��� ��,�ʕӼj{�J�Sޥ���QxpH)�Gh�M�n2���%g�hS����3a��������Q�z!��{!�-IĪ7L ����$/�4�zF��b�sa&�l��2���b����l��C�p�Z���k�/^��J~cg씯x�8".U�#Mi����<;�db��%}]���[Z�[K���ǰ�f,�쳽ףQVRj��?�};�3�ً�[:�@�&��c���������$"�fUn#�z4K"���z��\,�a�}j�=����.)mx��������O�1��6j%��G`*`e=6�V�����l�%��%4q�&V};�5I��e\gό���.ۈ��8�,��à�w�V�"��J�.���u6�n��c����{YAb�2I��%�w36/hp\�P{(�T���O��V�~}$�^K�zT���å��	�U����n�����d�n�������7�%n�19�"��4x��ûY/��]S��G�Py��Vp��[�ڶz«�*8%�p�eg��K�3�6Q�_��is�\�1vsF��#�\(��	�|�j��,�h`�����a1eh�M4%o�c.��R�x>��䵦��K�I�Ϭ���f�.�d���[%>��<e�,T#:�QV�OX�F_��v��(�/S��%�o��!�H@Vbd�0^��P��Ŷ�����w"AH�{��S�k�jC����u���e��}����NHy��c�&���G���N';'U[v�#u,���˪�Pd]�>��h���.
1�oNeI����yI���d��E�qv��������y�K����o��w��brt����8�]#y�9���M�l!�:�ͤ��a�5c��.Z�T��H�[x��$;|��vx��%*e������̕10��f���S��_��DLd�tx�,�B�\x��ez=�
}�hND&�TO�w1�3�c��J�m��DNs;�G6�=���v�������97��*7������u��7F�R.����?@w�rV���ǎ3�*@e�V���J�1��>���R�9��'KI�(5� ����0$�80�Q��G��b�z>�`q��Z�M���K��Ӫ�,�
%���(Wvw��h��A И)�����;�PZ�2��w
�!_㑺�V=�bM>���ԃ>T]��\r:�������p�Ac+D����b ����`�ߌ��GNҖ���Q���̒�r�H�pt���w'&�9wD�5T�{j�����H�#�b�K�o��(����G���y�{�[�7�4qBˍ�������b������k~��<��X�
e{8&+���@�#��@u��qd�+k�p�q�T$�������ھ�6�sa����+~��T6�'����h��irz��a�������"5[�`-ѷC��������������y���У�&Xϓ�`����g�X�t�;�,�- P�*L��QL����4��}i���"�ֵ�K���A����m����`�nT��	�a�>-EO0�z�	B��8�y0"���5+��*���
#����.�~��U�,tm�M�:��$K�@�.DcY������j[r�N)�Gg�Z�핝Zmh�����"e�x�T��0�~�P�R�O}�&o�I�gz�p�n��Ը#��r#i�lT+�"N�{�VG��d�N%M��8*����Ƣ5	h��\9�JG\��W�g	�"w�we������_	�uK��!d{�D�7��zwt�&��ߒy��Q�-��0e����w[�?1��y����?лm�R���P�g<�P����L�9���!(cӷ@�h�LU�69=zG���,��o}3N}Upy�P����ᔮ��J�"3�H뚷1>��C^|`�A���T+�vu�0ѹX�tع�m<���O1��s�p��� ���п)Whr����S:P̈́�g-�/�kÇ�ҫ:��x��+
S�p-��k|�C�R�%#��a˻��1�>t6�X�.�U�6Ž��w��G���4���Z��b��U��ޑ;�j�G#n��EY��W�Հ}-�='�����ګ/�2���,{ð��Pb�QԺI ���7l�[�z�1O��#A��/��I��`����|j�1s���5%@�vba������y%@��i�4��p4�v�j��<s���Dj��~���L� ��v�g��|����%�0��*^�WWn����4D����O&2�@�����r!]�]eD�
c
W3�E�p�g.@���d*��]s�R� ��	�=>�%��6�x� {�|�r�7l����"���G��:��^�=�
(����8���eq���^�NGDQe	8�c�'�eB(QS!��k$���zcEl�* 8�­L��/L4k�~��Ы2��E)�Nܰ�A���ѐ��\��ǡ�k�7gG5�σ��ţ]����ò��orɧ�`��O�T�{&�~�u˨a�X�g��{^NGL1�"3{W'V�ё�Qs���jx�Jfr<�ol�n|�,T�P�a4��(ƚTx�&�'����@ܡK`6dE��	8ʽ�;R����M�pə����P	CE�<�q�a�
�n���E�_�8PLg�� ���WF�Ѣ,�p����ߥ��M��P.���Q.�F�����߹��HLJ
�E��4n����i���з��_�^�5ȳ�~F���~z� u&:�iKӴf�)���k��f���3�~k�FKF����y2�G?�7�N�fߚ�*@߅�����܌��`8P�d=���G#1�pOp��"/^p�ƙ����^nv���̨o�f� ��NX�G�+Ym��pJ�P�:q�B#�!��s�Qi�"�s�cY�S���{�>������٥0�#Ɔ�l�mꌤQ��sQ�^RnQHE4�p�/�l��v�$gV��3�M�B�J��AJ���l��d���!�t�(�-����3���?�WT��~�^k?�&��уq'9W@]!��Q�;g�ylU:4�5�W2&r�&�Y%��̜Vi�j>W����8��سІ�h���Ig��Me�?�P�t�	��̐ݭs�!�A���*�l�b�RH��G�̼�<nǌ����?�n2-�l�A�g�G�Oh0�$�4�@l��|S�?��&���
;{�2^���y��^{):�`/�v����`&�׵�О[��t����� ~��w�v!͍v��YT�Fs�Xr0��w\V?� :�o\�=5�B�;e9l�=u��Co�Gk�"y/�n�T�Qte�\Sy�O^����8��{x��%�����]y��0�Bo����Rhs��8C�s�BРC��?��I¡$��D�B�ȍf�)iH'r�ꕾ4w=Gt�W�8���p��2�q0S�w����J1���Nz�>q�cˍ�����-^}bI�+���;�>���Ǔ�$R�\h1b��`�Gy5Y�k����ݶ�y��u�kkx�DA�����xb�
Atn������#̍;a?�a"�uꌙĉ 0�����I����Z��?���#LB~�x��sM|Y�0/�tO�7�qc����F(#v�'�wLo2�U��%�	�s�
G{�=��_Փ�W.����C���|�8:��E��|u�y��B��
�¼dI�g�Ui�/�/a�J0���x�S����Vp�[���~�4���A6�j^Z+��83�#H)1g��"���qt2�y�-�t#�؊�ͦ<c+�2�}�i��փ����^&a2��i�h�s�M�
�)��:#��W�����.�����;*����;�	�����Փ� *��^���=���L���ųGQL�cp�	&9��#7����,vۼ' 2��ؤ�H=К�v*��4��B��|�2�������0�9����ӗ�M���r����vo����A��8p�&�Z9h����~�����/$���C3�������23�/ "���C�j7����Ux�)���>rH��冹!�eL����Z5PC���S�(ig�26�.&�S e&��hB��/�6*uK��*�QG���5^�@��`�;�e�ر6T�[�P9�<�rM�Q�S�6���Tf��vK	@(z�?�V���"F1���F��(���p�L Lp�ń�u�е�:�Y�߅�x]i[�I���Y^i�|l@({��tx���Дf�3smPK��S�M�YV�+\]�����x�~γ	Zc1d�n
f�gmH>؞�Q->�RB���t���5:͙�Y��ݨ�饙�6d|Д��v{	�s�+�L��d=��NjH�XףѱS���3����rOm՘�&"𧅵O� �4ˑ��c��`�Yr��@e"��ʦx����؈\o��}��u�mPg�D�s�"T\h+�F!�,���}Z�B��J�����z|��[�⥙{x�D_H�=�c��x=��<\ؔ `�	X]�&�p鲙T-p-�<��3������_�|����E����^c��F�֤��Qi�����T�w���V��wb���ğ.cX;H��:��\���;��,��:��s���qYj�ų�\�0��1�֯����t�����!@[i��b��X9X�V�&5mԪ�s�^��[�P�X"R��N���I,�NnA�#�pL��;���ļCze,�CI�	I}�����s�]f�^f~89��}��q��{:9<��	9镡m��*_����TNDe�_H>B"