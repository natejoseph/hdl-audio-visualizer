��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���֒��&�ۥ:��Z�E���fF,;�s�dK�����p�����X����iN��+��/��D�i|��K� � #3*�[��T�����v�`>�h���c�d��pho���/Jz�׍�P�)JB��OY��vwd�=*S�,�>\�:��<�r 08��y�ݼO��V�C������5bG��.��iG�|
�(_q�"�o�֖�3�Mb#�ð[)�����}^I4+��:w9��\7v�(ސi0U��W�@A!��4�ʵ�o.����v4]�&q�:��Z���$��N¨γ� ����Mqm
��"��q�V0Q�H�_AG�L�b�>�;�."&��A�-O?~�����i���ϧ_�7�r���5Nx��n��Q^Kkj�"�&�ňh�^6Eǅv+�b���{/��y�+٩�4\f�k8�Q�n�o��&�C��5���D�h-�8���2$@(`�ZR:�#�SYuF��K�>�H==X��'I��J��B�Y�xK�u>ۋ��X����+:ƍ��x4�qhs��+JZ���}��L o�ܣ��zy?|M�}_�)���á7��V1ԇ� /�׀5���:י�I�T�:Tt9��)X翩�zx0H=����Ͽ|���AZ�e5�A�}�ZO�?���p8KCli�uX�y������6m��/ԩ���㫅"�2��	\��QL/�l���~D��k�!�@v�",=��D"kmh�����%i'	��@�T�^�^谮���2H`W�\��b� w�
Rnxl�ݤ�_�1�Ҭش(M
 퓢�-�>Y�k ʚ�7z/zZ��	��i.�����S�Z>ܓ�G��KctHn��*���!GJ�i��o�`O�0��W�M�����6˚���fS�; X��@+d���Ⱦq��#��~������F͕Ա�φ�_�ۅ����*c��K�L�;YVg��'0��Hz3�1��Fn���ي�=�iE��l�C�[��j`ו'��[�(k�����r3�L`��7	"_BC�oί�U�7}�˹����b��E3��ļ��h?�T�i�}��޵�̼���l[����~p�[zB�����+$w�G67m�I x� �6&t��f�DN� �T������J^r�8,�/���dm��b3�߹�&�� �x��W�g k�H�Q|������Fݲ�3����f�O���{�"��??�8n��}k�&z��Lz;vDf�$zLЗ���Z���X���kV�y:Q��7.�2�M�
��yz����;총�"Z�$�>.��F�Aq�]ǡ鳶\�)Z���ˡ�!Jy*
h���S*��kxOos:e��NZZM�)Ѧ��w�n5Ӭ�Z!�F!oV��@+�̚�)j1i�H&%�U�M�\����M�.^��mZv��G�� ����@����3���P�4�9I�R=	ZV�Y���C5Q�n{�"��>�� �U_�yѬ��[4�2b5���ʾIt�o���s��t4?��p���+12��V�r���A���v
!z��#.,1éYE|�P��n]��/�?�9�k1�&��1e����w�/,Ȣ�ر�������pr�����?ſ�} �ьOwC�Y��e��g������=��� Y{��9��(}�8iL�>�M��V�(���^�@����3�K9< ���\����k��8�p� bn��>�;�T���������2Y������*�	p�d�;�r��wIb�u��2��ό+,ڞp�{tV!�#�e�|���&�'�B?[IRT]�s�$;=y�	��E�#&	�x)^?����Rx���HX����W6z�9k����8�p���^��B[�����}E��ϟ>܀ϗ�Zb�z�}0y(�+�ti�[�M�:w�>:[�Kr��A=I9�g���yA�?}R�)Ɣ�0����X���U�#�!�S��y�P��4sݗ=�Ȯ_����5���1�ͼ9]�����ZK�mj�������<�ImÚ��լ��!��6�P����Cԃ<�$�D�1%Ԑ���
-f��Y����!����'�8������6�>}�<|RF|w�1�v��E�0L^3�+������ ���s=�Ә�;��l��������{�$�`�|MwB^	E�7�g�Φ��^>%k�Z7u�{&��q�	�М?�˿k]^�٬(��f�3�0Q7��<��x���;~��N
Ԅ�$N��G��C������D�_��G�`�`
��\=�`������"�_�88�d�S�T �b|�d
��$����������~���������=��^t���/���+�~	p&����oo���i�e���;`|����˜�@k��Ux������?F�����S��دD��~}W{ˋ��Yv�O�ae@5o�d���Eۑ
�|=��v���`	a��H{67��J4A�X��騯�Ns��q��B��U|�㯣��(�܁��Z4<^�`�e&�j%LX��e��=MC���XZ�����*c���E7�ww�%b��:� mz���b�)�t�YM4@Y�t�Fݧ���P�v�����@��G��w���п	���b�2k�ʘ���R�!F՗����Y�����>�T�Q⋅q.���HJ�R�Jc�|WY |G�n��|kS� 9�}|�j�5�j(R��M�X�&m0-3���)��i�t:��X0�ajea�g�e�+)�c������B#��2����沄<xJ�����Z7���TE���������X�Q�����i��~�	�lAa<R�'(�q��o�{�"7E��ŵFФ���� %jw�)Т���oڞ���N��+�� J��k}��'F;;j\[����-�PU�ȳ�\�#��PA,��=��zT�I~{\��WF���Fd��XELgiaH0?�C���z)��(��/]dHz{a��i�KY����X��zUK�fU3�%�L`����
�ύ��U��%�b�e'Q%��������2)B�T�N1̏*������0�f�&7��|&��0<�֣u��J��$g�ʇ�ğ����: ^b*&ώ�QQ�"�y�o8�2((���Ͱ]�x�++�V�	��$1$8��	����g%3�B��K�b�	����ML���^�|��b�n>�/�I<��m���Mմ���%�2�C������b�,eeP_dv4��M��I���O��d��կAP�VTG�\,��ے���ʩ�j�J�JB_Z��Vx�_��ȥI�]T��7�����и���^���b*�u#��x��3�w�jG;�2OJ6��y��ˈ
�7~�:�BL�����U��6�-��>��I'��K%���sq�~�ɇ�n���0W�iW�EӢJݏ��r�4L����
ؿ����u@�R9�A���w*�}5E#L�vr�[���{l�O%c�>Ȯ� �i��;�����|�eJ����<k��eQW��mG���}]�����Ok2�|``�0��7e��.���񋩐zm�zdme���y�Lܺ͘2��3P���߳�[$>�s��N����<kC ��p T�a���H��!!��s�0	�^:i
p���ڏ�@�F��V��:��JE,A�V���U�m��xm!uy�1�	C�(�Kn>Q{���;��
���l��ӱ���yAy�|�*!"p&��1xΆ�,{�r��[�S͒=̙ZN5�GF��y�m�N�Y~g�"�N�5c��b�$=��Y�S�l�^+ŃW���y#U(N/�!M�4=v��o]��}�d���
F��lY�}�!��h��vyA��}'�HY؝X��=<�X�?�b���G��0�������.U�Ӓ�GP�A��	Ced�Qe����$�{ȯ�>X�o&�Ž��f���0@܇R�Ռd��'U4�@���Ș���_=:���85�ۈ��'o,�pSI���ǰ}� w�w�_pZv�?Xv��]��.��Q��C�3!#��$o�>>�03�s	sw+~-��n�Y?��ȣ�Q��q[̦�i��V.+y��q	��ܨՐ}H pq��~:��z�Ô����\����p�N�mUCO��u�>�ʢӚ �=�h(�q�ZrN���pS��\@�tX��X�ކ;Q}h�� X��E�kWL8&�T}M\�����`69��o���;C�kQ>���O�w;}3�8"/���^�k)H�D�v%�ޱҙ1�l#@aj��I���^}$̎Q��"�X7n	���щg?&��kP��%`�y06���$?V������ց#c3t���@
�LG�J��1-�b�J�Ŏ&l�݂o��SS.�d�~��pHEC:RS��씫{��$i�Ko���I��5X!Sy��.$����o+��	�<����`2��@a�?�x4&�(DŔ�K�տ�����R�p�-#���
�1l8��u��!x�����lY/����xp��أ�H��`��6����]�7dpL�
Ufܕt��Q�����{=�׬�"m��U8�X��`��9m���)��~Dvc�?�E"��7�(����`ˑE�h�x�}���� ��*7'��9b���s,)� �Nʢi����&AQ���N�I�ՃT���B������|����,vҷ��o�{8��9�����ӎ���=u�	���j�-����<E�n��9a����&��I�T��<�K��vSLKW*,�In��RC�x�;nvz��Є�妷D I��T�ALK�?:Q���k ��zڻ���J��li�skk��.��V�+EʇT�.I%]��Wh�f��.ό��Rp��WE]�ja�q���6zKz��Su2E���i���B�E	L���N��-��oP�,�b��6G�d����d�e[7���������o^�؄,��٪�;#��)�w��~�
J�A�E+� �Db5�Λ3Va��Ǆ(�=��T���KGD��#���܁�c���p8���B��=׵�LWT�����Y)�'�뭵`�+>�`��K#d�F�!�8I��k"�tv)#'��XzY�=���`9��w���iK[��q��0��ڹ�M�����:��v~-�B�~�EV��d/~��5���� DS����������ɺ��<!S���(H.�A��uͬG����6��4'���N�*� 4��tuܫ�����.ܫn��6�Va�d�G1�coS}��������$���g���)bp��N.�~2�xpFxfbt�(�j��^�sO��T��ZvG�Dɮ�<t��֖D�����.���xmc&���caywGL���YܻX._�{ϯ������&?��a�!X�0&��ϟ�Z3���J�H�5�?���w�	eJ�����OND�$0��.�R<�h���nX�m_�s>��B4���}�Ƅ/�Y�x�q�Vb2�,b�W���� u�6ֲ�a���PǛ��:�u����q=�z-Z��%��1�=񴜐"�^��{�+e�_q�H
E�Ԋ�
8�rt���d�ǄE=�_ʤ���z��ѵ�>.aN�A��5�#��K���|.��h����7�уD-jj�8��I}1dF��B����Pr�3k�� zhw�:?��9J��b���K������eE����f���`O&WϜ�Ag��*���'����<Қ_Z�����J"��y�����03�5�$��}h���2����=D����Ǩ��*o��1�c�v�w ܦ���r0����a,+z�ʶCܤ5�Y>��֐Q_��1j��h�xQ�@:V��Լ��Ȣ�r8ɴ2�h�0/y)�o��J��F,6�$@����JWr��O�I :!��P
ԩcf����D��H���JW����Z�,��� rA<���G��6�c=BW�j�����ګf��I���cXR�=\H���!|bф�2�	�r��6ЇbW���q%�©�X.�6�"I�Ek�c%�i A�ĺI��G����LT�qDN�(�8��W��$1�6������j_zV��1��bn�L-��2���y��=��D;��4{&��+�,���p��\,d��6�SG���Ć�+