��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�p`e{�z&�JX����{������ǄTfX��Իz��O� �FG~-��H���������#��M�7-m�
"��xx�.]�Y�{â�� ���/�߇�����Z��0�Q�"j�a=e_gZvV�F$R�6e��>��)��!}M�*����.�k%��W�}��pe�V+<գ�W�G��T��*V�)��\�������V� i�+�@��+o�(�ɭLP��?������H^�V5�bG;Y�1��hZ�lٲ�Љ#�䱚���z�;��kD@	����|vEYn��-��n"��9�/��Zf�HQ7{~`�V�9��Kqf�x��)O4��n?6��T�m��ʊƆ�\��=��G�^��9�9@P#[�<��l���@?�0`��?71=��ؿIY���g��X��v�x��TmŦOG(=sj�J4�o�v�KO��6�� @'�G]��[ �C{OF4���1V�.ش�p�n��#A�&y�׫JNW�b��[�r���������͂J�_� H8����m7�j~i�H���9PA��Yx��4��<MV<�7\����^j�5��52�V(�mI�V`�w���Ú �9��+mF?�=������vOD�MVN�@?$Ѹ^2�l��>�����m�n�)WF��d�8YpTQNzJ�)�B2�4���O�&��ސ��4Ʃ�M\�c���Mѻ�������|�n�/�6�|��K�4Q^�Ǝf�m�������B"�[`��H�Vǣ4tZ�/&4&���]���Q2� �VCI��ݽ�������o�Y"����	���`kV�)U��l�Þ�Ƞ�M�Ǆ/�S�"}\�n ��x���\Ț+.��V�ࣶ���C�Z�������/�wv�"M���0{��kv���Y���a	i�=�#+�D ��-7V��@�5̠�^-*:�r��v�0����D)W.B&檟sӏX<���[Xn\H��_3s����F�� �������Q,�ؔk?U�Ge����W�E���u�i���:v�'���j�M�y���ώ����8�ww����gt��8������!X;�[A���D���g=4�Dn�*Z�=Rq���WN�Ɲ=�ώ�\i�fhi=�f��\����\0��vnY����E�U��(.u�-��򄭿VMR�p�y+Z���p\������k�paZ���7���^��vm���d����C�CZ����[��JD��Y�T���tN�P��5���	��34�K:�9�9�Um`,���ؒ>�t�A������Pf��`��$}����e-��ñ��|;ft�Y@�c �����^[]�@�@�����*���S�V̩�U�%�m��{���o�isn`�PlP�Z�@��h!3��)�7�ifo�b4�૸pW_�jΏ���GA;�Dj�gdT��G�o��TӮ�?b�&2��M�kt���Z�_!F�XwEMF	��M���[Y�Ҵ��	�@`H���X�����2�e���ɪ�>u���j����T��yM����ׄ ���r����	�C)f*��v�*���.��qp����T�hB����}��*��8�>��O4�|��U@�=B�q<]p����F�6��V���T�R2���ȕ���fd��!�����f�l,l�z�$�	�h�7���Զ%�,��TO� ?FzQ=��?k��4:��ˀ�6��5OA��g�]��",���CI�9{��mf�ݙ��׶���O8��d���txޕnFby�y�Ni<��:���O�1G��d[#�u�tKE%��}f�+=i��4z.ͺ
)��>�@ڳ7��*��t�7��V>�M{h�FNe����c.HD`ћMv�d�vQ|����ki��w.~�b��4E�'%��7#�������N*O'o5�I ��6)j&��MϘ���/NO�'�~�ceV�Й���V.3춝�弑�x��'�\WR(�����M�}K���*��>�Z���O��UP\�rZ��K���H�h��OOȣ�?�4٢�_���c��
�ڇ�eݘ�F�&��������3��zY���Ͼ�.�KCm�c9$�'�����I�W2�h	ej��*4�./� ��W���t��U���)�A+M�����i	2�(Jw��_!4C���|�Ë�lC���pF`8������j��p�q�e4��&��?]�z�����ʗ�3o�sS�dsB���F��R�:���>ű�塼��&LV�xj��<חF��eǑ.�:2G�����x��?�*A�ɘp=�AAz�U%�l��y�՘>�7�_��!�[�?�Z�\B.0z��"����~��c��,A�M�2������施����iqǗ�A0��y_`�e���Y��3�eF�^a�����5zr�uC�3��> 3)Ȓ�7�Qn:���l�_J��B���@~�U���qbi�:��{�Dh�-�~������"�p���<�������!U���QH���WD	9��ĎC��()�|�O:f��l�91c���;�����z`�Gʍ�m��O�O�/ �qf�ݩY�'#<����k{NXϐuLw�6B�l[{:�}��ʌlƜ:8����/�fjd��wr�f����g�o���� G��-��{�ui��>�k�)�d
�1�����By�
������>Û��a� !�0��8_����
�_-���,8Ե�T�	z�@����Løgڐ���e7�����9�\�T,�]8�n3@3��H}�x	��2��f�N�=���K�G����,���m�o�hW&�����L8R�:��!��
q7�e����n���E�1��Q�|2�c�:O4|̊jȀ��t���,�-kDc���s�@����l�>���\�QJܪj�s3��%�=r(�4�`=+�0EX�ZpQ�a�31
�V�G3��>oP~�~�9O���/��	�"G�N�??9��������;�70n�i�Ȯ�W��I��O��3n��&��.�,���:���f}��4��oXI`����� iǭ���a�9c��5��x>x��&/��/�e���c�	��34��