��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C��Oҷ�$�S�u��B=R0R�E����X{W�yh�)Y���ȷ[��Y94Z�|�cLP��!��U��se��\���?��C���k �:5\�,��I��l��:H���C����#RH�t"�qͿ�ǆJ���F�J��↫���������_��g0��?�/w��Y�?'�R���ئ�m�T��jmdK7O�0���\?�m5&ě�	��];��v*m_�#Z�M�{��f��ٜ��ʬ �&�5(�^=�V����kf�|Y��H��Lz�w��kD�4����4P_����ΐ�l�cS���x�W�pl���[��n9�{�dUp�2�߭b���G�~���A��?c�i!T�4Zd�$��'���.�v��g�y��;�g�r��cGb��_2�r�qP����t~�4 "��[��[!�<%9�/�GL�)mB���CF��B����5q�^YW��a�c��GB��I�5]0K��R�.se�+##s��W��9��'�o�c���I���<�Z^ŭW�Iſ�WꙎ��-y�"�:}�R��t�މ�C[�����3^��@��+ߏ��þr��5H=��i���� � j��2U�a`��T�m}��&'�׆��Wp�녷��®��X���p�H/gJ,�ۆ�ŋ^���چ#�3~Qn\��Gs�k���
�[�E����B:�E��p'���i6ד��z�(�z��^�/�R@]}��q�����/f�XC�Z[I�ڧ��6��w���7H �K��$^E���&6�F���r�g=��s��"25�u-��\X,D�ư��Aԝ�#�]H���n�
�+Fx)ϊ�m�"l����L_]�g�'\0Jz��J�ώB���QM�`�3/Y��=�Ws��ǰBp�g��sd�K��Ԩ')�^7vf��i��5�C�O�;Wnk�>�b��� ����"iP�c檠��e)*�(eн�`�-��D��"�.�.e%:"��}t���5Ka>Z��LG�s�xw���dmm�[�i�+R�W���a?�浳
>���G>X{9������Y�_m,Ӫ��m��"E:b�X���Q��ᨼ%P��h����J:���o?jCAG����R#o���.5Md�U�6Y���W��=O�@�Km},�,���6�4���PGzlNޛŲ7:�h�wF1e�s�H� +����{ᔻ���Lb��#����p'��^�_h7����D��O&��Ÿ��P	�{���]�ysǆ�(����l��kn����7��1���f|x*bt�֐pZ|.L���>���#��2�鯾��{L{7~s�A�"�xgPǔ>C$fP	j?�	�9�\Ew�㏑��U�Ĕ�Zl7}�P���V{R�ż	C��P� ���k��J/���Uݵ�5'��H��*�Ȳ�M1�3��א�y9�2���ov?v��'�����n�V�"�1���������/���t{��[��F�ak�	�k&���U�7F�/c�*�x�a�{�������M:���E���x�ͤ+o:LpN}���>Ƭr��Kz"C���O�._��iVN`	Q�"��?���Ӷ�3i-��Qړ�|QJ��[�|�o�u0�5�8^緩��I��A��~	(�����^�P��y��]�9�T*;��0D��MW�v��b�����鲟����\m���f��W���^>�(�*BD#�72`�m�!ۑcVG��(�����ϖ�`�L������[�"��s��>/I�{�Sh�U�M[��~�u+^1?eC��//1�H���]"P�쏦��]�ȑI�����^����K"dI"�m�������7Ѷw�J�*�	�$�uu�~*��٤Ec7��Ȭ�&7�H�����DN�4�'/G�wٶ]�jZ9���&vG���-���OO�D�#���1%ir��p���F-�U���3x�_��>����C���Z�W���v�<�0:�4��yA4�N�.��^��ic'&��鐳Q�oz=�����D�hG�6�I��!�.������Y��o��J����-2���~fԡ��#�pJ�E���9�ɧ)�����z�o#~�0�h��� t=R撢U'7���UP-��a�D��T`k#��B���Ұ�巵LI�y��p'�T�Y��r�b����Wh:V��u�}�e{����/�w�ޣ�m�~���fј�#O�?uO���O�X�c;c�(�-��fX�;ʗ[.���D�.������ۥl����ݩu��/�<ҵ��r�|�c�R����ǁ9�{��q�A�=�ƥoݬ�5=�f�L�eT.ker��-<"���ύ[���iڱ�a�9�VL3�y6�}��t;3k�R!����}s�p@;I+��\��<~~K�_�;Z��B�$�ݔ���"�S`�N��Ҡ@�$&��Z��#i���UI����_"�$R}#��Gݚ��ԓ��=����T�?U�����R��b����e�2��1��e }7�5������/s&�w.`Q�ޜ�:I�n�oϛj� ��{����u�������%���Y#�v���7�J��w�%>���Yw�OI&T(�A^�ήC$h^c��K������&���1�C\W�w��f]��6������;�T��6&�mi^�s�n�ڂB͒j�BT�]gO��!��#K9��������/a����`��*��<��ݩ�4�&3�W���:[6�&������;�H��nZ��I1{�҄�>(~ø�F�S�I�3�P�v��sq	���iA���m����?�W�Z0L�ѧnN�!{{�R��:��Y�2-k�u�ո���|���Li>�*6����sm��o*��y�埃" ��w �:�ך����0R��X��ŎVk=��*�j2�Q�c��>��Hﱓ �DXc�I<����JY��WAX��s����Mk���z��;b"� �]�Dj��&�`�ǵ��DI�]���i#Ǘ���N�VF���EO��+���U����hb��Zx.���D� ������l˽ݚ�@���*t��0?�1A~��z.����#G�c�?�Cz��
:�ŋ+��fj�$L�)Q�UZwjP%D�^:s7)���h��%���b��`��WlO��g߫I�4���C�U����7�3|�ȿϸ
�!Q�F!�D�~FƤ?E�9�[�RGт.�R�{i]��v��"w��`��,���6�/�����Q�i���<�6Gx��M>�'x�Y��8ʏ  ��Tk��%G� 5��uМ&���)�ي/p����y	`�"���5��T���vɹ��ၹ4IpN�-'ZE94}��G,�t�A�O#t8e%���̃g�#ڪ8��m�&�z�#�T}��e.*2�吿i�W��[nr���� �LG5NS��̀G˓!U�"N�*A�{�P��ћ�� V�]6��HZ,����c��s,'��a<�y�}��Ihb�m[�@�F4X��J�x���!���N5�WX՚��%'<��������W߈ώќ����Q��N��Q�|�_c\����ӧY��c�9x��"OT#��O�M�1��\\N~�&i3��ДcEoO,(ǚuUXC�6.�.�;w�O�P��,욵�
ܶo��W��Op��Tn�����l�
r�t���$�����ԥTqj(��U�xm	��W���5�62_3�^j�ѡ�*�Z	*�6��6�{��&t��l�}�����	�?&��n���&N�U(?�D����lVE+;,�q�̕W��<	�����Y�pzu��s��ßN��R��ʒ�q��T�g2��Rf��Q���Q�Z���^�l[zL���X&4�͸J��R_�"{R�j�h��DPk�|o�m�9ARz�����Q-�BV\�������'���V�>��N(j�gGQ�-�`�AH+x�gJN^k�G1���2Y>��+g�,G"�q�?a͠>����8��5h&����+_�[ʅjf%g�S��Z��s���L�|����۠�E�-�k���Td� ������z�
�\&��� ���t�����;�t�ڙP=��
�r�-��|�0A*�pK��@�S�D�f�&�T&T55h�뗋n'TW@dVe�����*��EM�x_w�2��#`�gR�#��������7����~S$�GnP��V���<3�s�ĆV �Һg*��֚���k�N�ގy��ǁP��P&����w����W�mp_"k_h~Y/�������]�,�Z��}�U���:�HU}՚��b�d�K��ܪ��9��s�H[��gj���P�>��.��q�TK`��7�Yt��ƃ�Ovo��D�j@�!��Ϧ����O+ ���y$!{RDbBn�K�K����W4N�`�"�y߰TH�:s��G��$@Fp�)��=��.G[R'`*��Ǣ��.�I�/���ځk�.����w9b��ω���`����F�y�����+Dj�(3�g��6y�I��B�LpA��@_ґ MuJu� 6��"��,�m^�0�1�$����c'�.T���n.�2c�z����L
���@s��b�E�������Rj����������)���j�J��y�&O��]��.u�����3p ��>���%�M*)�;�Ջ����ZcIo3�mƤ[�wE�����P{���e��XI�޷!;M�T�v�4�b�_l�_~�}�U��$�>� �/���0�]�����.�9㒾4 8��W��y���qa(g3j���3&����TD5���I<��g��M^&��	���9iOa�������x��i����:t���~"�αn�#�yr�/8�hM|�� p����Ck�[`<���,5S�L�:m� Im�̔���ܯ!�j����q,� �OC�o{!�x�]� ��G���t� ��(�F�A�mV`Riv݉'���B�E6 �9�O�[iw�x�L��C�EdoVO�rdi���-g#�S��gS��e����t���>�1"�h�>U�����i�I�H݅HV��p��iۭ����W����,����iz�~�a4!�M��nB�;̹:��Ц��Ԭn����(ˠ��������R��D�����Q×���1��u<M:"'z:+Dʻ��V0��ҹC3gd�5�ħe˓�'��T�ʮ2����'m��޾���3�z���s��O��	*��s+	�wىlP����vz�5ӞP��S�N/' 8��A�.�R1���j�=�HC�|����aa��" ��d���#�6����*s���"u2�Go���y0�`�P��e���`��Vu�8?D8#��X�<T�&��yOq��
y%�bߵ�Paz�A!��i ���2'�����p�U���cS?j�?O�v�fv�ॼ|�B炵��5Tl�����.���jXG�p��#�$sk�o�SO�S�}�}�C��t@$���.��2�c5�k�wp�R���dT���$�����-�G|��m�[�L��(:8��.*,��$؂����h�]H�:��m�x�������pa���3�*�%Q����'D��<�ź����X���v�Ѫ?�w���5]hQ���C��]�L�Ҵ�U�T���	�s��<g/90�.C�0�$I��5g(oWN^1�)ĳw�)"Fy�|a@��C��(�n��Ĝ�CG�=c505�̝����k�pgt�HdY�ղ�mn�NG"�3gv�>c��>����]F.Jox$m���&����E�O�A���/a7��9��k�\�E�b�	IJ�{�aZ\��$��-bEt%�:��Ju����s�m�ݐ9�a������Gs�F��0m��J��˪�d�Sŋ� 7`8�86t9duɥ�#��K�/1��RO��y+��i|�!��
+��<T@����d�L󭗅�I3�-�������ɛ4�n�g$�+�0�d*ob8��L�y��=;���~Ě��p ��K�ހX�[f���tٲO[҆hϒ�2��l��mr��]s���������@�>�(g9�\=��<!8� �������<�[� ���aY�88�b��pC��Vh
6�j�z7� �kj,�s���_i �~��2����[V��%��!<�����/�13ߤc�VodW�_���$V"m�Â�Z��].u�۠�VP�1��]
_z:��s¨���W�m�[U��!�m�G_�YJ������ͪl_��=2�e�W3���S!��[��%��䷌�8�I�#�uC$��L'm_�zy8
^i�E�d4��AĒ������f&�� ?y��da�{Ai�Ðت��o�%�s��%��dc^�֍4��V�[�U��	����9�p���ޕGM2�.�:���R�T`"7�֯������W�5� ���+��[����h��/:g�l	X���ʫh��9��-#O
X#��)y�8ƀ��>�{���YH
k�9vg%i�Hs��'R"W^:9���cxʥ
�	$�Ͼ(DP����M�{>�	X:,H���rx�M`\�z�9&b���+$��,E_m�?z��p�i�4�g�,s����ͼ3!�.����!�7)��P$8��Pv��J"�='L>�R�W�|M��:�B�񯜇�O�A��9����V�3���*���p�n�+P���4:~�̓\PcL���o�A����4������h"2x
�8[�K���Ϋ�TS�Zp�l�k5�S��=oNi3]=����)��d�؏gmμ��ȩ#���a�����Ӓ[�����d~��Lz���u{���<�7�C���ɨ!�jme�8�?�s0�1C���� �axm��wv�w�bc�q�p��3��#:ӿ�Gkqц�x����m���;eH��1�{�z���k�E��"�yw��6���?�r݉,�dd<�
��r�hԉ^����>H�q|����Ui�,w�������e��GM2O�ː�S��'<+E�x��`�W��~��z-�\�<=2�&BPV�aع��S
�15������w�����ש��c�����Q�7y���2�N�����Z�ٺ��$b���4��}*��;T��&���Cp	� YdӼ|�����~�7��n���RԹ!�	�T�|���)_�8`)���N؈C�j����T�Ԍn�8��r�^s��$��l��K��b=q�-��$�I�!#��0C�8l��#u���1�l��&`8��4�4��i�1����Ψ�\�3�?jr����� Ԁ�Y�}�m�g�5!J�'ԣ-9��"���\��v���}���6����pI�r�s�[�{(m슡CLy���\*ꂹdO���-����!��X���\��ۦ�]v�q;#� RX���?���)�q�L�ۧ\0g�����
p4XBD��-��8�������������o��X�^��AWq����4-��C�P����@�8�/8�Џ0GF%�`�	chI)4�0`�Aٹ��@��$~śƛ��,��9&��V.k}�Z��ĕM�jCBZ�@�����ZF|ƈ�� µV��y�L��
X)��-޿��G��J��XsFn4M��LH�A4M}���A �1d�a\�Bl
�_8EΟ���0ߨj���T��hKMQ3�}-�^��'T��T�֗�����
�N�e1�__�&�KX��ݲ���)!+Ϳ�e�D���0_�"#��8fr�C��:�����?x��oui#���ȧ���?�~���߻��Y�;ĸO?s��L#UY�V>;sl7��,{闑�+�����H�@e�)m�Wq�c�I�9��O��d�+a _����/ty�������zt�̟$�C����Z����	?n��R9���x���;��M���{�z@$�-EZ��M_���ެ4�
�£<���g|tkYC�/����̃��2�9�|��F�Ӝ�_rA�[*��㰪���U��f�!��f\�^�k4��u�T�%�Ilq�~9��n߰@�1�?O��m���IFƼq����i٢� ���?��q*Yސ0�}�j�MA�κן��U�����.���6PQ+�����lR5���6v6��(�/��=�$FWq]<ש�eT_�S1�
�F���08y��A�=������G��#+�R��A\�7rͷ�u\���v�"�2f"o)U�B½?aَ�M0�ʎ��!�;7��ۊ#ঢ\<�W�M��톨�r˗�զG��s��M� ���)B�[����o�*���MBK ���Q��������wꀇZF�ڃ���G'!j���d���iTXc��5�0��A�Ii�6�'m�Q�.�?��UfSY�ͼ�n�� s[\�.V�͚fJ�/���?�'ߢ�#g�?ǘ># ]�Wg�}�������s����8�&�S�jO-�|����*&�)SR"I�(���X�33��cܶ�Q����DyE�ΐu���!ň�l�BZ��������W>�������50���~ ���_�����޴u�����J���M������IǢ���7f(��ǰ�߆�e,?�;JR�H���}3��SmbĐO��TZ�TY^'IH<f��,WP�o(BE�-x��p=W�G\�> ZՄu
��C�)�
�HҸmg���0]�_u�I�
+�İ�|\�i���ۃ�ؒjz��_w��nG��F��˗*����X��?��#3���q}����r�Ь\E᥈/�U�g~w�9�LC�n�ܐg�(tQ 9���� �ċ4M�ŒfG�=��RuFZ���n�EC�>
�j���
2�kOoĠ܋
�]�,�S��'�N�$u;�'��Ik�Jl��yL�}~���4u7�4�v�}S~� �����#5	0ߝ�#'�p��sy��V凣��dpZH�z��IZ���`jw�gQD���MO�|�>��8?�&PrFe�غ�0_��"��N����q�=���^� ��� �f#R�t�����$N��O�fJ����YO}xg8t�v��ԵQ_�>j9zu�l��0�G�d� �IJeD��� �+��$�m�������=;w��~���(�}�$xu+��ap�1�d��%�͙��v�}�!����j�X\���W�a���E߲�Y묕%�k`A�����
�8���=oPO����r_���Y Yw�e��v��#]�~�1X YOJx��D7+����.�F�P�A�KR�8m5���V�e�_��Z��<��ڹHѬ0�X_Lk!�s5�y�$�x3�kG�Ǉ}DXG���4>����Fm_����\Ǜ'�܇2�Y�J���1]�NT����'E��l�.F����w�_ OJ�
w��*|f�E���p�&gw��
�y��p詟ߑ�) [�~'��A��@o� �<�Z��E���'8�;~~T��U���)8���ł�?��4�G�_�i^G��@=���Y֣��/>W2��oPAۙ|&�@��M	"�3��Za(ܢ�xĚ)I��:D&��u<��4�$ ��v�T���* f�%tW��P�s������� ,p@�L�i0\_Ą"Ǻ�Q؛�9���=�H��B"�-quU �S�ƾJ�B�e0���v�V�[6��nH1�j���	R&����ݷ���Y*����b�ߓ到G�2��/�$S�.���A�D�E+Q�',G�h�x���t�T��a����q��Tb.�n&`4��#��>��hGS��!��ul��� Ћ���I�}�:V[x4x]��Q��� ���'AE��@G��B�C6�! q]�v�,lv?f��nU�ͥ%H?�Ҥ���.�-�� �h��,QH�X��U �y��jS���U�%ΰR�b��Ȋ�._�7��	B�Vm��(����^}ʹ�tV`�h{�1�U��4������T�Z�BI��M��+�El����g�G�u�Y��� r���(Pq�/K�V�%e���Ԟ�D���s5Aͼ�)<�%af�;�;���*�&�>�3T�\�
�o��z��ET��Ζ�����k�\��x��<�t�M��B������h�%!�	'���{,"s��ҽ��8��[@Bdb��t70%u�z@`�s���1��ݵ���=�t�Q��E�?��F�x�~�u��
-����᭓$&���A���Ю<m5��3��=ˌ����(�BR���J���^�X=!�	�Cl�K�k����3"�a���H3���I���ꦃ����uz��''Q�9^8��ǻ�h�=�5�H�z�-�}�����-� ���Q��u�y<ً"��?sI+�"� u��	�	��>�;��@��H�&rz�����|W%��$囍J?�AU�P��m͖��g~"8�1����>�+}�ְ�h���0@��F �p������)��J�{�Q*�"+l�����N#_�ue5�D�~�iۗ��{v�b�dY�w��G�5�&Hŀ��V���{�x&Ō�ל���]��b�kz=N�SYl�6����Ҫ^I&�2Ȟ0H�	�`��h���������㊚�MO3�}k�Sw������ʦ�_ԣ�_�E��f^��|}�q<~iw�].�p�^�+��������_Л�o��CurB���l�A�Cf�I��'�;����B6B���/�a�8ߋ���|˴|������u�����t`ᡇ�;�Cx�;��Vj/�q��gXga���Ě(��@���Le�	^W3����z0T���va���i��CYJ��2�V��eV�&���řY);L��G�3�ڧrH��2����4���<�Y�U1A�lZ�}/��ic_4P�A�:�R��KJ#���jYy-�j��F�^��KY�Ǳܳ �Zm��(��1��w��K�Z��T0�?�<s�r�d�[:�$�"-jɼ�Ya]��ƻ|�"=n�i�J��Pٍ��A�nn�_��Q$� �mb�������/&�y��2���/$q�����%㨡�!��w�� �;�C�~�X��%���ܘ�dT*�E�T��j6_�3�H����>c��F��(�&�}K��g����WSZĈ	i��d��Ct��8�*�h�'�&0����S�}�$?d����i]�Ik�b���R�|�`�Hs�r�+����۪����j
��W�A�J�OU/�&(PF��ᐣ�XAE�����3_I��W�:4��-$���mN]6�@�ژ�h������*�s���<qd�U��U�v�4�U�N +f<�va�*��캚4/ȳ��������:}`�%���1���U����4f�̾��O]O�Mt�s�+4mcXȦ��T��D�?��.j�kF<���N"^�B1�Sl����/�����ӎ���n���w��Ǘh�[^�<�5S�_��w�t�&���,V��6�ma5�[��Exn�����/���6�t��[j.l����(11�{�8]�޹���q����N��A!�nvб�<[f�IۄVqׅ��{�dQw��H��%5��(���Ȟɏ����N��#�{"��P�m�y��P��Ay��87�\�{lO
~G�l�!UO�0��d'/M�0={k�3�u$�]hj����U��F��?�D��w|��}�	�������h���~^���s���Z��wD����
#�&�+|Ϗ�kۖ������fx�R�"tʕ�U�����i��V8�˽���͕��q�UЮ��-5�n�ׅ�D&E��qG�p�M�����eMĻwԭ�/�D�-=c%�7 �ػ�gj����m�f��Ԝ�΃�室:r�ô�T0��+��K�%B�O�*����̨��;7����k�Ɯ(�OK�BSc�2���A�!�s[�|�g��GT�����/�*!t�D�5�n�����nJ��7+�Þ��}{���]��������Bw�3�P��7L�Ǟ��"
8Q�����}�{s�J�0��q�`�72ڐ?��L����	�hrC�3G��zލ|6q�:A�oJŃa�w�ZR���m]-�b�?���ű��V�P�C܆�a/�}Q��2���~�!N�Ī@5��᱈EH3��<VX�q.�797��+�<Ȫ�޵C������dU���a���op�*b��d(���L�VL�*4�h��	�.�2�a�Q?'���{e��^F��S��ZR���<G���!P��,�a�T��8��o���:���Q��Q����ߪ+ ���uA"��B b���� 7�����Nh��^��E}������Vr
����y�ć��e�>p�h<	45�����$�����Aa�q��~f����|k�~�z�o�?��}#���Wwz �ԆwP�Bc�:��/2��w�?A%bN��.�b�"א�1��.m�%�*���.�<�c�$�O9�'ja�\�몌H䕵,s���Yӡo8�o�J��x3��yj�5q�v/�Ƞ¼aOP��ِ�G6�Fs��-Z�L�!_�L��	qW�?�q��o7���t�E�(U+�y<^�DuR|HF��,]��� �YK�W��N�eZ�~�n����$(T4�<����R��0��⪃�q�Z��P+gǨ��$���V�g;ށ�y�~�D����{=�U%R��i���H�%V�z��跕���z9:~����z�d��\s�ޗeR`���H�z��#2�5&Z�/�@�-B7E�=�Ҏ�@2����q�Zc�𷀍,m�=��<��e����	W_�:A,������­�!̀C��w<[Wv�l5�G��:w�+4���g]���i�r��eIqm4+��W�^��}�G�}I��~����I�9���kU�]-Ǝ�q�)J��_l��m�z�?0��t��o�����ns�?9����K��L�T��P�˷��L+������z�suNZ@�s�~i��,�d��"}e r� Gt�UGO���Xh\��eu��?���W=vW�/.��e�iƟ� �8�m��"~���
�$�j�9
)�!�jxI~I���+oVw ��މ�'n���I��'�Н�^��Xu"�P+�#s;T�#�A��t��Qۋ�<�UW h/�a�;Bh5ؒ�7���^���R~�Q�|� ���y#��qY���;X���;Mٿ1[�g\-�%<�aj�����,�x��C�	��� �3k*�w}#uaa2���/5m$��`��p���b����}t���=O��J=3���
9�e*��H.]k��,�����6�7����[��0_1>FU��K�Sc��:a���KB5z���L��@�.5	̪EC_�J}#��v�fK9̄e�A��ǋ�߶'�,$[�۵N�<���ʩ���4��D!��@7
�֌>S?U�h�!H%yu�T�}�?�{�C!���ج6,0��@t����]ݒ�-�����`�2Mۀ͇��g��u��6�MA}CI��X3���Ȼ���6���a�����oGH��m�R2U�p��'�e��&&q�gzM�i���>j�X1�	�>���7P1��˒�22��`X߱�
l� ^Ңrf�5]��.]��(86@slH�ظ��*�YO�$d�7;�e��w^~Z�99"�����>�M��'���M`\�5A�q$�[GSA�
�2��ܕ�S�Nqoݪ�B�<��u.��I���+�;P����馄��`�Id�ެ{qH�:3��T�z' 
wc�pA��8�.�uE��;_R�����*��I�����;�ln�� ��؀��9`�"/U���7)���=_�rOK��G��@�A6�ŜZ)��w���#�X�ZUfq�����p��m���'=5�|�Oa���7+�\��ۄ�������X�pCNd�oP,�&�m,����6�QG�Zc������伺�k ��If�-~ sw�]9� �㤦R���!X�]L	�c�H)�Wb.�:���ƍ�N"7�gB������uGCc!��S�?����@ct�^�15�r�M�`(�s��z�����QO���9D,��q���E��EZ0^�$���퀶@/���K�\Pg�1t��dw�����ƴ��:�����{U���o�^�H�dzPK�f ���U��>�o�`{��:�4�$��z��ɰ��RĽ%)8l�_�ۛ�*eϯΠLu��{g�1=Y濇�pǘ�#[3�4�X j���&q��HcC�_N#7���{F2W�ϋ���#r��@�M)B��@���Đ�U�
�m���W��S���� >��I"v�l�g.�������HV�{�1|Z��&TN-���X���$¶�ߖB��܈xj\\C�N��J��4r�N� 2 �5skH����m:m�����KNq�7�C~���f3�/����*��J��YN$n`����f������$�Ecd���ۻ�V7��oV�Vj���j�x]]��t��b�_מ%u��؈f[b����Bǥ��t�1�I}N�&b"~_�� �&��X%Y~E��p����yMC��!�cj�]�vw��NA޶Py4�l�/��|I����;���TPZ�,j�&�k�2��P&��}�k�5A�+��}�*YmP�1�V�����C�͗�ʚ��i	-[�2��o�շ�h�@���Ƥ{h����y�Ӧ����I����>�4_�?(n:=6l�Rbt.��C�h����5M��p7��wg���(�����V��|f�/���ZY�H�Ԃ��=5�K_S���2��?�"�_�y$v���h��7�.^B8���6p ;BV�Ԕ�{2�y $Y�P�Ӂ��8��qֳ��ì��G~n��k|�&��0�#S��,�]?n��g&�ѺH�8�Uf�[�M����W�����D2��"�����0�Nb�������ݏ�E��U����!
���VB_�cCWu`���)ިb ¸}��6Ԡ��j\��3��+뎞+�����g����f0<����oa���0�-x/��q�H#C���0�=F�e�?�v��.��Ѝx��QbK���|�C2V����ZH��� �9�ES�T��r�aE����O�R����dZX��,�0�ӹ�AU��$��iTǙ��#j/���e/��gֺ%:Lϔ�k7P`Wg�i"�� �s�S1=Ob���%Y��y�2e�ַ�6�L��`X�F�a���������N��Z��P��Nx`m�H$)�󄕺�X+S5Z<����:4���6�}O�f*�a=�.f)Α|�?A��)f��6��SD� OpO�A�:����ʹ�Y�\����/$,�@�����9 ki"*	�����$�k��+�m���|y^|�^4b�H�k����%;oBc$_?42B0i%2=)_A�H[]L`l����� ��cU%^$�)�<>�ޯ��PU�v?R����C>1m]#B�M`˸2�+KyN����U�a�4�N���[ey�^;͗�SUe�3b�h�T��;	t�-��<��� xm�+��� Bƒ�R�V�����;��^�-g[�{F��|�w&;>_�	����M6,�< �)�<�K��,_���Ք�J�
1���#���P������d��b�*AʘU�aFf�<V^�
S��S|/�G�{+�6��q@n��M ���l����j�^,ok�䯮�ʘ���v���Lsh횽�j��/��dY�nE3g�."�"w�z��v��*�Z��%�-�Nٮ�wM�dy�?��ܓq�/ĭP����|� ��P`�|��-P;`yX�swƢ��^)o�]x{$�T������N;B�Ɇ��WG_�h&�WR��C�;�A�J�l��<��K<�\9ZTZ[��.	 ��C�1�K��s�����I�=QA�.��U�k�y��	ID�Cac��!��#�WAOP1�p��X�1���
�t�A)f�%D���*��Z��r�[4�J�#��3���ͮ㩄���_Zc�Ye��m�"�XyYl	w>���5u��2�0}��S���q.!��'��? <�?^C���' �d�5�b�����p�x�O X�q�s��#���Q���p�����Z�tuw��Dj�`l�˅��A��Y��9Ɛ�����Xc��ڣ���7
H�%i����<ZAm�C1�rĭ��9��I�=��R�c)v�:P�dƥ]J�ڥb�H^�>b^4���$@�#aDۡ��K	���05����M1ʆ��X�`H����D��c�z����Qt�����컚��_��������e--e&6�}p�~`�J�:S�j(��~�?�Z�O��eE�Y��xK)��5��G;4��۵����|i Y�*\uE�q��븉 �D�Ck���V��G�֍�{1i�EA��ܱ���&y�8��pS��#�1�q�:)`LK�3U8��oś��n��	�r��i͖�D�|J��V���?�=sGRi�;���"vJe�Q3�2"���]���#�����qy%_�x��v��q�y�fƸx�#]"??B��8��X��4 mZ,��&�䁜��e�!f��n�規+�=�+�Ҡf��}*�ev���xEP?y����Y@�P�o�	�w�@��Q�Ħ�Oi����d1"\%v�kղ�q�Ps��mF0���4��"5�d)]���*K �t��R�#�0��P)m\Ed�������P��T>t��@�������O4҉�8��R8��p�����v�ΰ�Ǹg�	���l𬃳�'��elꉫ�p������A����/�-#>R����r�3�E[M��>��$����{>,_<0��i�	���}Da����[o-�E�����֐��M��\�(�q��t��"�G����^�ᭈ��(5:Ѻ������M6��=s4�3(��WS������4P] ���L�<���r��� d�
X������̠��Ť$;��{ZF:{�ݩ���4��[���	�Qz�}M 6i�u\fc=�?�"M��	����v��1�aT�	��k��]������zX=����~,�ˢ{�yȭc)�I�5ŶpQ?�l!�;�rL*�����*45�iP�����]`==����c�S�.��;w���@uC���j�+�&�M��YO�C�Ƣ��77]��x���6f</�6�K�bW �3�t�9"lƿ��Տ|�R��{ �e�Yl�:�m(�W��*GK  �C� ���)y6�|��������+����?3��6 ��xrp^��J�ߟ&(���\���D���1��g]9�wqQJ��+&���K_Gɓ�mC��[E�pS��lJA������ѣ�KU�:u�:V���Y,��V<p6ö��j�0{4���wS`�D��r��-���Q�̥A>[����=�[��>�������Ҵ١��X�!���������"a�Ē��DaT�fEާ��� �UU�I�w���Z��Ƽ��8�S>�Kk�@�D��R���ļP�{�񠾵l	2V����b�0T$=K�@A&���W� ����\��b�7�����GI����?j2T��S��x��ﻭJ[NV��+��R�o���ŏ�[*?>�n۫�����C؊���n���J]{Q�5H�҇� �o)6�"��Z�]\-��� ���¼O�b�轪��\�#:��t��B	t��Rpb�b��=<�uR_��,�IK�}!Yw�A�$��搊�����<�X�Q�E��Խ��o+�d��=���Q�ŌQ�W!�y�М�	^*��G�b;��bY��D�V�}�Y3��qM�e�4[�xZ�{AQ��l�<ہ8_������sq�=&���:��l@�ۯ~�������yu���F��,hqmSUS��6�ڰLSxCuϝ�hQ��:O�+U$�X3l�XQ?{!��K]r���*�z@|�碄6�y���N>��4!âN�t?�*�?�bH������
��J���1y$�dl��,1��I���r��q�x.����^;�P��('8Y��\�):����[�� �kS�H�	�T�~�jDE
�<�3h W\	;W���O��ԇk�e�Bc�2vS���H�p�����谄m�
�di:�}Ó,�}�#�|ҳ�,�*�n��(f���QxX=8����+�D���3��A¥4M�;�V�K�
��&�_�75��5�j��	W"��TӀs}|���鳓�;?���o��0&/��0fN�%D���X�[.=�oSՋ�I��/��k��ee_��%Ὕ��>i��t���,�$0+��H��M�O�ԭj�~hKXA�`^*H��nVl9:C���)��*�R�y�d�`B���.eLN�e���ͨ�r�Bp
�RyaȒ{g^����:D�B�b����w��n7|Ü���
�H�;�W�P�4�a��]c�<3��G����}�] �׾Ls��ˋz �� �d����`E�#��1�P:�\�[���?�)x��Nˎf�~�k�\!>hQl�p+b���w����-��W<���&�$�u۶�a���22�S�ۑ��x��aO�7����~rs2�Oi���J��F�u@�:/8ڕ[|	f��S�F�讛M�!�~�OU(����M��*v�t����MIDm�6vH��Teh���5�oC�#��N��ԟ������քU�5����Y��h����"ԍ\)�8O$C�ϱ�
!}�y�G9
��p$�p�NN쑴�&l�f��-K����Ǣ1�)�ͤ�Z�W�W�b*Z1�C���qc_��Ǘ�l �f��U������Mܙ*��N:pI%��kE�dO�%uB�@+��W�c�Re���|(owB���*�tiS4�5X�4S���K*i�wi �W�����'b�2�����W�
,��UH��% �*vM��t�J7����ɖ���sg����F�%R&<(�=�u�d�@�F]�I��� �)�7�G�,�ӭ�s�|�S���T�B?�e�Vݪ����z��G�P��J�������f�q���xf���c(�Ί���b,ݙg��n��Љ��*��o2��q� dlU����B�5܈��&wa��
|#�G�����#`�m(�������y�_ǿ�t.�*䐊?T��AyOjp�^���K� ���^��2�R��ɉ=�:�t�#����h[�@��Y%���۴D�*'vvrwiS4Aͩ^`�{ux����~2:����[�����2����G-V�H<i��f��b�}cR���<�L	@��-�y7�Q��߷/
�ےR�7��X�aI#��f^�k�� !H��Zqw�t���[��5��[Cz�l�%}�P�����NH�g������訇�[wf���k�2\WK�\Y��ߌ��u�,VX����/��.�+�+(f��KZ�n�T8�y�k�ƕ��Z�K�R�~j����b|�)<�Mlʘ�U0�PBv�O,S2��ܔi4\�$-'������� �n�[�t=׌B�$��r6�&x��4���a9(O+�6�/n� �M0A,�b����� ��΁]Ø�L1���H��U�2�Fh�`Qor��P<���8pTwΩ7:�	`i�[���ک>�[S^@"��%J����jIpO�������� ��>Y:2no�%uv(jJ�B����\��>q�mR�$L�d��_��3���\43?cD�9���6P�_Nw0��4��w�A��{$p&?`z���aTc\�q�\}��i���Y�ԾSB�hS���#��4s�-И�B�(�ӏ7˯,���{w%�fik����Z]�?��� ���&V�<�-���O��Y�?����p�_Q7�مE��țc�BN2���^CGQ��T`�׽��Ju@j�v[�+P���j5r������r�rm�A�H*<��P��9���w3��{�.U�#������	u5mr/�_�Ш>�0y������;�f)������ޒ�ȤA��K���3�w��y�~㟢��u���*�ܶm��L�p����۬�٪I��e�kH9�����_��0a�����Sk8��"�(F�jA#tODW�$~�Ks�Z�2m\�9��!w�$[ҫ�S&�� z�����6�t4&�����'?zͯe"��;(�\F����]M6���2����w���B+ä,�af��=Gq��Y?g0���i���9��0Wh�<gXq�=����9R��З�R��ݵ��=H�=��q����א�@�_�&��m>�����@'G�D���,���A��&3gLFc&�}IlQ	���ܽ�;y����Zr��-]��Y����G�'�%.� F1��Xe\������n���f��Q�,q����M(\p����x�x�����C���Z�o�A����AN5��� ��/���	�9z�%�p������N:��L+�#��֩Tz�&;������V�N�IW�qi"�Öa�g�8X�N/����7���~��c��Lƾ+�I�i��;�E�E`�����e&Թ�HDuS���r!��K��P�<��)F@S;<q�-�8�wI�7���2��L�/J@��j��[��x�^=s~O@L�Lcͬ���#�}\"Q��>��s!�Y����N�\i_N�da��,�a睬��ލ礘�6~`ѕ;$>^�ڪ��8s��n�~b۪����+�hߜ�xPA?�~Ƃ.��6[6�<:���-6?����'&���- �B&n\�=͞�iA?����C�6J��DeE�A[�4XIs�X}�)����$�-��y��<Ҥ#�4�v b:�V_u���G2����"T�Xz�MǏ�i�ZB=�&8����Xo+�n极��]%��ݓ���g�Ȇ��	� ѿ�y������ʾ�~������aq�	�[N�����^K�$�Q����@�	Wz]����3R�}�M�?�v_|B'G����K��0^�{wd�����\W����$����{��/�Ow��*AMdj��������d���L��
Q�bGg����CG�8j9���0Füu[�6�"��2ܴ �E%��	��N4?)5�`�(U~�7���D�|�#9��Yw��k(,EeE�H��:u����&�m�<x������&se"<r#Y�}i;�G��U����e[ItX��.�Q.iNa�j�^9+��fMj1W��iQ)C�*�>z4�V>|8�R��Y̍(N�-kj�J��b|c�B���E]�zQ�^���|�	#	�jK���\y;�$I�b���krj�B8�E�Ƽ��y|�.�!��5;��Zo��M<��dh�\����x��+h���e,L̫��2����h9�1>��:t�a���j�T��5�X��u
�c�P�X���ڳ�o�.ה@>P�߀����,ED�yN�G��1����&ڽ���O�PH��s��I��7�&���|&7�+?҈�)����T��}.��>�`s:?Ɂ~+��XO��E�m;S�q����4�7�=r3��Ah�d� zv����?��o���w!����%7+1�4�h�I�a�do�&�6Kg��K�57�3���6p�RR�����fW#�M�g�]�!J�uj��ͨ��
�j�>#Aw&�!���)�t7��!���me�ۼP�O�2]$��[ � �t��bV��¬
05�QPL�7��.z�*m�J��jx�斞?V��}/*T(ɩ��wC�Y�w�/�;���ɪɊ(	�$�I8������?31��ćo�3sgp����*��?P��=�E����AL�z*F��O��Ѱ}��#�b��!*�Z���ɓ*�r���	XK`��Oͽ�) �CثU����o�;��gĻD�K���d�R��g���u�@AF�I�wmuH�2h� �xj�x<����D�����\�Z�ՊZ�s<�ۢw�� >��%��6��{��<�y����vQçk�Z�z)�U�)7�C�"����Ŕs'pf���{�g���M/�4���{5���Y�G�*naN�	�~{���^��� 1��"��:H?���yO�3�����G�<�`�l�ug:��y�Zq�)$�Ivv�-0a��@l3�Y_�{6g�%��*b�<]�x�k��#�^���	��}��R��^\�]t ��V�oe�|��������C-i�Q�Ft:�ׁ�*GSj���aFȲ��|�(L&ɲ�wZ҆�R�Ě��1z��bLƙ���
: gDT�k.����]P?X`W0�ch�jJ�����=��7��Vmt�\о/e�(T\ߤ��߷[�x���N>d�Ӥd��׺�Z*p+nhӾ8�&7�i�)F�ܝ��{������D�ֿ�S��]w2=颣̞{[ܦZ����8DU��֌rE�1U����3��G�R��s,�$�zD�;����Z�\���K�.-�9sY+	����vzT)%U%޻񉏚�4쥟�됒 L�+�{(�b�?W�o�Vn/��LT��C� a~ׁ���eC ep�O�x4���(�u��%%�{"O���4kXV+L4��S<<�����H��) M*�X�}���#[��!��>9
��O�����76&ח�1p�%[�
tU���5Ő�̏@��9U�e� �D�R�z���8�Z�)�����F� AQ�����:N�����7w[�S�N}��NܮSF\y�Js S�?6Py� �K��f�3��O���[}�Cl~l�R�~����M�W?�%�#d���m���ț.)���sA$3�[����&�à�(�h�r�'QO�I
H�5�|^i*��b�?�4F�$���4t^S��I��5e��j��_�u��YW���tW�IL/�&gZ35���&H�ebM��ʳ�8��B�nDHL����u;=}�Ŏ��U�T}F�z����!Y�?�SzY1���(�r5�ұ-���~{���㴁��֊�wY�{b/l)1�nI��=Q��W!0���0X��#�V��a1�%�HLb9"3��ƪ7���`��7Y�ۈI�HD��5�@j_�����J�!O���}��"�nϛ�C�^Ve��`�����C��2J+%���3r{Z��΄����ԱT>�ݿ�(!Tu���\�(�N/r�?+&���Z{u�%�t��[m|p��@)�;x��!"<!aˡt����@���d�͎Nh���k��dg��1������̕����c�Ϸ��멚��V!��.j��҈��f��e�@�D�-g	/���l9Cì�ڕ;���Ի^E��K��J�$���ܔy����*j�U�HjVn���{Q�D��0l�����>4'�b�w�%�'=ڳ>;8%e�P��`U�n����cG�����]�ډ!���&��wx}H��%E4��46Z�Un��եbq(����k&��d]�ܷ�u^xɲ�0�<�_]��1�`���_��8l>J�Q���ѱA�g3}x�>ZͲ���,�z���mT�}�We����E�Y����zE.�� ����`t��煇譜�P�+5����V ��3� ��;q3?y49��g���l=|���%�����0񓲉��4j\c�9�� �z��q�Xw�q��lR��	�e��a����v�t��4�;�0EI)vⱬ����Iʇw�w�����|,�C1�C$�wK�R�Ќ�-n^p?9-�DRH7�H//�)%&q���+��c{!��ܸf�\Y�3J��������g�ؚv�U�����/u�=3��&�b��.z'x����,�[�үK�a�<�U4t��}�Y��r��+5���h.W�����(RG,�p??)�X�t�����]�>��i��q5�4��4~�ɊS�[�)ξ�c0���r|&��#���V'Fuu�b�Y�ԆV�8���,��=P�?(�匞�8B�Oni����c%g:�#"YT�iZ@��!m�:������q�V���d�R��:s��5cMեtqpU��"�,׾½����Q��"4���\3ʁ�!ڃ��mV��'lHpnו�*���H|D���4�p��((%������۾X�?��G�l�ZSS�_�Y���"ǀh9GC�P�*���l~ $M�B &tqF%�s�c��_�F��>K�jT��Ŋ�eA�/���D�m@�̒�9D��D�c��r5A���|K�*v{-�]�}Aпdށo�[���%����r�W+Ē܍�P}��i�6�,2-�P�H�0= ��
V�<gNP���6��-b���T6C�tju��,�+Rcz�V�&�ջ~(�|,KUѐ�#l�5.9��lY��T,���'�(�ͮJ�m��D�8�BC�,�}��[���C����pH|��i�O"P���l��Uj/#���x��u��o+DO�,v�\�d3G���Y�A=j�Phz���ar�̃���g�7!,PK�1���+��E��E9���	����G �Y�B���g�#	ޠ�o+�n�~PS.�'���۫�s3k�����1 �\���i�E��o�:4r�}Q���M (�����eR9 ������n���g`�'�n5T�iHԌ�H��8�k_�}7i8?��u���l��:+�i����}�����ۥ��8�=�݊ˌ5?/=q7*�����D���<Lҫ"˵��}Hּ��F�)��u�E71��Ҡ	�M�kZoL�
��i#x5��8�L�k�U
��0KJ|�4ن�5�.��t؀��hq���?!�)����οඞ��U#���]�FA^u?pW��c ��=��;� g�]�1G�N�%Mc����L,����E��Ӹ{[܆nq`S�g�-i��u�(�M�����Y(l�\�M�t�c/ Z��7��ҵ��:`�5y-�>V�Zm�/w�8[�:����LÞ⹈R�1��	h�Pj%j�<b�AQ)������x!���<�J{�G�ۤ����?8"�,4*Q�1�dG�SgV�T��� �����L�2c�/Y=K���k䛹8���?�����g�s��h�b$ �H�X���>h��R�Vy�L; AL��f�?>m�nu�BW*��ځ���h����T0��y@2��t#m8���0hZ�[I�)T'�P���s���}55��
�V5hbal��!�~8v�y}�'�W[����Ly �F�S�VT�����e�&�����9�:6
��pɱ	�kr_� ߍ�����)6x�	�w�I�5u]C0қ���{�����_PN��/+j���hLC	��[.��Sm�Eie��<�5�W�5�03?DΥ ኘ䠬�[��GEvc�n�}�mȱ+�yaf�C�Pg�䗈��Ĩ ֠ZXq�a�F���l��f�f61����O�F~�!���x"z�BD�		2���!,:���X�{N�!��AX�����B�s�ݤ����,m.%�us=?������n!��C��A�˼|m5p�т2S����'�K�+������R�D���#�z���zÝ�3~����f�p_m[n�|`��
p�B�C~R�Er�Y ߟ�}6�[�z{f�~¾^p�A���ŊSY���n�LϥkN0��)�;�� @�e%s�a��Z�����.�+�g�	vt�~��.�C(�T�v�2��,3�N;��=��B��h��,�-2�ć6�U���i�W�gW���1����c+'iŷ����P�邭�?oy\�f���C@�\���OĴ�g<���	ob�x\��gH�
h"|��al`g�֟�a����ӵ�+KV��8�$>8�oz�%��~4<���3'���M%t>�����y�a\�u��2��B_MȎ�A�n�.U�J-�dv?�u��}��^�2��6	��Fп�yZ-�4K$t&Ji�i�"8��m�	�Ug<��p����!�H&���8l2e?AƖ��R�N�<���}ٶ,LmuK�`E<:xح<� ���O����5�saj�E�}y��hEy�?�j�y�.�C���t4���]����7�8�K�B���=�7>���Jі\+qE8�V����Do���+7�O\~���2���<�jWk2z�ɀ�1C$޵�-�m�0��\p<��Aw�U�ǈ��[c�#Rk)��J��Zn�'��7��"���1�^	X���d��'�p�����$��H�uC�`?1��O�QX[��0�44�i9$�Tp��>����� ��aSԦ��P�H�/�O�/俕�O��q�F4�Y?���5/rD{.����jh,Y�y�a��֘mDg���#���	�v(<�X�F�I�2�*�����T������|m{� Os�o/�G�/�@�#��٦-)iJ�T���潃%wo�?v���kym��|���	�S�KX_��D��w�[�yJS��4%0��֏�Ԇߑ���+C(MJ�
:�C� c��j��ʹ��.Sp�;[�%O�)� ���D��� 9o"��ؚn�G�ի�^m��g�j%�Q >�H �!�Rz�NJ��rV�iۂ�D�b����4��)��)��S��G�Zdv�� �?��e���:Q4��<�"�M6�̤�*����.}�����[��?�x>מ�^ 7MI�����ߞ!6��iP�>}�+
�9b�X��02��G)�ouؾݪ�M�����&M5k�+Þ
m��}�Pz^������|�npI�bX@�v)҂�mJ�2^�>�<���n�*�Yr̿��~�	�f�����7���e�U�@�Y����e� w	�m�!$��y#�62���k?#UР����������m}+�����(�y]�ܵ�!�M����F�tJ17$���-pE��6)Ѫ�9�ׅa���f��F����`���(`�-E� �����G	eH�� @�����U�--� �lTL�j�JXpԭ�������%�Ð�v�iB��{v�El%��Ɋ���i^V<�7��#t&$xt*yj�{?���{*f�O�*WFu(�coE<��G��Jl���B6�m�����EK�g�[0h����³����!��0��#j���7,%U��0+�s-F��!88$�[�^��uH����c���A�U�H�8�٘� v&-j&4�YpJ�� ��L���dU��-R���B�*��v\����5����q��׀/��r�H8F��J�?xMjx�w�/�Ϳ��WM���d�/_��^=s� 
(&O3���g9F>5\�p��{P���Q9q�#�_ܸ����r-��)o�z����� �� J{�b.��1NK�Z��^����<J�Lx�;5=��H���sO�x�'���c񵢓�aT�.����&~'�9�0�zQ������CJ�k=���Y�[Ɋ>���� 	�@E���dT-&���;��zåF�.���}b<���+r//�m�D9+jx��}΁�����s�Q�tiP+W�h�;�X���(3��+��l�(��'�]ɦ*v�cP��y'k�fh����	�H�{�������=�务=�H��Jí��3ȱK�hYǍ���7����	-��V��!�'T��l(�*�)�k��y��fd�M��$���N";yݞ�\�胄+�u���14|��lT0A�A�VA+e��:q-4�\3e�C���3�����վ���W��+gg@����S��R�.8{G�?��f�]8�\�A�fZ�ئ�S,|�����I�h!��leD9�  ����P���T��nprUv��(�J>��ɧ�q	�L���a������D��[�ؚgjW�r�y�@�D]�: ˻����ʻ�a�])LD�U�Q�5M11F�P��{��e����:�g��P�`���_;V�<Xb�T�;�݅ZÇf:��¥�%�8{�=K���9q��$���/�a�_�v� &�Ru1�GsG�)M�Ph�G��Y�A�SM����=Y;z|+���S���өQ���͖��|$o�A3���)݌x�_�}ce����u0��H�E�Dn�ϧ!�J�f0�3���_H�n�'���f_��������U�k�#�)t����\^��P�ޕ.5g�Aeb)[o���2�ُ4���r��O�37`�Ս_��}̇����OfOj�-u�W�TTH������s?+�C����N5&��^����R+jM�j�<a�fW��^ȿU��t�:2�����:�2LY<�Yk��5����/�� ��2GF��5�H�ۈKU�R�[fl�w�ˑ����?��rcm_b����`mx�=����93}�@p�.��BR $/[,#�Z3�)�Dȧ�b�a��Hx�|ۉr�}bGgq��h-��\���%���Qǚ�P�VEP��Y�jw�����;�NW.�������9�醱ʉ�?w�}V�aH����N��=U�t�K	�̪��9Qyo4T��X�Ϗ�~��ǡd9Ry��=�p����@��@�z�����I'}P��g'�w&!餱���_ؔ��H������K��k�$)n��:ퟱ�綩��]Ǉ�)����=� i�^J�D�j`)$n0��C��$T�,D:��!.�[�7	�t�� �2a?}?�+��1�ƀ{+�O�)��Bbf�7��j�z�fY?��A�a���
���>��3Q�?$k�sw�\̣(O0'��|������<��4�]���U^& �|(%1����&�����+K�.u˼V�w((;�,O��cq���-P:H4�G�\S�Oc�
�A�ͯ�I��T��}%���m��}�=.RV���AX�]y�9�p�#�L��I�m�����5�ev���f�r}���>c:(�XTVp�BI�b����U[�j>A�M!�חv��Y��!�,3F�vf���-��9G�s;�e��\)!d�ǓX� c���n�	Oͪ���p����c�k�d��aYܶ~��y]�쌭���|��A���I}�5弄�����V>J���!ߥU��md�~`[����aڻ���-lX�����m�Rj�/�I!t�3��� ��0��w�R�W�k4�����M$ѷ`�~��*��� ��I� ��%BJ�7趃|�`p�^�J�S�ʋ�����'U��C�y؋���y���?��p�:zUIQW�G�H/�����-��ނ,�oۆ�����f8!(�1�i�o�����*��II?�=����,k^͜�g��5��D!�+U�?z������j<<��~����0�S�{]�F�_���x�(B�\���鞩�k�G1jG{cr}��b��e�WE���	s*d(�X��jPa���Y��r�f�����S�#�B���D������������Gt�ݿT���<�Rg����M�9 ��H?���A��}���G�m�:ņ4-�~_f#n%���x]F��h��+��cb��[n�pJ9����5�0Nn���/��9+(�����t4�ӧ�X`��8Z�R�c�Kb�xB�T�`���O;"�λ�x+�(2IJ�z��u������vM��ªZZ]l��#����DCbY&�OWC����n8�0�Ko���+�t=�z��$	��Hz*�8��}�
ʽF����E�(�M�xA2V��*P��[W1�2	63ϳ��Q
"�Ae��3%)��4����ϊ�[~��RQ���p8EѼ*ű�3ȳ &���xD��7tt\�+��Ua<8�~>�?�$ S�M���Y��S?��Ct�{��HOs���>~V��kI��w��;h%�^C%�%~��a�Wr���P�m��"���t�#G[�k��{����v�YĶ||��e�c���%�s~Fk.�ɩiZ���Vλ�b�cO6+x�I��z�tC�]Y�Ӊ�Pg�b[n��sځCYC�w�i�̹�����4P��P�]J���1�2w���;�ܔ�y�����;3C;v%��M@R�=.1����]��6�xEV�:/;y���`����u���)�j>��!�K��ߔV�6��DcÑ�\>��(�O�M�y0��g(�l�g����ގ��ݑ�[�A$�P�1����������3|�7^�sK�Z�!��JJ�T��]��p��#�h&��j���E�1:g���ҿ��!�H�#�OCK�e����M��dpF�)P���+J�S���	�q�]IS[[�.�{FT�B5�<o�ץ$��j�Q�{�kb���I5�gﾮ���k@_�ӆ�'+�,�5��5���b(��|+T�^�������@6�$>����>��_W7��B�K�Ɯ͉;-�ae`�u�_z4�2�z�����gc\t�Q��&Qv� I`)/E{z;�����,(��y��շ`��@'��~��	i��YE�K:�:����;�=Th�� �YWf�}�I��8��q�~���Ђi�kf�!S���U�Gw��|����yw]�-�K�i������#� ���}��%j"g�
��K4���L�W���E�w+!X���>��w�z7�Q��~�O�8����*�sz�]9`��l$��e��Ac0T�Lfp�~U�L޵��M�8��g�,����1���_漄ޅ�Y���AVi)lj�%��u�]8�6��}E���M��A+�vY+��>�j��ҏ�|?g;]����b2P!�x~S��UȥS���n�8e�3dV��V��m�i�!���<���֣�tg#�����?��w�ԡdř�xEO�dA�w�������y@u"�7�n�S�m٪)����Y���w���A���̷�՘�㡩�?V��ӧ�F����Ό�6Va��N��� ���ϡ.1��V�a���]�e��ϢC��t�YCM:E�M�]�,yo���`�05��0��𶪐�����Ө�A���T2�!D�y��A�-����N�
�y�voV�ۭ�k�M��t&v!s�ɵ����[0�6�R�H�����:s
֎?x�賦�]������ަ��?~�0��J�𼆱��n��G��j\���aw������ź�����A~��Ub���)��.q֩�:_qW�B��L�-�$�����Z�ɏ���=!�Îm���R��~@3%	H����u�Lt[~�JME������OA5�ؿu��M�qu�"�Xŷ�T\I����ɭT�W��l$��AW���jo���g��3��jg�fޡ=�c/�+��ΓCa��i�wkPo���a�%��|pX�	�Ld �7py�3����§�L��9��ʿd��o!$�������.m�3�.��	�`�?c�!Hj��zՅ�G��Q�Ee�����?m��'O�p��&'�N�x�NM&By�^��¯č*'�Nԃ?D<[�Rb҈����ԚI�/�y���E�+�} T�;��8i���2\e�Qχl��Bwx@�z[������C�����C�& t7��a�Gtq���V�,5+�ݕT5�[]����l|]u�eg�$@ϸ9`�<|��TT0���Y�Z�!h�9��2,a���X����71`���$���L�y��,��9�2��ʈ5�Ek��nc��.�Tp���ED��rѱ~�u[P���m3�\�F��GƯ��H�)Z��U9�~��*���>�����aG�m��a��K�O�*8��MpD��%��mH=!����M���3������E���eWKJ[̊�|$�hM*�^*��������4�hw���P2��']�Y�pD��A�c+'H����y!�e��P/��r���5 �Ys�����2�-b�:D�/}���K�!˹�>c�]�i�Z˘7�9�e٘at�y��ߔٿ�p�qKy�L��>.�����I����p�k��:�ó��j� Q������up9~jM���{Bu�~�v�}�D��[GT�C��_P7���B��RF�:��u�G{D+_�����/J9$���!�}�:d�91�Dp�z�.(��*�o�hhX�_i�6#�[Az(ID0����*�V��bR���A��#\+���c^�!�ߢ�����,_���mͽz����M�"��߹�k#�����XJ3���)�ޑ�_���� �n���@�Dd�:d�f��"�n7SVeO�%�n \'2P�%��1�����ʹ���N7�kš�U�5��������5�ݺ7��Oܓ�lK��:P�z�Y���
�i7��������Y�1�[����#���@Y�=E��B�Z<V�*#�Ϩ�:z�.�:,�Թl�k��./��I3��n�[ST5�	�6����w�+���U\��p�b�]λ��v�;*��!����}HO���	���9��|/���
����Q_�`i����W�b!�}�I�F���2N�������^���Y�W�d-�!q��+�@��������MF��em�G�Q\�$��0�"������
���}����o6��C�U1��@���6�t�W3�ݎ�^2s$(������b	��Dv�^ܰ��[��ؐ��4�>�ȳ��<�.���c�ݽ � ��!�9d`6�bAf���q+�o�!��Q���_�*�0��w+n�05%(F?({��E/��,���Lv�H,��hkq���%����F�|+W�O��P0��Hv=M���+�
M�DN��vx�����d�U��*���*D=*BUi#z*�&S�S]�lU�	�`|b��mz����^Y�o鐚&��̅��9�U�{<X��`(�~<��5MZ+B��kX�p��c!v����5����L�a�Ȃ�G#��랫vT�������m���%���T�j�6��tb>�B=���o�ǅ��X���2y��;�iY��v1)�F+�H�g5q�y����i@�ϗk�,y]�F��&�(�=h&ɥH-�Y��6:|�7�����z7�;lTP�<u>��P�9��E���bh�҂��E����2��V��h�<>�K#�ǜb Q~b$�n.�E�M�":	d�	j/=��_���H?�fdX�H	�C��:�q�4T�~M�Ş �e�J%����2C��߀�y����bض�?��ܨi�fڞ�W���:�r�NfB��؞�� �c|~���,��%��۾��-�7��SU^}�P��[��Yos��fc.�ߨ�SMᩰ̅�]�"��'����\�%����W�c&u����"��.ֈ&�������h��H&��˘'��k����;Fl�V%PO�����rU�Y��С.Z��kk�3�P�T6����"x��f�n�v�z�k`*�˱��˚�H-5�����,���e"%ߟӹ�-2��q>_k�\mP-ـٸxlh�n|�v����������$J��k�N���Ʀ7B��A͆g[�!�A����}��b��;�i88��)��fO�I���X�8D�;*�U\�f��K��W���Q��4h����q�A���Ĥ�J0�h�[�$�Q���������L��XP�I�c�c��ĥq���EŻ$�y=� �ePq�	�A�'Jkp7v{�.� z=�s�v2%ӥA�� 0	��@Z����^y ��9Jx�<z`(>Ǡ�qs-�z0/���w.�*������?fv����,mDxǔLL�O!c͌SL4��'pRi��m�p㛀�6�?$�$�+,�5��W/�G�9���\���/3���ɔ]3Ƿ���=�U��7��<�&��=�z�]"���{՜�<�R�E~D�}� R�%g�[Bq�U^H����F��j��᪢��uR�w��ё�Pv�)ˠ%�U?L�:����8̘k�/"N���6�|N�	)�����ʭ/7�t�|�T���a_��T�.6�
<��D��I�{j���9�N�FI�7����.:]�gv����d���\��E�i/�D�K\D5��\����<!�"�!_i�j��(��M�5+�2|m=��9\(#�֝M�b`F�*1����j������i�>MJs�xfP���JZ��~�c�?�_:` �ͧ�t�q^��zw��Fj��J|���).��p=����|n(�TD�!_�a�T��_����h:9t�nXJ��6:� �=xG7�mI�և<"[��
%	n9�ʲ��k\�yC�Y��i,�v�p���k\�{��;"o�-M��MW������񞠩�B
��UP���A.X5�â?�+d�^��(�iG_�Nx�,�{�Ӧt�BԴ��2u����!��Ma
�f�b>�h/M�[!j������\� ���^җ�OMG��B�Ǫ:�$�Ջ��F>FUSbOm��]�$��g���Q������m�E���~��ͮ�م�]���=�/$k|!(P�nn�}�c�i���e��%�����eT�]N�R�I���k*�{� e��G��	{=i�Cb��6����?l��v�X��e8��́�R�Ŝ�#�<��L\X+�G+Y~���m�$��څi�Z�!w�|\ϐo2<�>���7�"��6.
z윃C[�%��#6��m�A���+_`�F9�*���+�y�k����E��E�c���U��Wq�uŽ������C� p��B�ގ���a�Z��!t���CߟNAwU��0��]E֝ϗoHe���s}�5��2�OB�a*��PV�>바��N���.}�M~�W��U�h ������r�t��	SA��	�o����nu��$����9�B���Op`d?.3��;c�+,�'5Tǀ;�/	(�bkH�q����Y�X<\�Ӗ}��VJ�����T��䊯m���\�����x(6�����ޫPe@�Wg8(Ej��&O6 4�����ɉ9ԹΘ?d���"�4zn�,���:s�?�)�P�{#�����˺�a�Сv�M�i�]ަ7I�"sy�>���B�����P^U>$�AG�;4p�Vf�tZ���q#�?T��o�Gr�^4���s�J�]vo��{N枅�T�E�Gf�jl�֣_��2�4}��\j��NZ��6�����o��(�')r,"���gn��_���r�u�c�O����&Ŀ���͠ru
?�B��AWn�o`�G�C-���O��$�S
�^�yV�f�*�2�1<�2l����3ļN�	�UN�i��=��I�FFpi��ɨł���ZlA��xLg��s,�G[�CkE�W����F>�|�4G���h>^����r�E���$c`!!�n���\R7�t�N���d���^8�d��U�Mye
�AyS!���q8_9!^�$z�pytw�JS��Q5}a,.��b`#�*���4�:x�YX 1��O��e����X���k-�7�����j�mt�����<�`ZV B?�h�J��A�S�f�}���='��i��.�Z�6v]!��%)b�<�b���&���[�-���s��n����������X��0ȋ\@@�OFFT1���?���\i�X8���g�fb�z'?sT(�+c���2��ȝ��������w����Z�0E�b�墼�Oek�3�Oogm��G,��fϒRV�@��U�
6�5��;Uw��|��$�_2��%~�ȉi	t����bx��	"t/?u���M���Tc��e%JPz�.=+��)�#�g$�od���ݏ���C��c=����oӢS����D�y�g���� ��®�/Z|<}X.m/r��\�NBCA�����P]U�l���x�x̢ �,��������+vs����Dv�&Td�\�pº���N����?�ֽ 69�Q����|��2�Ár�H):Y�L���Z-߽RjWel[��.�}_���%���::Cb�^X�gN��~��r��a�����n�M���F�����ՙ��@�O��wM\<Z�S�s�w�:v,Y�T�����[��E}�0�K� HI���s'`��%,��A,�H�6���F����+�.�&䔡yD��{o�Kڒ3��F�U���6P}FWSn��C��̜�K���-j�F��V�GS��Z<��������%�6���̴���>6�?�v&�$,��cg	�|t��ƥD\��~�����]�U�X�|T |#	�"���L���U�ǖ�J����!�Ik�/�s�!%)� ��yfgABRT��k9`V:�:�x���j���f��4
�[E% �L�G���#2bC ;C�'��M�[�����k��W�0�s�b�������>�'[r9��/���v��|a���~�W��C�U�3t��Tc��7����?C��m2A@	�xk(��i���H��c�. ��A��Y��S�䏌?��]8�����0�Ba^�����&4.�@���-��v�^7+�.�!Y:̛A$��Q�V
�ZU)<t1���9hw��[����v>Y���ktM_������
"sd���:�Q�h���F��}/LԂɓ����֐j/�k̸ܢ�����[��n9i�'�;�,\;R���}��8��!�k�b�����(۷�����پw蒒/{�iW���b���/m!�8�d�)EI!B���8Ü1m������I8mMwL�7���*3`�J�ˤw>+�M��@k�ϗ�ղ�������&��{��)�)�zğ6gé�ڰ0��OS��fs�P�iR7��9_�P�r�"Ny���"��3�l���v��]�S������t"p�yS�]��rn�yfUܤm~�\(C����0�h��Ε���=nBۅ��ƍ dd�>6�狺���T�J��jM��k�w��_�'#˩�q�j�������K1H��+Rk�|��Ry�sǔ	W�.*���c�0��r��qr5 *�A��ʢ�]��J��4���)�)F����/8�M�雗ݡ�%���v��U�������.߫���\
D��SQG��^�X�#�� �a�+R���hz:�=D�9��x6y{��9[lm�+��μ�DM�Y���M`s��W+e�;�'�D4{ñ�#��2|Ĺ�j�5��`qۣ��d�8A��$�,*����Y9v�_u���̄@W��G���� LA�f���
��k�b6xoV����@�W𑥜.+��m�I}���46��g�Y�.���=2���7�D�pd	��D���Yt�2�0����'��N�7,T}�kd?���	��G�*k���>���=ⷈ�4�AlBj���\��h�6pnq���E�i��;J��f�`!���E��\���LH�mé�3@j��ÿP^���4�w0�[J��$N�X�� w���o̠\�pY����#�D�)''�K8ٶA�E���Wզ�7p�z�����}� �>z:O��]͇:}`4/�'G�v����Ay�y�7���)Jj�P{G�y�&F����%ȂTV;'m@k�z�pB�F�"*��)��s/Ś���>���v}����H�=����)�Q�/
�U:������$�G*F�{#��ښ6�c��,�M���=c;�{gZ�W?T#iO���T�E���V�4�o) ��vAɸ�(okh0O�y�]R����d:��VQ4��V���.+#d�h&FM%a��JO|�0���
����J��HZ�}�e�3�P����4���	�����5����1_�f�T1i�\*�B�Av����>$�g�m9K�B\�B�b����=���6����v���n
D�}��Ӄ�6��� _�huP|��bcЇ���XDDZ�������r�6?l7�am_<bZ��5��QH��Ŵ<������^99	�qw�X/���m�юF�����Q�4�v���J�gi/[ت����UX����d��jB^�S�y�)X��_C$Ԥ��--���ք�#b M� ��ϛ$���x�>B;b���Eb ��|_�4�x�Y6G��Nܳe�g1d��K7����q�|�Y-�׹�����*��౫@"�6�^��ɋn��@]� �ۓ�Ʒ�u7�\;�u��	r��M3��2� >�d��d@�N����0W@((���T2�@w�@�d{��+��E_7�'����r����m ����4�ȭ;��-6����"�/Aւct}���� �QsE���\�����	-_"��և��<��2�d&#$�'V��g*o��y��νXg��?h���k��2�6/�dE�h�7
��^��t?\"�Ag�uO���W�R��1mޏx�~��&U�&�4�*�{��.��T��)카}Ul�eK�p�m��]�	��f�y̦����H�hdޕX��
�2�jkw�av;�9)i��߼>�Y�����"��5Ϥ��f�$&K,�̷�!�'K,���e��}���+a����!!�t.�ҍ��g������=��y�Ϭ�Ɖ�8��8���Hr��}#���6N��╁jZq��G���S�a]t�:/_k��﷈k�j�p�-�h����L����iFZGt<jrf�i�I`��x�T�x���V�k��Bl&ל�:t�7Q�F4Vb��K��n���pG�\OH^�UWב�C[dm�́�]<A������)2@��N>��3G�LW�7�ݛ�l�_�������>��B횎��^���C1~�nGm�e�=%�M)6���^�W��8Xڋ�z{k#�P`��(��$H���"�l�ޕqdK�yeҰ�L�tBkB����l�k:U���͒1���ve��~��0	����kH�@?��3-�UHD�λ)@�P�mۊl[�ٟ��3M�rΎ��-C�)nUX��B��hŨ�G�J�@��,j���9��'g21:�E��f��g�)�~`�wq�"�`d!h�6��p�=4��o��X�yR�%�;좄�ă�j��g�l��[\+5���(��[���p!o�m�՞��Յ����j7k{�{ȕż�	w��̕*}�rF'\-+�
Q+� �k|��0|�JP^N'��B�RT��ٹ5�J4�>p�uJ�3*qو~���t��O�ã�皥>��LM���\Qr�7���m,x/X�t�{��7M�DD��nz@�
��Gvo\#!���~�{T�ᷯ�PԈ�ɠ�V'}�1�� ���(�����0�oi� �\�����xfZ�Z7KsE�ۣ!Eo�Ju�fѶ�l��@Ϣi[��U�l�W����3�����d���J��iR �&�'y3�ˬ��9I�z�թ ��5r�GF���v �؜����ran��������fx�%�g�aEɄP���%��>�p��ſl^�\���c��%'��쌵�k7\�y�t�� \\�_e����Dpa��>�L�":�w)&U�
X�W���ژa��8:���-];�Ʌ&wd�2��h�	5+���%�A���Z:�D|;�z��V�$�c��W߭x��u�P��v�ʆ��ڣԲ;f,�o�Mؿ�w�2ۖ$}Lmt{��ld�x�c!!>���
d�� T�3fB�;g�C�(<]cF�.y��˖�w�2$z��%�,�&�uǔX�a�*j����%�~��{��F��A�O1���]v�OT5D̴=٣D���	B����Тou�i�Jp�c��N{�A��q׻�w��c�l~Ԃ��.yY�� ^�����a���V(Pd��3`���lL�)�:Y�9�2���cZ���9Qȣ�O2-Z9�����[���I���<�X�9��*͆��C)�,f�,�n9���(c	{+�H%�[����c� %�~��q}��"�=�z��I�;�����f��R=�}+�D��ѧ����U�a��
��
R��:�ϻ{�z1�ԥOZ�*R{��ؔ+U�I�un�'1�R:۩m�)7G2��a�����oQ/'"���1o��Z*Xm2t�d���I�2nߟ�1|t9�gx��W��yeQl=.�)��b�2I�FP�\�����x��23+@İ�l�w�{��:B�T�B��
a*�Dב��t/��DJ,��f�AfҌm�b`F��;����M���1慷/�k=��R�z-mT�VO�����)Sb5WW��S�����3A�i�mm6���u�i�E��4����pA���8��U 6D<����s��7�X��so]��~��	��'{�m*��(�aesy*�1Α
3
���  i�^��;(IQ/(�W{[�͕���c��$�߅��d��@�	R�ZyD�6��9̜B^����eP���c�c��Rd�1[��*D�*4��_�(Okx�[Q+o����9��I�/H�(r�D�㘍�4|}���aI9=���Ī�Km�6"�$a5@�i+8z� �,@9,��q��i/�wh�����粘T�	�6��@�P4��'�C|k�p��s;Ȥ�~8���(�����P�x{ �ɤFf�q��W!@&inOWH�����Gl���X<��^�%�+����~�W.��
?A9��d8Y��vZ߹�8�}LB*��^�,"���2�o�A=(z���ry�+�~�y���������Dc��*����=�PK����]d�O��h�8����LH�t,�G����Wm��.���vT��=ɮR5@��T%�r�;���%�#o蝒Y� ��'\�r��y�n8�|{�<��N!�\%t&��;���8n#���m"��6����+É	�N���*�A��7Y��RC����Ū[/rT8�f_��Z=!Q���) ��хm;�e�>~��0�����C�R�c�H�*pG�/��_�;h��58m��V��,i0�H{�����c��{��i�-3ʨ-��HG�1��~F��1):h��������IJ)�	 �5SfN�m�y�}����D�"�6Ǖטּ��g��> �Lp�q���^��JuҤ�85/�f�[��{!�{q�HjL5"c�uA����jş�+~�IGx��TV�g�j��='�?A�f���^��?�}�i�>�3s��a����{�IT2�
=�Q{�]2��E�~b4ޱ�_�'��^w�p���� E����F���þ�Ta*�F��e��Xn��t)��OF$�lF�� �w1��{M�Sr� ;��Y/R�o�бx=�@AW,l�MZ/4Bwh5�����Mm�3v�HՎg�	1l2��*�i�d®Ч�*vpW��H��DK)�G�ơ�c�,�-�V��,Ҩ�P�?�=mo��t�8���\�Pdvo���*�ϒ�T��#2�2?7.\m�_�ӮC���T|���8�@c�8dU���T�()��W2Wxd	>uR((l-�B3�8^y�Wt	�l�:f�\N��i�N�>D�z�w�أ`���]�!a�c��226R6@�F��t�
ʕ�2v��Bf�
˙K�D��CZ��WQ���r���R�ݑ�B|xB" � oD;���0�vS�h�0.�r�պn�8�q ����g���1��I� $�~cC4\f�P��m�LwIv� ����Q+֒hh��M���57�W�_wpz�^�����h�>��S�1�L��|�X� C2+����� ��|�ta1yf>V�}�{}:����5N���#��)J+�-��\5�'|�b�c�:I�B�N��K�B	�����U��0�	��%E���A�Ref�Jd�ծ���r�ߥ�IF`U����]&Ě�f��S�gH�e���`?�]�u�u��G*�Y��T�u0�b8��e��K8��!\��{.�*��k��{��!����wN;�N��+�:�|�Қ���<1$���G�p����6t�w�����h���8$�ت%ɮ�Hw%k�����X��&���A��yœR�΍���m3�yz,Y� �|=+"ϰ�d �5�K%�R0���IYd�pA�(N}���]� ���H�Ε6�L�8�/�]�\������^+7Z��߯��9l���[Hx�e���+3uF��Or�0Oa��T�,��jgv<p�^/�Α�&����-�]��6;g���ew�01�o~��,\W��g�2�g�,=us��)h7K�{͸��S#��4���jAw�7�H�m	Y�lkW���:<�]+6�l�sƋ�����Q1�oF��.�n�:1&êBH�ߖ��`@y�Qg��cٸ��I�UU����LΚ4���-�Q�[���_�4׶Li#�~���Q��wq���8a��/��i��Y4O�Cf�A�`@)E����B9�r������� ���}|ܸ�S��il�pN2�,Bq�ue	#�P;P�M��u]�Ut[T�=�q��E��êŌ�SS�`��Ak�KF����SX#�u�6u���,W����>�J�
��Wŗ��/�7��\xv�@iw>�j�f*F�����;؉J�5��`�0&d�Ⱥ=h�灩�i@+0��ʈ�ag �χ�oV��s��&���Ĺ�9����S���KW���g�:��WM�5U��fv?\��#�{J�j�`��*(a,O�T��v�Xs�q�6O��$1}]q��M^��5I�"�>�s�����%3�Y�0ۥ�1��'���A�B�
�H2b��p_�q�a�ᩡ���r*A�f�k�7;ř`�O�O|���Ϋ��,�w�a�|�O7�z�,y�D�)�����m5~0��?FTŝ#Y�Bu_x
�p(!��s��,Q��x�r<��Ыҡ����T^	�CĞ�b���CG���d�v���� ���HDN�1T�6�L�G ���N���`n�
_�g�ˎG���r������a�A��J�VҮ��������"jD��(��)G��L�b���4�Ϙ�
ڏ؝h�B���$-�f�t��LV6�*�xX�X�d�YC���g�����oᩡ����A�h:�$�Aب�C�~U:c�!�~�uyF��jc�۴�^Sxk:��e�A�#b��K��p�w��c���CEV�	��A�+�L��U<@�u��6���L��ſ�}��;���� �Ж$��+׋Y��H����Ik}g|ۼrX�T����W�Z2v��/�!v�B^�7c\}�t�zԵc{=�\�+'|j�X[6x�|���0[��H�Ѓ2�7�iLQ�����]վhA���ⷍD�*A�����2����$)V,$*�ͻ���=�ҍ���?����s�ǽ6�{,G���a�q��>��}�/��P1��1�
y)���#{=�:�?h.QP�
�~�M���e3��ѐ���<��������*�c@P�6<{</�BZ��"��c����G��C��d�ZQbߌ8�+��"�$��t50
����Hi�OK�è�"��c+��JL]�0��d��.�|��l����,�Q#+��ۘE'&~����?0��eG������о]8IzE���K�83d��K�S���x�؁��{>9��f�v��&@z�B^�40H�����x��U�V��� [��)�ǀ���5���B&�9�Ww���.�u��P����}JL�V���!FfB��\3���QR��/K�g[V�:	���V�CPL�~2�G���<u6���b��a����T#35_�n�]��4j��0	,����K���*3۸��Bv�]9{swᓒ���{��_X�J���Qz@���j������SkS�;[����V�%�Zh��Jy�֑̎T�D6J�բ<��–��~��&�t�2V��R*���4�Z�ـ�Tō� f/���q�n?���V?�
�Ex��u���������vA�sm/i#�y%)pjc&FZ»�O�y��xq���?Aٌ�A}A�:͙Ӭ׏e��68��$����Q��y�q��̏��#��Z��`u�b�NI��B�N��k�#/�&Y/������unū���[��&�L��dp�M�-��SZ����@�����'.$��b\^Z�ج\�s�݉�W�h��}D��.J���G�A�ڀ�k���R���솶�qX���M�3iI�e�� ��F5�.���V&&+�gƣ.�|�d7��S+��$�f6��4P�$)z����Y�H�%'_�W�E��v��"J��B��bd) Ea��hq��T��V��\�3��M�2G�̃w��V���+Α&����{C&	��x!���!�[a�	kg}wx�ؾ��a�Y��pYA5k���ۿ���.�3���5O�[��v�6wr,4>��Nw#�Bf��1�%��Čg����,p�>�+��}�E<�ZU���^mI�1}8 ��o�5�Ep��W���<��"����c�o��,�K&)SOi��܋qƵND�=���N2O�Q��('�gX؂!C��� �����P�y����m��<$Eg�`��^�Z�.�Q�s����_�(e�5���Κ�u��<���z&:�׍BViV�'�ԝ�����	���,�s�zF������~ʲ��Fƽ-��rߔ&&z�����w��py��vū�n�ㅕ�!�� �B��r�� ?�U,�]fPW��1ve����es������y1�$Ab�9�*I�|�g�'H�f�ĬRct�š-�y��τ�7X�,_��ʋ�m�=pݗ:ͨ�.;��O�{2�h�O��3/����o��<$�z�#�t�y5rAr�t}{6Z{&��
��*�DZ��l��߄��R�l�9��)��=Ԇ�L��L?�ϊ��Z�}�z�:W$9ϑ���!#)�A�#	wyh�}L�#�|8���nM1��N�����)9�.'~��֠���Z~#<�5e1	���` ��P�6��|v���5���uO4`d�\3��_��x��p����=kej��E�q�$G�lM�>�q!y3���$|���=W>��U6���[�(���\-�k�@���4�֛�oX�D�d�d�\3$�.���etTu�q���־��Cp�GT~�r�&vN+����Y���\��l��!�h�5a���S`[�%�������؈d�)I��|�玣�㛵��vg�͡���m#T��&�T�7iFYK�8I�W|"�z۽��eD��]�?
P��=��t��u�Th�~$Qo�'�6r�=t�5]��9�P}X�] +0�b������2r<��n�h���A�i�6��H�H�'�;%�@�����bS�Unk����_��9]�}��L�V�ډ�;�ڀaOM��n��P�/:Q��gF���w��B�`s��k� _Uju�eh �݌cxF�MC�oӮ�Qjv�%Wd5�����w�����ܝBW4�ْ���h8���|�(��փ�����7�A�es� :-S��)>h�_��ҥ�?b����!:�lP>��ʰi��A�d.����94g��2���=D�|�GC�����p�ND^FD���(��N�~����s�!�
F���V�s�<q����"�������܂ɭB����c9�^�Z���Lp�jNy��tO����#0�Po��%u����]mN?3^�wz�ʸd�H
[;v�q�[�u�+�E��0G$�����H�����$�n���:��d"�H1�Q�+�3�/�h�Q9��nN�����G��U$`��Kq�AU;�X?���2M����6�Y�����K>��γ�ͶyN���z��&�����;3.���t��y`7�bm�=�C�rRf&��vz-_�E A�/�6���-M��t�ғm�|�UJwFF����/����5�$�s
�j�������3yG��O���K���cR^��O6	��Y�Q�*f�n ����F({��bU.��@lncV@5bQ;���]\Y%0��m���Y�I���8[�)�z-2h��BBd�OMcz�-�mJ o���{@�5�+S�u:�+�і��/L�G����L�o�= �GY2?-�VW����^˼V��`g�bG�FZ�)���`ӫ���_�Xwt�U�g$L����7���R�k��V�5�thz	u���=`���8��6P'���p��$P��$?B��t�`x��`����7�n�E�g��A�X�6͙�$L�K�j�c�=�N��v44�8U8ס�r��	�H��F���(D���!H�;�Ƨ��փ�������J��}(�~j�%^�I0&kU���EB������C���V���:�,$��+4�T��4�%G��Wdb3܈^�=�]]�б�
 �г�Sd�'޷�R�@�y�!��=�'�^�{��a�Ĵ�.�h��_~�A�;�t�}���Ǜ�/0�קj��x�rj�Jo�;	�6b�C��t��9=�������w��k;�����/Ob��������}���R�2`���y䇛�He[R�ѹ�S&�/�,6o�Q���f�_�l!+r�Y�\���>�����x������!��S����M���5�'E���ŗwm�S>��bԘ��}�*� @�?�-Կ1�o@��\[.޿%26�\B�c:�os�;�H��Yl�u;>�R�|�Q��X�� .bAY�!\6Y�6)�q��TIw�k��.\*���洞���ŘB��P"��/rU���(o��E�a��m�����m�t���
$Nk�cT��\�ݧ=i��;><5����0Uq��E)���a�7���Η��rEܮ}�	���$�c?����kX�K#>�q\P��l�V0�zh�l)K�K�h�ku�"k3>��v,����yQ!�eZ`m��|�E����=�����i�w^*�%A}g)��}~d��+�_$O�t9�+�����G���-Cp僝�h����� �m������5����g�l�G�Kn�#�0���y��-�L;m�F�6�%dd6�wp�#g����V�`A���D���_���geC�*��x�L�P�c���f�y�ڗ�)��%,Zo��x��BݑNG ���oB�Ş�MU �ə5�:�>ꐯ��x������^��A�-���u)<���S�UFd���1$:m�!��V�#��`��>P;w�:�D�����Ϊ{���]塁;�J�y��q޷����p�2�}�f	WN�x��(a�����}5��^Їx�^��-�Ѓ�����`�I��Gm����n��X2E:�Y�Z��`/"URd�"#0I�dq��/~׫+�B<��-�����k;���|��js3Ӑ��y7�Q�?���Ĕ�q�f�܃�#}���JM:�T���D�3��*��|�@�+�O�SF���!Ȥ2(��&��w� �M��t^}'L��o�7'���K-?��ö�W�kX1w+�Hw?��2���J�:�NA"��09C����C��,aODs�!���w+�6p�H���~�֜��N��HUu�*A����E5-%N�톚��eQ�v������h���]1U� �i�G��ad��BT�g�� �L@Π��u$�CF�%bDKVxF�z�{j�H�s����̓ߓ���Lȉ�)1\м�62�'$�+"�'O��5h%��X9���В䥶MҼ�{����m����`)7����^�V�Td�Q�`<����<�8�^�+��q�?^wS�Z���|/!��A��<��N�8����@U��7C+�E�L�I�F�"98�&\o�[���ҽR��/ieTX"�\$��$�1>��ǄXC\�զ�(x� H��Y�"���v��RRy���6�} �.,��?)�@(��e�8�~�kù�`��l)(�@.�L�0��@x��-m��-�=�5Љ���H����O\��3pV,��xg�y���0����4{���Ѻ���3@�\�(ک12i�u�X(&�4qgWA�%��Ȑ�=2��U�.H� 0!h|jQ�D��U�����*.�w�s�H'��U