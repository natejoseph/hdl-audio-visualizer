��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��E����C�5�_8�'y��>�1D� }"�^A`h5�d�fWG�R����T�l��2���0�oI8���j�{{�4KL�R����H�πY{�hh�(�lQρ�mˤ���_u1���[�~W�N�Zn�Q�Q�7~�u͈�������F�n�Y9�?���Tץ|��ӈt!ZfX��m���Yo���+D�"#�ܔy	�Ko/j^.��		�#m��]�˺�}K�L8s�<-�I-�(��*�|��vȘ�0��y��j��[%1�)�wu�mi���$�O�e�GM�,q
�w��|� ��"�:\c'��|zB��P�h�3�V
�.�b�*~MV�Lբ'R%�,����9D���X1x�1�RL�g��,����<[���2,�'���.Fr؏#�	%��}	�Ӱ0��١֮�Q�Ԑ�ej�i�K;
8ן|������u���<����̄���f��G�0�Tr&�6C�i���c�:�-�sݓT��ۃ���H)�J���|9�yz�_�M�o�Ѝ��M�'U�A��(6=P7�5?HثX�9bϮ���H;�uTa�` ջ�0��U��M �����?0�o��Fm�����zv�g&K��5�9bu	޽p����!�h�y�xJe^EVȃW'�<x�lf.r����i$m,m�ʚv�r��q0�Ebs$�϶W<�\,kX��)�J��eC&8iE�uT�~ue�����ɾbR�.6���l�|�(-�Py���ٙa��F��n1�3���D��̇j5/� UqR�9�X��{��q����Y
�%N�_y.d���n��y�h&������8��ど����1խ�D!I��=n���/z���R� ��W�n\�ږUg��,�baâJ�����$,מI�t���&�;M��s��4l��]���"��!��sל+����%+V���Q�y��hb'�����}nO������+_����D!=�on�};r��Y|"ʞ7x�v�c]H��L�7^c���W'�]x�=�D^����������'s�|smȀU�ɖM��E���) Pf����j�;k5��<��fD��ʠ4����*f��7z}��۪��.w�}��P=#��o�rʱ�M"�� ?"�Q��sƭ<��fT���u?p�a���O@_�p_4�h꘨�8K�2�PcOP�Xr; �B6/G���W���m����Сe��`�7�r����٘҆r.B<dЃ�I�ea����4�&��"/y'Ґ���T��1����U��g��������d6�0���+���������(~���
+�S�g��|��kJ�cE��*Uu�ɻ��~�ݛ�Tzv��]&A����e�J�AV1/~��Cӥ��Bn&����BE������^m����iD@	{��.�x�#����ġ��t�vV�V�^�W"��F	�J�l��a���~�6�I/�r����z9ȓF�}.T���ԐK�ۡ^��
V�S{��o��!ш��^��@�]{��&�8h�+�<!k��iZF���
f�>�"�u�6�)�+�I��a�a�N���ܛ�I��2:�G[lV��-�Ԭ�uρM(̫�Χ����8�2��j7���h�%2ƙäɩ+��1���g�b��|}���|�qϴg���1�ZrG%�JJ��3��Ȼ�P�6�˓�Bi�&�$�S�&'��.Ovo��l�������3���ˣV���M:L@Iw���^���W�C�;0�v)u�!���9�"�n��A��z,�,�8FYw�6�쩅��t'-.yF��OpOh�|)�IYy�,������YV�_"zx]"�D���V.0z��o�*��:�Oū�CoH��T��B�!����
(�����CTE������&�W�����o�k
�k�6���Si��M�Ѥ��9�(١۝�1�Q��k �\��G�A4P�x�Ŗ�>>�ԕ�pf`	��������>w�ٛ�g>��]�;���Dz�G䞵A�*�.�9W��w�dO3�ۇ�ێ� w!�]�Q˻X(+���Fn
�����y�Z�Z˕%{�W�^Q �/��I��Q�AA+�|�46��!#��;T�c��h/y����1��+����H�.k|~	��P�u���kVm��*�۸�j�$�)BֶS�4��,î��{�ο�]�L铤v7�K�6���s���w{m�η�e4��_��r8A
�Mx��#�U���Ճ���N��%��Tc���W/��	?5�*1]�ٔ���9���Ap�{vӆi}����i�5k*�甯
�>be��^/�xj��o�GK�%?�/�(�>]�~���T���S��hH-Ԍ�"l,�2��K��;��@�A�����EF��'EZ�RssT�|7WǤ�K�S�K��J�mű�����e�����C4Ͼ��v#C�P�#4�P;*��$��p�4$�<��j��<j��pԳC��*�9s�[/k�U�����"��{,2^5;��N%e:p���
f�/&e�^+m�,f0[��=�&�m}�C�H���9�<�������+�XCL��,m4G�8�9�z|�u8u�X���]yb���K�?@ )*�Q�~+�-Ss��.��?�w/݌�+��ߣ"�E!!){72	��J�:�~��8���mn�ΞZ�z��S���((��R�=��o&""��\����sp���r��jP���y��2<������<���4}m���厸sCt���H��yZ�I���t�!��Z	��#����a��xX2�@I��,�d���+>�J��^��	5>� 1�7�q9�I���,W����7FL�2��E��'׊%}ܩ�U��	�1���R�Lx�eIR�F���%ˏ�9C����	U9��#3rI�:�rǕ�#4�I�RXc����e$ ���YS�(�}Ĳ�Zo�b�Z��JC���(t��	����F�����`��/���C�Pޕ�u�Hq����Or��b��e�>8�;���Mu�<E�kQ�J�ɶı�Uؐ4�J��Sf.���c�s�.�͑mP��{��+
���OSV+��}^<����C�����q,����M�q�Z���U��8{�D�E"��s� l]�T��v��&"��(��_M�SZ�`��B F�5��k˜CKp]g#囃�o�#�����iPC����{GK�#��kUC�${��5��K������"VVΉ"�&��k�C���-_��������W �_
�q���ڻ%�(ާ��vs�!�g�+�S�CΉ�w�ꈃ�oTO�����`��-����)�G{G���W�A<�U�d�v�_��o	��c�V�nQ�!�p���'f�������-�&��	���k����t�ޝ�c�dYZ�AX;p��\����V��{?�܂�st�T�j�&t`�k����u�d�K�w����,�L�.��y���k�����G�~�i�����^=g�A{�-q���L+!��=���CRZ��E��L��rͰxYc�+^<�#�_�j�\֬6�N�-&t8B�d�(�a�G-���+�����၂��� K��O	�xI_G@�D6���a�kBx�I��9������l����f�����hR�ۭva�~���XZߤ��2n����e���#�N�.ꪀ�^�.���X�r�w+�/�n@'F�`�����\OT�8$�s,�����\ה�o�dh��̏��Hv�w��Ԯlk��bu���J;dEv���w���~����`B�,�(�i��xF>�i$8��a��T������"�\�v����=��V�F���4���H`��ְ�{ǡt���Cã��O����/>p�ζ\���.��H �ݗ��~n��*�'t��ۂ��_�ֵU�R"��ir�	}���$�4���&F�ws��s�U�J ������D'^}�q[���-�ᯃC1]�U�غL��"墍g�DW�_��e�n�Cd�ctz�ײ����6�:x�Q߾=���lkc&��r�%M������*>�z����0�WIO5��!�.���i+=0���X��p�ҝ-�S�U�y�c9�N�ڿhՏ�
3NÐ�ծ���J�����C$�^��h_����MCxP�eϚ6��N���;2L�G�?��!<_�pI�/2s[��M�u�L+JO��hX�!#|�F��������/��)��>�����"��ZU�Pp�D��nlY��^�X���u��T���\�x76O$R�ՑeZa�2"}\�.#�����<���q���&*|X:��a���c�~�s;3N���c�d�����P����~�����;��d�<A���0��a�[&bt��z��NV���MJ�μ�D�-�<[WRu���&�(��N����sb�Cۓo�Σ47*��&��iΙ,�3�r��<{E��h6��|��D@�R��c���������e��F�Ӈ$�ؒ8�������Mi��z�4�d|�$ζhLH�l�Z��A��Ϛ�g�4l�n9�&�M���ho�չ�:3@�(��S
�*{Պ�75zcX��(d���3�^:��H��xN�n�m��eG�����b������q_�7.=uL���p��63i`�lV��&���� /�w�$��[}�V��Z�������tG�5�@Ř_ѥ��G��d��ԈP��$c�=OF�R�m�~D$���*,�_M�e��J��BH��F���q�u;�������w
�����$��CZ��<?�\������t��S��	6��3����Tx���̾m����V݄��T�{H���xLPn�?�~D)�X!��x���i:p}�3+��&�|�yj�G�=f���m�/˹�oߨ�]�dW!���P'b��P9�7�=�e>.?nh���~��14c�ک�������䊗#L�S�`/d�x	���J��n���'$���2�EviQ���I�H�ZӸ�x��r���т1��
���n��ԃ6��C��L��ä�c�t��J���GPզ�7�B e��#f�fu�O	i�:ʪ���ρ�\�modۜA�PA9f��&yw�%OLZ)�y���ׂ��H�g�bάk#�Uuw��V�LrE�'1��Ę"mQ�U0?>���O��\E������j���5� �h���5A[��RG�{˼h����Upo��>�G�Kz�c-��R�O{CÊ/�|!hZL
�໡�|a��KONA�nz�[b����WB��!,XYt�4̣��JU��Cy��4�����i�
r��!�D2��n�{Di�c_$L핔�[���0Nt� n��~!��_0NS� ����޷�F��FQ���t��Y�!�T���,�"����'�]O#���Р�/��鰛5^�+
�bC�ڣw�?�Zc�9��@هD��բ(�8)BpJ�%A���%]�q�:tvp�j��9<���b{ JY�6o�~l�1eN	��ݐ"q}���������q۬¤:� ��/�m$;D�˦����Xz�$�qz �&�/�L/B��D�m��o���3t�_���P�=��ف.�[�6�	�.]7���2^C��'{�JMK�n�V�7\z��j�U�����
��A+1&�B�x ������5�./2F�~����s���_�%�D�V���˟tp�2�/��LG�RaoBi�(^�~���O��rྡྷ6�NXTP�+�
�{�crlQ�<M&�С�0�B��t?�P3�r�K���"#�iJJ����C�e���I�����G�zO��I0�a��U�?�~!q1�M���#-ِ�&H�F�(�(�IWȕ��)���^�.�`Z�������L�\�@}#<t�zn¢`���5�UzB7��ȕҊ#-i���f5u#�h����� K�TM^����L@ef�Z�d�6�˨iǇB^�����-�S�2߸翏��7Z!j��׌IWW�u�$�J�A��Ο�w~
�-��U�4ϟ�q�p��k��3�v}#ya�_�E��8��i�K��+��e'���0)���sz��E3W������=5	J���sܨtX�����K�-ʺ��X���[{��~��@4E%]HYs�h����I�f1�VŌG�Ờ�}`p�c��2[�Q�T���ꓰ�@PT�6�r�$\�c���]�	��;��JX>n��/Dw��>������J��V�?�mɠ��*��D�Ｄb�&���8��=zgJ%��^�~W�"��C��m2q��w|�[BԦs$�b��
��m�|���'�¤G7�ЙX��ǒ��%�ɺ�r9�e�x�^e��N�_��Hl)Z|�a�I��Q��V�r��xQ �����m4S4�'F��EW�O��"_�M0Pmɣ���#Dk��{�*3?�;���m5\ӥ�rI��������fM�߼k�BF��3:��i��(=�e���5?���l��{v�@��0ld���|b�CD�����5�T`(�(��k5��_ͽ��9���߱�d�Z��!�^�N�\��Y49�I�K�H�|���E�)��7{^i�#v5Y�H:[<S�#I�,�!�m��Z�Z�-�4B2(�tat�|�g3�;�76B�/�4��+�0��EC��t�X0΃�CU~h:�}����K|-�2 
��}@�T���K�_�Ɋ�H�����8�Y�UP\m�1/����c�}�a�l1$MGxݍ5��	�x �.hI���c��쏚�U��y�]A���:�wN�rP��.;�VƢ�ִd-�]O�Sq2��]���'w�|Ţ2</�hv�Evs�2ݫ�Bك*��m� ��ј�H�5_TD��=����b�]�����|�)^�M?���{-��~ם�tKW9-H&��:voٙҌ�>v�I��,��Mố�����#��ũ`�����8�O���C��F�Y��e�Ra��b��r��B��D.��뫬���=�Ξ��2!L�vf�VrZ��F1�J �[=A_���8�m}")�R�$ڎuW�� /���yU���m�䝆[�L^<�L��퉎�nU.��Aj�j@R�y�пi?�1��7)v�H��ϑ!U[8bUe��� ��
�B�Ƹ��O��7�H7�i��V���	!�+�A��v^Viom�}��g�o� �p��#��D�ꗺj�Q�O7��*�K�Bw��
?;���wɴ�������*�Y76Z�>V��3�;�GQ�"Y��T����x�����Qa׼ ��&�(�`م����4�9o�Z�EZgC2V���QV|���X1��*]F������~�������ܖ��,�q�,su�ẗ̰ɸ�ܺF6�|�^c�	K ���6�%��y$�啓��D��p9ӯ�B �Ն ��g�%�̸�*�ݡ��#\�c?r�A�T]��P�8�ˊ�T&@�$�ww��>ۢ�[>/�"��YFkl���E��]e\ޔ��B2�9O�j��B"^'���Z+���I���HXW�Tvhegj���Z�;��k5��{�Ēj/�{%a�g?�ADd�2O��{?����S�B�ݓ,��E���|�9\�����@�/�|7�(_��c�\L�y%^�d�2��a�����[�Vf�M��9�+��B?\�Z?�:��6�
"�r�Py�����FL�H�8
7�>�.dP��Ś���8`�4Hޛ�ռ��h��|��ɗ�-JuiW�(x4%_2��ͩ��B~���J_����J��CHʓ����B)[�kH�mS
�B�P[\���!�Ő���$�/w������Gw�h�6F٠t0}�v0T�8��%?R��I��p��}懀�6�a�6���K��5p�fV~�wY�߶��q��5(��4+Q$�o�)��A�QMn�
�4w�ӱ3n�Is�W��#�a3�ԄJ]�-�#3���|.R4ĪͱY#ꌖ�")]'�-(-�:��Z�i� ������:������/�e딃��*;f��s�QŶq_9�%%ؽ��sX��E�H�#�!�{�sb���Z�c@�T�j��{Aq^a��|�\B�Q��/���b
����ǯ}6K�H�ѭw���^	�p��
�:-Ut�|~��I��t4rHW󻴌�s�Ab���F�2`��>�E�N�U�߿aޑ8�qrDy�9 ����ؠ�����LY�jYFL@��������os���ƍ���dV�=�&��m%2x�	��J�XP��)�"�>��~�z�*ڸ*	V�|(Ö�T a7qj �js�� ]B�\]o�bsM�i�U�uː �$&N�OO�1�=�>!��&�~������#Ch��UL��5��e�\j�S�t�5$�G��a��z>�A�3XQ/n#ڟr�GY����+��C��\δ�ML�� ^� �\[qe�%�V��ih�@_��:B�KE?ʇ@�sC�&���B<juov0��'��H�z��H�hK�n�@'��%�[��KݫUhg �&x
�+*Rb��>����c�n�|�|�h�%�f��ۛqN(y/�������G��A#�ђ�4D7ur�3]���z���2 Z���*��ͽ���"Hͫ!�͂;Q�E񏊃�gA�²��&U��?#�	�����F"9�/|�Ѐw�m`'���뻱jG;��7Mmm�{�u�v%��"�H% %�����M-���D�w��A������(�oK]`l4���� iC���D8__G��=�~������Xc��E{>�*la������mz�u���Z����.3��j���o������H����M�t:C��|�P	��~��c���t�|�<������i�9�>��XiF&,&��E����c�PG�)�
ϩ�����l������Ji"�4�������zE|ڹu�*1+��ΗuPY=���w�dX�]궅Ţ�#v5�*4��/�O�I�>���y�nj뻘)�&٨�v� J;��"`HԾ�R��1O�(���1�C��J;}�O,��:#J��e��WP�CF�}$����z�س��o��c�9�{�����=I���I�<��2��i��)��=��a���Oݨp&���/�yXe��SX�qV���� )��o�3���7���k��l���N�w������b��bE�H&�M����S��dn�(g�vȍ��RD�&���������-��2����g�#�4�6$[�dߒ��y�$Eީ��$c9c���=�2D�7��[3+�_^���5���J�H�������=@��	v���csr���?��zq+fxz�����Ҩ���i/�0����3vŢ��
���54>Ѳ<����:2�ɬA[T@k��d��T3+��4��־���}�fg���n�'��_.�O.�C�קz]ҭ# ��|�[�j?��'*�x��+�F_`���IH�Z�g�V�J�Vk��e��]�~����Q?��� ]/�j��p}-l/���b������G�b�w����gY�"�rc'T�p��%���>$6�84F�D8�7�¼#i�K6|rc}"��;S��R�����x���K�c��C�^���&z�C;+ �}��9#|����'���4IZdst.Yr*$D�\Cb+7��������1�k�o�dF0�w��C��f8�l���@�S!���<���}�U�����k��Y�����){'��179/z�&�¼<F��vK�d�zZ�DI:+a�_��Fdz+��Υ�m��C ��k�iE��?���4��F_LJ��8�t���'��,!ة��(�$܈�!���g�@���������(�y�S&��톖���"��z9J�Vz�kGG�/�N�P�i��tG�W�㚱�5�V�Qˮ�p�t���c�=>���d+�(�m�q��WFy8<�����E�;��:0(���>Q���Z<V����m������jW��+]�2���#�`]V�uߓ�\��٥8�pP7aw��B���H����)��iK��X��%�����}�H��S�FW�1�R)�$Q����K�ֽ��Nv�
����A��6F�jjZgC,�̓�=�r Z����
��ͫ2~�R��z����p��c8�R�DZ����oO[%�j�� �M:�xB�M!8I�C�Se��D�I�.9��X`$�Aw���}?��8��� \�D]L/�7��eg/S��m���x�ѯç����g�Xˉ��'��r����adP�dumk;��� �K�n��9:�����*�
��D�x��N��)��x%�_��i戅�>��Y��nH;���I���D3YA7@���l�E�^i���ð�2�����a]�Ŷp�$*Gc7����%���{�=Pq���{���2��#=����b�5��v^�YPЊ9Զ�I| �i}\�)�NF0I��zLM}�I�P�}T��qBK;|�9t�ɸK�-��Q6����ӹ�X��X:-�� l�R��6�V����5��� c����H��bN�t��f�٠�;b�t��q){��&���\�<Ƭ�]��c�8�O�P�o*�!��
|�?��������R�t�����<����p��fa��ZK����I�<�������ҺZ�tq
	:'���}���%q}��	�'�}f��x�P$�p�/5��#��S��S�jf(9��e���k �8�|����?�[�@f�s^ȫ����Tq>'0�������p��Q�K[��]��I��s��H=&����"�2P�.z�����<�D�{i�GiT�e]ߔ���xI�'y����ڠ��ngq��'$ʍ�b@��
fyw��29VbUL7��oS�{,L?�7F)�1g�$Ů�5єR��3~����Llʨs]���ZK�a���k�=��۬���k"�$��H�R�k��ܞc(����Aoo�[��-U�	g@7zW������5��]͋�����v�Xg8�x���.�84������E��5ZD���cdV���;��6R ���4X�r���9��
�s~艕�� ,r]Q�Od�ѕR[[>}=K@���=�������.w����y�s��&�Ʋ�9Æ#���ф#���ދ�����UH�)�gO�3'�~O7���V�U������PH�D�sc��@6k��L�h�B �
���
�G}�o��j�Ӎ�_u&�D�N�2n�F�E�$��1���!I������KҔy�CQ��U�k�m�|�	Oc���A-��oy#��d^	ofb@L�&����֮�}Ev�M�i�X211�f��U�I�SIJ�g�8��ay����='�XnZ� R�)�!�Rz�ԑ�A��!��Dzɢ�b[�l�`��H<���{N/P><���S��l ��o5�Lf\�p���k���B��*@bY��9+QoH�����1�����I��mj���/���އ���6{>�ޝ4t��_��lԛ9]m���`���V�g�
i_�e�[�#�uo���K��\X��K��$Pj�r�\l��*dX!�f�	}2��5�w�-����1��+�l(��q��5�拧n�^�fG�L%DS���Rq�t�Q�IlSW ����[��Ek�?�Ub�2�?bcLC����ŮS/8?$��C���+&5[��: _�У��#\<� &�*_W�ǆ]8�/o�6�&T���^Ӛ����c_���H�q[�WY��4��.1�?���&o�:���4�&|�?��w&:T0�c9S�QN��~�9��#>K�G�'���*;�4��q�fX�b��I��i��5�X�0׳8�9 ��%P�n��of�Z|1�t-�Ō��$�����U1��ǘ�듯HTŀ�P�Y&\��=���L�y��(�O֞�U��b�f�k�/�YX�_D,'���טALv����D	��a�4���m1�h�ٻAI�:���
���H:��뀗[`������2t�7y|q�ۊ�Z���4b�lD*˧����?,�^7v����JS{Z�ls���X�u��1}
��<�����%��g6�V��5��8"��+���}ek�̹�j ��A�i�Z�m%RT��`	*hcQ/xy����״j4����
��v֘LQ��{Vh2����H��H��J����;\{0q�^�(��J���X�!yN�������J@ԏ���<��sZ}T �ʀ��B�'?��gAiK��9�Kao��6[Tjx��'�P����Aõv�;K��?��z�9�Ǥ^�����l�����(����ʍ5S!l�����B�Ԃ²B;�MŴ��$�&�B ��ᵫ��}׫J�8��OLo��|֑�-8��m�t�m������׬��]�x�#���
}-��x�YU|�B
��T��.{�E:���t��\�,sz=��Y�y� �A{)�;�P\!�~\���)%�[���	?TFP�7!� ���u]�v��=����|�6�zGE�^92���X��,�!%���,�ۭgi��9�HOS9�[�~��%���Z��`aqw��>P�Sܪ�:��c�H̐�Լ�'[j��k��]Cz��oQ3�ҵ���I�W	���CN	F,�hW�ȼ��DΕz>JA_�����}86}�V�Ws�N�YYgl�=�[l`�ƻ�������x�mkP��&�V�͌L��\�a~3c��6X��i:J�s��n���٩��ļ�T.ϻd�Տq���ecR��Q=ro[_�+��ֲ03�2m�Z^{U/�'�s}��ގ�~^!�m%F��]���#@��`�=�FQ��r?o_񨪆�y�����X"򖁞�^f_E�d�裓��9�*{:Gػ1yc��4��p��/�8���J]a�Τ�%"<�!Ųӷ�.��]�w���T7mG���J� ­�h@h�J��Ʉw��wO�~-��owl��;�W"���D��������ʮmx��@:Ӟ��~V|{���[�*�Ɇ���->�»��Q��^\,^�4.��9,�c4�ܭ�MKd�^��1�$�BAm��	�ӆv*�����P�r���|&���R�+��	�=u���D[��m *Gݧ/_��P�L�B�A�7ث����Qb�cռ��B���m���$����e�����m��^�=��g�Z�L�|���=<=��C�ОG�wӼ���v����r#�ؒ�a��I4�Ed��Q���K߻� ���ݮS�Fԩ�B��P⭅ȽnZV��y�����71j��]}���F�'N��I�f�}�wV3Qj�z�%��^1�7�{�7�|h��Spc���κ����
�D�C�ѵ�<]��h����"`�8{Xm�R�t�Z�,m˶�Ō
B���G�-k1�<u;��X�{q�:\p�ƀb�{�Dr���z7-�
!W ^��
0b]nu� �=w�ɱ9����sl[��Ͳ��k�3��	���?�7�$�?O�??�d����L\��������c�1��(���y��C����M9� ��P�g�6�\s��f��=*,6-�bZ	J<�-��i��뛝�J-��7�}c%}O�`����<,h�4xz����m ;]?_�w�!+��t�JVEdK�OR"ވ�6w�]�,�Y��#>X)i��a��6G�D<�R�(���̰]����0��J��|�p���$�0 ���Q�=�*{ "}\d0���0�%���W��0H��Ý%� \p=x2�( ����l�T�.u���M�@S�B��T�-�OTl�\�ѣ��RJ���8DN����n`7h#�t�cꆵ����ӣ�;���b�/a!��������r϶I��H�ϳǳR���{W�1[�I��������5�HK���w��N�-�M��̐Ӏ�����Мc�]#J\���Tm��P�,론n��c:0����z���B���	�;?�-2�X'�������п����y-�	Ƈ_����/�市��<1��h0gV0BT���!�=���� ���%l��k�����A�8	�?�Q��f4Ӌ��K �p���d `TB����܊��궸��k���6Kl�Ddg�l�V��+G�Q��)��AqD`�1�BD��� V�<�?D�	���;�M���/$�.Ĳ�&���?vB�D��|=gT`����=�{%�3.[��>L�[�@�I7�g��u娤�)���
(\��C��m�2T	�i���U��8�z�X3��O������|�9�"}��OJ�뺨T+��稯%�'^��Z�z�$���a 1��P�`H��3����cfWP���!��d���/=�3����_��U����ɾDU:J����@�LM5V�e��n�3����^_(��iz�]Էap�=2@�e�Ur���#��?�=N��5��q����.Ѣ�~=�Yu�F�R�Ȟ��(�5�HI�"����/�[LÒo��Z*�D$C�H�}��f��)*�؀��Gmtf1Ǿ��;�.�Z�־S�ͻ��C}<��(�ДӾF=C^���X�ޭ>���)#��W�4�7ɥ"F�#�8
S������\��2��	�73���4Ȩ�w���9MH��(|�!
��h�ٸ��0sB^N�%�X�܆��|�o��Q��p^���)���0hwq̃�%�o=�#v��Fl0x����j��G�)/��~�5���.7I�����̐��
n(���ľ�@��a��2w�b��kN�M�uZ�u�Ǆ��`7�K��TÊ�Bз�"�r����}�qS�.�r���|��O��tx_8���d�� �?����J 7�t�v	�`%Έ�B��a�Y��$�V$q�o&�����D���=Z3�_���O9L�4I�1�
aYk�rڗ=�qJ���|R�H��	X�iI�r@=$#U"~��"���^{���,��G�B��1�R�B�Tw��56=�`9r�SwO��\~�tD~0U���+� e�_�3F���+^�R�qp.ի�(�ÌH�O�k����)�v*O�IpM8?��p��a�Q ���a�b�@�Q�6�6/��b_#�Cax��70�*���D�*���+��h
�� S����v��1�ֿݵ�vV��i��,;C�M�����>� Nh�}�
3o� ��»�K\8�n������&$�[�I1�e����6���âLG6��P�E�NӀ���7��eR���P�J}�@�YN_�����ʶ1-�֑�?�����֏��q���*�W>a��y���8K����@$�;=��E���~pG�SP����̞l��o&
��j?7�3�����+ThQ�!��}�ղ#�tH�h[X�[�w}��dpg�@[�;V����V��������څ�&�{�8�����/ڭt�N�J~.��\��R�d-��e��枅2x�)��Zc��jC�������zӑQ�Ia̤�V�n�}M�� ���B�9|�{m-F��BZN���T��˖����~���G@\.��t��4���r�V��Q�&7��M^�мG�[���9w3�2��=9j�׼�l�	'�r��s �����j���I���%�:#d���o����#�X��w>����p�j=#w<]Ξnu�*�W�("4XaG� :Zt�>_:��g{|�(�����.a� }DTV3�@�fF�~t���k֎�-c���3#,��F�jm�T���8�]*nG
}�$�|�$�Ϻ�vȆ@�=��\i����t�]�(Lx�R� 2	�d5��M��M���9ə�[=�����(SP��z�[{��ʷ���s%n���{e�X1y���|�� y�T��$��уU���"H-,��4CN�kF�c�,�&~Ɇ�����aD1��Z��kBn��m�����=�	���
�0ϣ�Lf�'��q m�y4�v&�L��i��;�5�~~�3A�3�\���O֋�>�=�eW2F���"A�N?�? �qw���n�>y�� ��,�VԗC���RN��ʄ���y�tb�����l�[�$Z�qՆm����e�m��t�8u��V<�z�<5�V����u�Z��߬���������3��n}��W�>N�lHT�L���`�������!���[kw{C�Ad#|�gkl;���-���������9l$29���]0R>r��-�P��p�S?�M$�s�@��I�� �_:ӊ�\택���XFo�-���V|���6��P��ţ%Ө�o�����(���C���"lh����09����]K�����<g��H����<0��!��@9p#����dgѲ~�kS�����%�6�Y�٣o�%��)ZʬZ4[[�bTR?��{צ��'F-$��;�u�G�FU�+Z	��U�����{wr �x�șU��B�1s���t���Р�	��zn�5�]��CoaFi<�ܣ(�cԈo�ֵ��w��j(2��5彅R�B�-�����Y�*R�d�6曒Ii����j����쭧1�H���]SC����a)V�_��\��O	0'��x�`����9���mSN���|��%��G+��(F>i�����y�ٮ|��`p�ƪ1��/��5�(�X����r���$x
����V�Ľ	��碏�����k>���� �G�jFI�A݉��S3ݲ=Ae	�U��X�]�#���tz+�YF�֪���<��1!���U���G�i��Y�H��P�;���{ꆢ��	I�}�/N���}��I�����5�2fF.�y�W��~��~�T���濚��AB�GJ~��oǟ=T�&�s(H�}�%�pȪ������v�,F=7|�Y��j;7�08"���+	��K�bwNy�
��:�R,��9mVk~ ~���7��ȥuH��{���2'�)�S�퀐�RS54��F�2t�O��wa&�ؙ��Ǧ9�'���b^?ŝ97�6�����$�O�x�4�V@���.k�n��%���,�Z��R����w�g֯sJhq��@z�9[-�ϸCz�7��RQ��X�V�8)��ĳz��w�kcH������&l}΄�	+�S��)XS(^0���&a�o�;�t([D�;��H?��|��=�
�ԩ��k8)aLK��HwoB�,K6�m,S���`3���X.B?�S ��^L�*�j�62Z���W[��خ[	Fp�w���*���>���\b���If���rU��w7g*B�0r5O&j8,:<�=M���Wc	j���G�a!z�wY�8Gf���~<$-�f�2PC4�z����*Tǂ�L�u�M'wz�Z �{�q������k����{ q�n�sEkNt����m����rc���e��p����0���v���	v�܀�>q$xB�Ɂ�o�f�2�:wW\�vw`B����F,�Sk��EdV��Q��W�8j�s�d�\�c���t�l�<5ssc��v�YG]���7�Xlf9Ѹ�e������n�z���6�r��B�������%������t %x���S}�!�R��F��#���G�1���s@v��K��Hi��f����������<y�)�.��� ����ҋ_T��r�۞�Y͑ c���{��H5I���B�x�3������#����Au���d���Vk�Ӱ��;�di�w\/U�E�/�O��}���-u�c�0=���A�Ղ��%U�6W�`i������oo�L�������R��
#@h���f��&~�^�&�yKhy��́�Ђ�w�1}��8X����-��ڎcֽwz�N$���:��8���#�ӽX��b�~����Cg�/q;����b�.�I�ʩ���h���dC��ŒH!ͧ�r��U2���߹�_,J�ѾrD��!�VmF�W9e��V_�इ���J튁��=��k��yJ��+��+>��<y�G��ȵi���G(�$�ű�H�����Q��ox�+��םZ��dTew釦�%1Z��2��L�e��k��ƟJ��#�S�E�2-{�6v�0��;���;^��ٛ(S:迹��ğuI`J@VK s;�]�-����έ�-2�~`�$]}�r�*Q3���!�/aD��� ��ݼ��	�tj�DZ����j����V�a@ˍ���%V���+�}Yɬ��d׌.�:;��V[wPS�er�Z�pOg3�j ʴ.�� NxF�O�p⨾�C&�G�?���b����h�RY���������:1�H	��g�u)�"9wI�Xz�gZ��|�zlչU1�;z���G�A��Fd�ɗf/_���)D��"@�LT+�;����U��W,��i h��)�g0�eT�1��z�3R��CDبwm���_Ȅ�����K�=�J�������s DA����jT�PgZ���Z'���� H���٩����ג�_ZW�gX �3���{ɮ�eN�ɴ���J)CJ��뾱aM�I�hb��wZތ>K	�m�_��*l��Z��5���(�>�a�#{�2��3�#}���7�CzQ�շ��?�gr���a�
E���J�R�\�>��##�F�&�,*ْ§��-z�k��0�:����Y'���0����x�sDxL6�K�Fa�O���l`~��c#�˯��b��O�o�����;_��Z��Sq�����P������*������o��t�/n���D��)��!�\�����q}��l��S�a��iNu������/��6��
Pz���J��u&�*�kxf�a�9±�MC�5��Ծ=O�0 �=��'��I��J����6���bl̋��Pؽ��'�u� @P$�Xq�oj�,���;F�!��P{���0jI&���f��*�����V�����uS���S��S��GbZi�!Q:r����T`�&������[=�:��QM��p�V����C62�1sD)5-DC���ٙ>�uK��)W�N:
^ULĦ�L��UI�#p퉁N�+OP;@���cf���嬲�9��o$�H��M߶��@�� ���Ow���m�ߩ���P�x�#;t��du��`>�ĀS�;���3�8��Gs��;f�Do��˱(nU�@�Uj? <�:�N���2�ͣ�K�W��\�3�gih)���R�W�OA�dP��ZZa��َ�t�VF5�����v�RgU���!�n�yI9G��z|�퓬z����r'����r?l�+D���y�O�����ZN�H4i���b6T������LD���h~�-㑉��t�1%����q7�Wo}[	~p�SNt���P�R�6��FO�� c^�Ź�_:ƿ���f�by-�>�(�=Z/	9��I[m�^�b/p��[� (�r1�e~.L6�#�s�."2�����	�	�8�1��Zm ��q[�B[���h]�w:���5C��P�7M+dՍ$��ӄ����_c�h)Pd�q��1؎W�e@�Cq2�(/S�Zk�h�J�!�������Ni��u���f�-��w!�6�O���Z�8Bou8���tԤ�K���q��v �V��\Z�������E��x/����6���󤀈�@g)�7�h%�3�*N�ʢ�O���Br�=�M�O�5��-�ȭ��V";�ueS=�ϥp�(�e����-�������P�.!w*��B�óf�<�����&Ĥ2��*^�c�K�rz�<]����SF�`���T؅���TI��-�DD* >��:|�(W3��U��dw-�@�|-���؊֊ ��ʍG��4���5 't��+�
�+}w0��lQ�.R�V=&Ä(T@ݠ�K\�����������g���u��qaN4��:w����0�����w�FH����:�ց�>�r]��ߎ�2��.����I���A��13$GQ?��l���ӿ���>3�e�H���X?C�pfTJwkIMؒ6.���%5��e�*eO.o�u}���G��|�.�LOA*����x��($�c*k<1r�w�H���/Ցh� �Ct�q���;�9 +W��� |�i~׹�/��Я��>[���W��ٵ������6���~/65��������tj�W�����>��,� �z�֞&��*-PS�D��
{�N��vP��*��L���bW��r�萬=�<�����D�DJ',x����1	�yߒ����� ��2 ~��Y4�[k�ʄRL��ۢ�*�a��&	ɣV��(u�B�l3f��nJ;�m�5�!?�8��BH��d���O�=�&� *)E�ȸ�@P#�J�8��#G0���q� �Vi삒��k*[��������d7�FXc�`F,�?�F�˔�&￤h��\��)�c�^+�l�g8K�_�e�FC4ɨ�7V`��ዒN*���XQ:;|9���!U4�mh8�l���΀��~<��@;�l0�6\�Kx�Z$�Y �M4����BL�H�����j����,���AR����]�ۛiA�����.��-[��w�<�!w}2�³	��fu�/Dv�k�<�@���CWrjQ��=�7_���{�r<9u'ZJ��}�o��ڤ>���aG���˄��t������:Iq�!�S��Tt��h���E�j�&tϸ�1X��6��~�����.��$3����?9���xu�C�w�.:恐kH�,�7#/���$���
�kԻ(���Or+�bK���S��>����t�H�����U8F�8��b<߇0�L]�x
=���)�e��m5}������õ:2��S�1���=�"��򉬇��z�з�_�K�o�.������GVp����Ǐ�� #qw�L�|3��@sTPz�F�<��\W��F�(�M,�x	���r��X6�Ь�x]U~���i������R��.�k*��_��c�7;��X	�p�d;�S3������[��u�-pi^�fAA�VZ:����>���*�t�Hn�B4`-��O�<l1�����(��I&�r/��Z�%�;�g�t,W��@����q���:04~����S=�(Ƹ�C�p;��lQ�%��f ���=K#�����"@>�D��ӭ�h��S��C�\����e!�#�_�KbJK��R�������kO�ә�ع���qj*�\���G=�k���@�eUĽ3��_H3��q���$�6F��_YfXSjo?�Q5I�lk4�}�hx��M�q�d2���l��tG���k�x.�Ҕ�cU��H�IΤ��3��D���~l:�) �bk�E��K�R��$X��$�����v
�ɰ*�kͨ^X�=��H�~���xq�zΆk�OǛ��R�$��Y������ Y�|��b_+����S�
�B��v�迋?��BF��� B$���Ŀ���*J�v	��-dE�9��_b��S�Hp_W�\�G�U���A�-Y�f�(�Y�v���jG�`ںC�Bc
�͝����k�š��Q���æw��"+ICk�,�0�-�j}˥@�rjf����ĜM�jS�e��_j��z�U���pq٥G��Sq� �*Tq�*Ŀ�F��3�k��j���f�#C{�ԣ�4M��d�z�9�����dU��3~)ϡ% ����eռd1�J�	�e91[�#îF�o]�m#��Y9�J�2��!��lf`"
�^�D؜�'�a��T'�w�X
�t4�!������1~�P.dG����	<�<�O�i	���i�������VX8��o(�g�S���FZ�S��4� !`8���F�f9�Q6,P��)Xv5�S.r��M���48�-_���+���&c�U�k�6�������A���2�x$��)��A��T_�U�2������c.G���2�H@��^�M���q���(p�H�y�.6�Qɽ�u�K�y��s)9q��E�M�-LU�u��o���]/�=�=���Q�sz�Ǿ��q���0�m-�����'��?��@��*_�C��8å��=tY�n��#� I��v7ݝר'���	gʓ��N�|AGzxݱ���0$�_%�����k��d_K$��E�sb�u˼�2	b}Ŧ�_mԕ��r\���x�bN��S�f_�Uz��ƚ4�`펗����f0�s�7�@�L

@�-j�1�#�y2����i1�ӱZ��-	ߍC���e闿Fk��:���h��C��E��"���7�ZI|v��]��J�1�ײ�s����c=ђT�y�ؒkcmLsG��N`��?��k�R����jx����G���86���-��*5ÃS�1AB��9
���`�U��E�K�[��U+�P,İ4��G󎁈��r{X�QɈ��הJV�*�d�/T"��d�8�;����e c�C�f/�Ԅ_�T����]yfh�c�c1�&7�:���H��T�p�;���D��ʩ��.����0�[K����t^�k{=6.o�3f>V`I��,~�����ف+{T�nn�̱p����5a��dx�%hj(G[���AI�l {?�! ��8����5.Wa�RC)����uu�#�D�5�t��9��g���<�{Ca�ׁD:^��qT��5и�5�C�R�)�1?D��Gd#�� ���cj��{!��f��$��N�<=�`�D�}�}P#����0B7�͒@�M���;BUc�

��i�%�K�A���g��jޘUXJ�eL[.b<M�� �Q���D�,Gψ���1Ky/��Y�����(��ɱ�/{
���_���9בEz�g.®��ԅ�r�	�h���[�縁_��T�F���k#ڟ���s�ʿv9�E�X�e �e+����]��i�����}*�o��lEd��1�Ge)tuJ4��dZ'5�X!��7�J�B�J�����˕��?~j�qJ����wb5>�[��Md�B<���DkZ}�k������g|P[���������~e������F~�5�dl�Dq�*��	~��
,�,�}W�������a\��h�^���s���T�w���X�I|��.IZQ,�ؙo�?% �.&�6�,�����6u��!���8ķs�/��]/ �qB�>n��6���0 ��ۦZwl����}ɱ� k/vߖ<d��ug���B餜��	|DI1��i^�NӬ �vny6^�����S*�SN�_  ���]��%�K��k��kL���q�oX��\�j��NG�8;�5:��M S�l0�ȗJhl
4���䠟h�D�ۓ�S�,��?ĵ��t�� �N��+մ�e�|�6׽R��Þ������K}�,PǙ�n)�����r۪!⠷k �k�]�&���TK�]1��e�V�ek����MF�!�/%�5sf����5�:�>[�`�ȕ�"}h�f���?2;w���6�H�5ܟ�K�(���Y�̓!P*V�[���K�lW��Y��rh��HWo�!]^NL+f��5��D�#>ݟ}V�$��ec�BHe"�X�V(��ll�j�`&��j�w]4JV���TÜi���!1�f� �(��� ��.\d�Ę��(�{`͵��w����$�jQN&}�DZ�d'�cInXp]jLԮ!��ͯ~
�OZB��@'�6�$Konn���!�#��p�ES��2aks�UGmݬ[�^I�-�虗Q�b\O>�VgHLr�4�����"^�+|��B�<a�n� �U�ei��m�N>�)�,I�?���]`�I@^���$�!m.Ǖ�4j�%v�=p��"쎡c��bQ��.�g��x�@��g?��nJ^���m���C�2�hA�����"�u�(�w�N6�>��v!���{	% �s�T���)����Q�ʙ��%�����|�hQ���B���:�b-t��MX�D#�«�����P�ZPx�c;�4}�)�����Zr樤֮������~}`\���V�ʰ9��mN�qs�L&�޳���~@��/�e��<7J���d�hK�D*g�Y׹��	���1$W�Є��~+�0D�>_��lB{��u��|C�IW/gz_�>�5�6V]9!����b4&z�}�<�-����	w-���k;	1��(d���y�d�3?� ��m�4jd}�O��V!�.�R��!�	N��Q�Sd;�M�]�x�Vf�uy���T�if�sdw��8ōQ��$�7���a�޿��R�Ül|χ���h0(螏-�@'�6����&��&��VR,u/w���	CBƆ*��g�.�F�������o5���saa�@����>�Y�����舰\�p�e	������� 0��D�_lxᄞ0ږ]�ݣw�7�Yǟ�DZ�r���1P�q�b����)�?kẄ�؆4a«��*6��9P�#�b��]�*�#���e�dI�xGd~ߎ��y u,�Q3��w�ƚ�ؐ^�s1{���Q,_{��4d�	�uâ8-�,�M�[kɪV���:��Dh�S|8(�o��q�f���q��h."Cp�!���~(�'0I�gC����q5И$%i��#H�%^��P
-�&��C����@��X��B0�J��z�b�9�)�X"I-���݈6j+؃;�xg4�����M��a�Q��z�&J�z�t��1�=Tp�eh�DB��/�;dy�j���͇+bT"�I�V��y���rA4e�d��#������H.R8c�(��2��B<=n.��j�CHk�D�;lf&z�#
u�A`�m��>�}�Z��37>�Q÷��Qr������ÿqUC=6t�|�=�j�ǫ��������Pd��N
�- ���`bY�`�Nܞ(G��7�����g�oR���;�!*mjz�H�%�D�h`iP���z�N��VI�.=�
C�9 Σ� �8����L��)��G�K/)�SW��mCа�Շv�4�/h�u��9��K��H���y�{'��p���R�0ؑ��n^���)Ά��?"��D���Q�sH���Zԝ�H�ԇ����H��K��O&X׌a�|�%#��H#�7KyI�5�sh�_'�;;�7�iw��"����E�JQ���b��v]Z��"�(2h��$�?l�!xsGn�'t\�;�%�Ь���d�E�+8xh�ܔMɛU7H+��v1��*�jr#�u6�Ӣ/Z��g�k��ٚ6 hkgO���&��b�V�Y��"\�mrU�*f�g����m�(�o���q��IY�<���ـ���{a��#]ۉ���n�+3�,'7ν��O��g,���AO~+��_bK	��]cR��M��(��=���\�xg@��fC�1�����q����x�*�]X��W��1���!(����@�O�)$n|7�~���?I?!D�9�~e�� �WYR1�_%���1�n�W�u�:�8�w�كp��K�3ŗ�a^�ʶ���T�Yi;��~���0o-1�6�������y���8,
�L
u�L^_y�N�;Nb��џ��GV�_4��?W~��N��h�$���F������`d)���-x��.������e"u�nμ�b���w���$P)����83��⵱i����q�;&��R�O2c}n\�z�p.��m/֤	����D>~�N�Y���sղ�J�&�t��N|1�g.ٮ�<+z<��4#&��Us����/�2Z���y�f��?b4�bҘ�����~
����H�m\E:%B��gQЂ�Om� ;��)M ��TVD���T��[&�8��h+�I��`H�5}�����V/%��$���?�q�$Z0�A��I?c�i7V�^jLRXCŸ*Ƶ_^��C��4�t��)����<���/Ë)���iN��;�/��4�nM�J胵87_	N9#�%�1|?���N�@2S.�`Q<�U�QV�첓���"���s�`�b�"�O��0�F��]c+��"���ϥ�mx�kyB�9Y��`�Gƺ{�S��$��)��{+#��H�ZQ�f���T�	�Iʻ|Y��Bb�8�����s�P\4!@!����8�U�M\d%���o��}�ji����|�HB�� 3��� �%��t�E��x��+ұU�X)9��H;uӡ��8�����uX��'���Ɖե����>A��r�ƒQ$Ӊt& ��- �-�z��pN@�y�K?y���i0�6��fZ��5+~o���Y���٥���9\���'ъ��k��#�\`x$tf3�`V�9BM�c����x���pdW�DLL"��h�P��?�WӔ�7�L1��[�9x<�����|>6^�!���.��e�J��
v?�	��̍*�Z;0@�ȴ�π�辸V�g�y*{�d�,p�D�3�k!J^2g�.��p҂;s��# ઀����m�
W��#��aB�"�e1P�(��I!�e���ҧ���`�AV.�J@?PDD�'���p�)V��Ŏ/�B�n�图E����WKs�.�@5�����;�M��p��ί�����yfPZ��_Dw��R�Unڲ��U�%2���O��,mp� 0 qb��_����)��֡']���4�1�/��t�@.z�?��W��a�N�z'��#m�9<Q���,(�\�;�,�VJ=o�[k��s�jT�͞;��P�s�0A��G��N�����'l�Q�剗,Ot� �b�	Շ��^U��7{S�c�2  ����H2z��J�Z�]�3�(�!�zw�;�G}/�����7'9��m�k�1Ò�U#$g�U;�F���(#�ݚy�1�QR~���)b?>�c�M�t��5�,����(�F7(\��љ1s�ޘX�-��m]���r�/x���t��SY�:�D�����_��J���g[�ۛy�~`��9��E�.��F���g�6x�֒��!��(��H+��RU���;/1"����� *!�3A�.���7��<?P4OH�p�Ľ���D�EP����Б����R�f���j�]K^�{0���#eՍư��ųz�[�d�?�����Q���;�d�/�u����t���V���g7��+6�#s}k��yb*�u/���� �9�������O�����@j���$� �^z�L���wU;pST �Rɛcjd��s7?
m����$j=��ץ|�},�b�-`���n�	�=H�槻Ʊ�
os;'��G{c�d�{h��`�Ӣ�5�꿚Ϳ "O_�\�+N�9�8{������P,QS����6����V&ȣ�<(�=d i�s.p�΂
��8w��;A�C��գ������È͢��F|��E
�\�x�GC%�?�Hw��V۠Ci��Y��q:;c�h��_����ɵl�J$��� �C6���g��{-���0)��P��I펈p�ODo����	 ���X��|����=oeU�A���/G�	��'D��闦qfXv�)�w��}������7W
nnf�M�֗�a�w�O�c�0Eg�j=��P�+k���Q{fk ~z :7�-��͙dy�;�/Cm�6��h����FYn����W�H�o�4�g��B˺����݅� �y��6����0��v!$��BA8Wh�9����[�Ϳ+��ʟ٠�$_�nW`F�����Ҩ�R�-u���}��Yͭ$���~6q��/E|������+��p�75��q�<�󘟩��U(7�fa��@�8� ,���� �䤐o:���ք���ͨj;�cm�ŗ܌ţ�`-�th�k���䉉4IYy�`l����5�X )���,�"�jcy3��P�ݎ�֣��'��	zܔ�X?���?Ń�o�