��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\�$���� �NE���D7Pp��\.KY��s�����F��a�d58Pֹ��US�{��!b���Z��z�lH%/�K4�sc�̙�qj[��������j�U9lwCOw��C���mdN�s����w�n>��A�Iα*���+Yq�̰`Sn?kpx��p���iU�"���m��0��e-1[UJ������N_Ѧ��.ht!I�p��;79��of!�=�n��Og�y�0������J�v�����<�Tfj+�������ZX�t�u�*L�$;3� p+e|Y��pԝ����N�gb��&�sRWiX%nY�4a�. �.!�_��җK_w ��3<V�DϤ�����N3�ZE�
��Qh�2D��N�Io������y���
��ۋ6���V$���G�5�X�gH��) �����"��S���4��[�+(�*S�jM�T������&��9m7��~�o{`<S'O�h�LA��bKE2=j��)�N�gD��'N�_G�D�lw�]m}8��)a�kKjhdq7'`*��	�w�	����Vq��GC�/Я)GR�g�X�N�d�Κy�+�8a�tS�Ƥ��0X��Ud%�{<�G4�=fE�R;wo������)ϓ)�l�0�Lu�68� �V蚕L}���zM$j߀`��q�(�ǯ��wꄱѭq�������84��rϓ� Ǹ���u|o�`���X�2�5׽~�n����J���H�9R;�J����$���]��F7�t\F��� �+4�cd�
1�G�E�Q�E���[�dp�I���v'q[+U]%s#Ѿ���Pt��{�����'��Լs��e����7��/�[�/�q�#�f�'>&�K��o;�iE�d�3���W�<�B(�����gA�62j��e�[��S���N��NS,�,��Ž��/J�ɀ P-�G���[��Ԩa�"�*�%e@_���x���{-�ۅ��+�e��P|F1�!=w�k�6����f@a�Y�����m�0���j�4~�D�l�4X��v0�[RZk�'�|�~J'����W�ۻ�KCE��Y��{��(,nshx�e-�ķ/F�{b�<�_��X{��WJ�8L�A"�au��O..(v��yW�UN� 3�W{���kԂ�l��$��As$�ʾ{�������S���>#�ƻ�g��J�{1�a�ZG����q'�ߑ�6���F[_t���|J�_׽B�*�Fq��1�->c���~^�/����&�D7��xi���5�Ԛ��������N��#��7u;�쀊��͕?��^����;-~� �d�VD	*�b�HbB��lqF�Z��rt+�
|̃8��;Yڿ��_�R��ٺ+���&_ԕ0q��Tk0u�M�z��O���q�)��s �T��Bp�#Z�cB|�Ж�Ji�&�k06��cx����j��p�9e$�Ƙ�1�K��G�le«�Y�*\�����Fy?�#8���S�K�Å�����b�vs2v�=i���iA�;�f灚��_RLicb�%]�;�V���Քr��Moź$9K��8#��L� �n�>'���MK�����nc(
���M���}ֲv��5L�[(�Ƕ�btv
e�ӳ�E&�T3��Q�1<��hf9���[�e��������q'Z��E�����Nmw�g�n9'H��3���w����\���[pa���^u�8�m�%�q����7�������@	�a�%��� Rq�$���蚽���۸rC�i(w7}?�o6V*���jQ�0��� T$s��{��?��+�E) ?����B�~���{x;�]�c�q�������dx1����*�Uu�5:�����)c �5Wd�-Fmi�{���4W����A�s� �t��������Ӓ�����e��`T�=Gdʥ�I�HصBY"��s��O��R�:�gVb#I�2
2���F��cDg�̄�'`��E^$�0�����?�a������W�ccNZ�S�lq�������ўED����?:� �e����Q���Z�]�im����k�w&6� ����ݐ�7a�Z�JP�v3�X��ɖ����ɨ��QK�*Y+0�J��Y��n���M��u��r�y��o�/<�K�����]����b���n~S�-%`ɲ� ��7j�Zw1��Xg>��y��/�A���9�CF����	_��R��b�:���HS?��e�]�������i����&ᭉ��ޟE����ϡ͹G��!=@F�M?G�2�e=~�z"�ӽ�e�a��AUB2!|/q�������=/�^w�G�i��NK#��7�>�ڭP�F�9�I+��k3���쵶8ߎ@��9�tR���7�Q+����c���~��P�H@�+�����.���~���t���B�5�m�$�S��wy@�:u[ݓ/�X��X���Qm��d�	��,�E�2�>�F=���[E��u�,<��3�
�+@}�&� �ª�`p+B�u�ͤ��/�P����!)�˘N.��$�d�������W�l�48-�$Q4$y�2,�MFoI�sN�T���>O��8s������\�3pK�p�/����u:Q�2I��7⡻���qW�v9-<�(�8t�8݀.���>?q�	�-�y�eO�"[b��h��`�C)N~Q5��P����\��3�	�C���tT���Qw��<�a�zav�4���~�ǩWnBu]�)��X<P�fm�����6��2�K�:�5I�]E��|b�#eW�ƻ��Ŵ�yU��"�%���(�U���d�錇����(l�b���ɐ��h.L����9c��)��1�Y���~�����em�a��s�@�9��0��%�g枮��P�qn�;���'͕,zY��bݞ���B��^������Ai@�7�f�(;�9���v%H[����Õ"<$d�G�kL��x+	���9y(f�
�LN/ ��8E	�,������11�a�lt�68%'���M��)�pk^�hŚ*�Z�Rs��L���p"`|��e¤M@�`
����@�����Rq�%����4o4#z۬�W{�gɰo�&���gsE&8�g�O�������8��c�0܀тu���e��WG�ZN�Ӝ)�A&��}ɂ}�!�CGɏ� ��[� �m�0G�*��u=R#��e_�R����q�g�{�2�8����Ĕ��ޝ�A���� �:*p��ٜ�����`�A^]�-{����`^Ũ]��n=��{> ��]�d54G8�Imc��7e�������Y�+��;������4��zL�x,|�%3�W%�.�D��g�3��}S��۠��r�vMG�QF�
+�H
� ʍ���-	�U���S�Ⴟ�V�Jns<�S����X,�tf��uܝHD���n��kP�U;�B1t�����?7�?w���ٞi6��v=+�pAW؀L�����A���_�	刉��Y������i�Kс����h��v���0��C��;�zŸ�
�QI�jQO~��������a��b4��X�iaj�Y9�̖ݻ�<����u�g����u(�e��{��wC�ť������d+	`JfV��UH�����[��8����(�2�ȉK�7 �qmn~����B�7SL�-#�~�):�E{���`�"��H�,cC�}����W��Β�"�+��5�>$'T�}n>��'��Y�w |��(|2�Q�)$�k#X�z�1W����AF�pK5{U0^U>� ����O��c��Z�B���٣�kn�Ύ�+R��k����$/��.8�����M*��M��Q���rJL�����r��{"P	917�O�o�1T�8!9�.#�� �&�W��s��Hx2#U7vS��<��J��Y*�.H���0���2���-�d1�k���4C*/ƕVȘ�W�5ciXe���O43��ll���]�)t�걜�4�i�`a��ͦ&z`��#مb<��	�#�E���RN��5@��s�3�ŋ�I������M6b�s%N��7�z<C�>��7v&'�I!R���s��+�!-p��p�%و����� X�:o?`:�t��ԣ�ǉ�m�����ok��W���l.�>|��1�wt�&,r���L�ʛ�ߚ����uF���I��/H}���옮:y�\������8!�d�4�&h`�C�?��?��\��e �� ׌G���r�#E'��E~���Qhb��
�ϔ�kě���kt��fó��5�1�ޠ��s��~�􉻮����k*>����%4"Q�؅ǯ��`�g�n���b�\��ˤ�,�߹2�4���'Z 2��z#��8�LqU���W�M���"��B�v���"�&��7.�P�-�~	�>&l���)�Y0E�PŴ͏���kS_8k�Q���j4��3:-�}�r�̵��)��c���L�"�"�Kyy��/9WǹGTV��,Y��w���qz��c(�O���f�?����"{y׶�\�8�w���0�.�m��h�<�GW�4���w����3��"�d���s�����å����6����	���J�U�J����=xЩt�O����vO0�pƭ�og�T�K���g�6@a�Q2�
^}�}�FL��"���d�.��0�b�j�pW޳�Y�ވ�ۂ�-������NFY=Ě� ��P���J�mP��_�j=b�eCg���m;���ڮ����1�IwIж?���9�Z5�#�`N�v*���������tt#�,������܂�F��W����˭��;p�iv<��� K��a��,#4�98t5f�~�zw�L�c��D��Yx+�����>��+��?�P���~B�R;Q6W�����2���D��#ͺ	�� ��1�21�b_q�%G�_�P��3|�qGr6&с���k�����߉CuՋg/W!$�~UT��9��:���J��Yj�Oʭ�q"� f={��-m|Vf�	���E�{���T��F���!S�R�$	�E˳vB�{+��}�3�%9�\v9�]��&��l���b��O��	���u<�D�yʰ�	�ܟ3N��޹���~zr���ߏi���pv�T}�>��BH}�x����m+a���6���W���>UQfLoZh\05�	čPE>��i��e�XT[�r�T���:f���r-��=�Tm}��$��q�dQܶ+�p9�8Y�����C*P�����ݘ��T�t!�s�	وfF��}���D>��OF�/�6�/�7x��dt[�� 	_�e��L�H�o&�Al<z^��<&���Ƶ׊Ho�=vYR�Z��r=�&L�42t�;95	��[z�=�t�ٷ]_X3������`%d{"����h�btDrV⊤?E��Fd��T� �X�m�~�]E{3H�\Hso|�~�&I(YH�l�E�{��p�9I�� �2�1�*W�db�]Y��z���vZVdC�y&\v�#+��z�T7�s����CB��1f,m��&X���������(�Dh��/ Z�ZO^C�'�A�	�x?o-�z`aRv�d��-�Ld�Tu��������D�'�eX�ό_0�G��. N�g��
�7NҔI�@��~��6��[zX� ~��������KU��oɲ���o�'�ŕ�8Ů���Ƥ���nU[_	�?�,b�x��z��4��t�g�ٷ��Y���̺('�%��?8J��͛���G�{[`�]-c"� c�|;t@�2���91��%�cj��kT#�Ñ�?d���
ZI���ɨ��.��B�PoGTX�u� �yJ�$�Q�xL�.�������\�S�H��q���4gH���m��u�b���?��g�pg��C4��>��В�o��j�~4�O�z��$[�uc��PM����r���z���sM!-yL�O�_5و���2���Z"�:˷�۾$�׀�C�8�h꩘�@jm�m��$�s��3�d�� �Aq��(�����(�do�i_�x��2����d�?�N�hS;&���1$���(��3LymM�Ҏ�u/����#���s��q�=laq�Э���� �4+B��'��r�#H���M���D�~���Pk��Xn�BL]!|s��X�t�@���'�,��A!���%�}�&��k��&����"J.�OȄ� ���5����4�L��]��w�r�U�n�>�H�8�ξx�L �Է�/�J�膄�g�-+�q���� �2O|�%��e�x����SB����^e~ſ4�+��K	�w�h6e�6ſ��4���(Q����!	�ͦ˅LB�P���O-s]�2?~��P�%����e᜔�B��,[N}��A��

�ؒ��J�{����+�3�UMΟv�!x1�;����FuKxy�řR ��i�D�u��� v�}��7�#%��.t��S��$,�`y�a�_����'��m:��q[�wA���l,���qy�����^�=�$�(��6�ȱZ8\��oO�@|�A�_GTs6 i$JR!j̗N�L�&g��	2g"�Z�v�/��T�L}�m W���� ��q� ��b:��<��	N5�]+��f�����K� wo�Mܖ]a4�����\6`v��l�Ʌ�����\b���N�������ǐemX�lq��0��ABy[������}��P�$�n��^��w�+� \�I��1S��Á}؟2�g=�0=�i�s�'m�ݩ5avF�A���ex��q8k����9��8IT�rl��K=�kxZ̪pL���F'�L��P7�w�b�M�#U?����	�Um#�۟hC�s��y
eM%W�U�`�b���]!}�m�a�h�jV��k�E�L�����V/�:L3ݴi�A�c��U���e�L�uGs0���
j�2�������)L�w���d&Q{�O�b�d!*ttO�)˸`�E<Hq�������șd��������I����-4@��I��~e�r�$�tUP��=��%��cD�?R��`��������QC���H�8mp���t��(�����T�}eV%��avV7vvN����)]��2�.4���zhY�h�jT ��?v��%�Q����rA֌А��P��:q~�=�}�7 g��,��MG�ͥ��)����x��z��.���a֦�P[`���cݨ���OP8.�R1��=@2����C���� �)~BN�N ��?��.�oZ'T�.�Я?�uJ�=�/�7�;#~w��=o�T�}��W�̊d�B
{�AO*M�Y��Fe`��E�1'��ޔZ��r�Zk��,�����pqgh}�>~�/�m|�Xr_�Y�z�6�©I�1��}� 3_���s�����r�肣w���P{S�4��8�$/���g$\���C�Yyۨ>U����w���V�TpcԨ��_,��
(���=Ӄ���UA?�x�ŖO4Н��3�a�C��h����i�|�5��ˑ���˥�R�%�t��O�Yan�+���$�2u�����3^��W4b`,z��@��Jo5��?�<j�o�n0����O�;��;ǧ���Gr�,ȨA�\�lտY�29���@��a��{P����	����fg3YQ�0	� ��Y�(qB(�ְ�6� �;J\�ҏ�$��]��m.w�R
(7�yz�|En�f��N~^� ���x�s�]���~��?��j76F�u�5�:;�!���5+j��Mo��a�$�
��0�,������V��O����Zq��
9-�3�ntSx�Qō���M�v2�/�ň?�61r�3�v�0	8d}f� mӯG-�y(�)[2K��G �;qX��i;0�)���_Yt<����.��ͲbL�HW'�#S>@�Oe���m'M�� �ȇ�a���퉉u���I�\Oy����E�Kg�O�v[���M��g]T~�^�R����4�N��b Y!3�Ո�a̒��H	U��Zl0m�%&�:^�G@��8g(��L����j�N�ج�f4'O�)�xܰE�W�$B�Ι��px�0TY}���񌇔=��?ѷ�9{�j�c�0��W�R�{9&k�W��[\<��z�b�|HWkQ&2,��+�O�#�u���w�dS���lPQ��]�R�N�0����/����]c�k@d ��/SR�lO���</E�b�+�q���BE�J��5���Tr5��
�T���`f�s���oR�Z�E+��o3�����tٹ�Ⱥ�Eܭ�żv'[�˾����=/��\J��wx��$���8|�*�ȃ�����Rt��"���8�����Q�a�	t�H���~���,�g2&��i9���Ҿ��	@�G�,5���U
^+��H�vVu8+�>���='��p6[
I
���)Z�wG�E��Xܫ]��CG�����Q�;Z��H]S��]=�X!�	L̏ßc3��M��.�o�`�5�Zvr����	�)L��]��[������5�>o�/�����"��O!L�@�r�T�9⥶j���4�-�%&�ta�Id
	ĕ3x_�K�&W4���r�s��O��`�'�*�M�m���_� [H�q,�tw�@��S�)'���b/�F|vlӴ�C9�����b��߭���NJN�4���(N�%�@x�����Z7l�#�)��y1��<%�C�is@���u���hRd�Z�.���E��Z�ElM�L�Rm�P�)aZ��A�23�yz:�?��8~k�uzS0Y��ų�k�:�j�����N���֢�#���8ߚ��"@��.��v+(�9x����k�t�)v8��X.ZC�/<�YZ�o):���A.���qN37k�'��#·�I]��~3�o�ʴ9n���/�6N���u����Y!Ǌo�y����V�10�@��9k�Z�7\4���wV�fv=+Z�8J���r����������#d`��2��*����gy*�7�@���k�,#���
):�~:BfG�:�)޵��1��yc$Qo'��jX��]�FX	7��J˨�{0ʴ�?g����o�=�\C����]9�Bã��_�N?ֱy�sCT�����Z�r���N(5�5_Ǡ����,�(��s�&3�^��di��7JO�Usr�J�b��{�x	��9_��J�b��M\PI���(��ۘ�n�74񍆷zƐ�
�j	c�W2�`&AW�i�@R`��	�&nħuaY�B2��E�d���J� ��d���W�5^���b&�*_6e5N�S��RT���S�j�н�_?Dɬ���PxW�(�(�g�s��DMxTq>z��"�1��md=�Bx
�q���y���P�
�ј�Avȫgi4�!���Ұ�cN��.ڊI���1�'_�?ɲ�Z}��E!�74v	�����.��ZsD��	�$!ۚ��|�H�FGE��
r�xѩ�P�L�qc�}�=�BKT��,ք)���$r��J@��kwΚ��R�j�K�<�;,#��hдhb j�O��#2P�Q鶯g�qJ�*ܧKπ�oCG��0(��	�CW��0I��'
8���X�4�մ��A���2d�� -�^�W��m���W[},��nz�����."_fP1]�!�*��@.6Ju�TgU��Ľ�N��`T]nJ���
��g�rK�G�u�q���%tV+�#�]�G�Zߐ�J�L�ᙬ�-�!�*�> ���B��Me�UY�~�X
C�� ��zxf����v�:��(4%ݰO�����:��*0�P����>�U$b¥3K�S��AQl�'~v�	�X�2����N>�~�z�����\p��!�T.��(���3k!\�s�;�Fd�㮗vw��)wp�;R�:�B�'�nTPB�Џ^��h�Ӟ����L�T<���W����&6��U~��щz�#�;���Z�x�T���af�Ni�}�cj���Q�� �k�KTrL,gr���ώY�Ť&d��Yv.�d[�#��_#�����^��DI��o��Q���1��ܧ��q\�����rd%��䆉5�9�7OF"-!���t������?m��?�Qr>_�O��O��[�,I�X)�W�ꃹ��i�p��[eWpa���Ƥ�-܋���t�]�?YҢ2��R�XϒÃ�þݨk&fl�zQ$�W��'fq:�әc#t�t����j�V���&�9�q�=�r"��=�:�z�ﹼ�?�X(r5 o]���
�S�v9�e]XVF�Q�~���>>� \:`ܨ#7=}$��g`��TӀ*Noi��7M%_�C�H�O2��~aP�@�u��0��6���蚁�}� �N��������`iT������ҘZ=Q���"�����e�ė_���:�v�*���K˘7�yY;�;���9��[��CX;Gޒ�*��wbxƝ��i7E�I+E�rKZ�Hl�����ΥjR� 8�"�2�ݮ���ЄC~���f�[׫V_a�clW���$p\c" d�<�D8V����c�!=gR��y���7�h�/����sI	̭8�d�=g)[��N]�Y��|�i#W�&˚�b����[�l3��:�;�1�wgY"_�>&��X
"O�6oH�� �n#�����sG�q�\�?�c�:g������p%e����eR7���KB!6SI:���Q��9|�ڸ���5�}��q?��n��6B�$.K?���::��w���Sb��	J�g?���J�M����Q���(��e��|��k(�y�/���0"ܖ��R�/�����́Ȯ��Ԣ��;�h�� �h@��~�"��1"�4÷|�'�{����'[�/
��vN�Cc	~�Jٌmg5��a5��8������I��нv��E$t�D@T�Tݘ�|�ފ;(���i^rm,���:��y�^�g��j��"�8�H�T��-�: J�$ˣ���E�#w���r�!H��[̎�w�'118Y2_R,���N$&jfK�7�IL
����*�*8�oUgҗq-����:��*�;��1S)�>�vN���'�,	��
��Sѩ�ij�Z���D�R��I��S��E���
��U}D:�N�P�+#���������|����  ��)'>e0�Q~�-X��V�#���sݷ9Ri��Q|�_I�Q�X����],�9l���Ί��w1�%��"�	i�k%c|�岛����v�%���t��+Ϻ��xp�����-6�\���U�!&�\��X�Z��ᯭ/Z?�v�6SnG�!��/�J5�����ߜ�k$h���"�Pٴ�Ǵ����♸�c�Ax�ʤ*R��8�ndF%*���Y-h2�o �_Kϧ��{�9��szl��}A����<�3jGtt�Hj_��-������������7�{�`�����p��KW��|%M���2��A�c�i_�{���j�c0����	��mGy�D�tG���U��8V�O��x��	�i��1�v�`�~S�h�����Q���$��,ؕ ��@��;��8L{b�W�\`c��7�#�E��d��S����R������dm�!�X��=� �ⓠc�|t��n�gu	]h!�CIZN�����.h9�#}d�����*���`��$�
�I߻B�z��t��[w\���:��/I�I�C[��z�K�L��x��Qxl|��:^
n{)����Oiy�t�)9�?Թh�|C��y����]_�T�</iBf�	�W[���(l�Xr#y�BK\]
��>WZ�Esy�K3,��fzF	��<\*Zu��Ryy����+�r }����C��5$5�JH����B��<�^xe��������/�ѤŚ�`�!f�s�$'�F��V]4�Y��h��4gN�9T�S��y>(�p��Q��<����*�U;�һ�/�S
�o&��yᶢ��<�(`lH�6r�LJ�	E�=U���SY�]���Y�ۆ��Yf���\�ę���O�W!�c��� �ƨ"f��rY>�M�8�-;tc#��d]�����P9�=�"b� %�תEbH����`���PD����9bMQRp;��f�&L��8�ɐck.3G�:��4��7�k�m�b��T�'�ei�A���w����3R*��8̾G�.�JGj!6Q��+F��k���q_6���Rӿ�$ŃEJ�y(�9ź�)�i�G$�]�)�hm6���V5����P�v�K�xH��p+\�l��/��}0�L<\ܡG��������m{6��b����������<]�Bz�r�ù�Ζ}<��g�"�s�y
��Z�1�x����;M#ͰZ������!Ѻp�j�4��{vq�UFw����*<�$��F����#Z�'/�Զ�o�������[QaZַ�N ��K�)҃�{n����s A��X���᝴�'���K,����Ʉk�ٗO�Һ��ƀ���p`�2�S�**�$���bxP$�}�3�.�^�"h��'�H�vz�,�Y��2��:�Sv��w*��#���n![��Vr
|��8�\��w�d��%��V/�����v%D<	�6�@�!+Zq�Ǐ�fԜ�B��<k̥
*3�|g��+����%���`����*�ܿ��v
��d�	p2Ǆ®mP�X������]��De��w̍!�G�8��N��!�ٱ�n	�[L�%�[9͊)�2���ھ�I��b5J�P��ʶ!)����ŀ�&�_�-��Gth�L��-���.�d�r�.B#S�i����e��jn�|��8~��+�W��Z!�(Pb��U��w�X��g=p�f�/w����m�y�'5��k��$���f7H"�]$!�H ��viX�y�$�*�L@��!T�Ů}�}ȩM��������;\T���& �I55v�,;�ۊ)�-��`��US�^��E��68���i�B�Db���w��Y_��t�A=¯���@�&P��$��	�PJ�g1�k�m�>�һjX�>�4��O�Rq���]~x������{2��-墪cz�6<+'ca�@+:(��F"$�e������B 0��6�,�W���w׀~
M)�Ŧ�V{�������Z�~�T;_�����\���g�i[B	Xv��'$�֣�nЗ�Cy��XG��E�S� 'g7}"����ZX8Z�RuE��q�S��Zr�����V�3�ʯ3���6F��9�8�c���	_!������l7}
Cp�eꗔ�s�h��e�����e,�o$v�8!�$Dv��f�+j8\aQg�qA	΂��s�d�7��^a`u�]v4��^ك��w s��7叺���!Gµw���C�I���h�J�Q㝑.�E����YX�I0� �R1�P����ި�2b`�im�$��&"p��m]O�D���0v
(�߾���h�\�̸��2�+����@>��P�I��!Qu��ݹ���hk�&!-5��?�� ����D�I�=��Q�5g�$�Z��XM�T"��R�י�ZV�G�>ƛE`�����'�Oş���9W�n�YR� ���I
�r��Oԟ.�����P��niV���p<�|�r��`g@>�}��Sω{�2
��j�r�X\lj��)���\�ˆ<�?0��!�ZU���!���+&��4+-fךm����Ϋ� ˛z�˹�<dzX��������2��8C�@ǂ̈�fp��������v� 
�)h���8�v�0g�Usi����S^w�Qe��J�`^m�I�x�ِ\J�XN�5e8��9p�W[\q�G��:�=���d�_�����̣`+�Da7��;f��'I�@���D�-���;��*�1��!�E���T�p t�V�b��o���Y�S�ɿݔ�{;��Y:��� ����Ixr�����`~)9�¶'��/�x����w�$���.�	4	�}a�I��L�z��Q��Z�⽄�[�����j�&�$d����(���ا��#ዑ@2�`;>��]�D剱1���B�ؖ�����.�C��: �bf�z����I}�4�ֲ aj*�4��F�������2�Հ�"����bĻ�T�5R�2�[�C�tIg{���7":��>My_?%m�S^��mm���e��R@�֚���������`��4�s�s�x��/_ѽw������/�פ`^R�cR��c����vi��	�f»�M_w��ZW�}xV#�?P�%Q�tX�tI�殟a�:�
��^�'��@��3[4���|�B���3� �ɒ����/�J�.�d� ��%����@�\���ãU�o����Be��s�([_��|��]��5�-��\�L�G��%�!5���N�r52� �_@u Z��i�G�9փ| n�wtsШ�酭w�i\A-�$vh?�|y�zm���l��\�W'`��_Ԫ�B�	?��0ImYե�≫�4&���]gS��SQ3	��ek�]����;�y�gKS�e�����]h�y)�Q;~C�"�/�k���4&��?�ʖ�ʘW�8MQ,�Z���+\���h�ŝ��KB�u( J�3>�e<���S��Yp��XGJid^.�,��&4gg�T�[�9���?
P�zȍ�/]����;B��3`���\�M'Y�r��K�u�*�Ѝ��ڃ�d�6�73��+z��H�C�@�x	/�^p/.G��コ�����$<�X��BP����뗥A���-Vĉ�_��&p�C���hbQI�S���u(#�2�Km1WR�7���Q�J���o�S�?L'܄��y�;m� �k��	7Ț`&%˃��L5��o�zM�ֳ�r2�-��f#�ۤ�z�ʱ��٥���k7��e����8�y/���v3�#�֟��E�od{(�Ҫ4AN�o�֗L���L��Ez�y
eU��l�Ԯ����l�����g���x�4�� ~�`Vs�l	�E�Q�\�mVI�G��Җˮf�Rk	n{�I�d"H�D�Vx�M:��'P����&���(���?r���"�S�U�{b^�z�u<���������j���N�j&�0�d��5+eM4W�E� rY�
��_������F�*#���J�5iA�G������F�5$�S*����,;bM#QFQ����l(���3�M
;l�m-c�T����e�6Ϋ~��t��	X��_��=���o��4t5ZBb�5?��I�bz�����Ur/���Gwֳ\�kd�U���t��m6ȱ��3�X�0.��nT�� O9�#F]<���K�Rr��C�*�@y��@͚oD9{�U '�GF�(�	}���`џT�mL��~;d�y"g�7�N����B����gЏ� ��;`�.�dP����sv`A_�C@�ш_��f�J�2^��]5�9�-��:22q�UH��ok�A[�k�T�W��dْ\g����@����ݰPJ��<��޺Z�0�95FyV�ע����D�4�gT�/���E=�4w��>8�$t���~��C�2�q�O&��/���@F6���~�<��W$�ؚ�ԗ���骲�?TJ���zD%P߯�c���_(ڲAo�'���=nE�v"k��f�	?������kȁ�O��b��hbO�_ug���i�����e* m�2��azۼ�,�����.T�İ
O|�Y��%�I
���Z;���ɨ�R����=d�j�Q[2@y�eh�tA��ҟ�p��z�}�,�i)�Ԗ��M2����*�^���#]}_���~���Fc ����f�-"�ٗ=�x�!� �0�⦗�����ݪY�?͹,�#�39O`S������8�$�{.�(���ga�!�!��5�ay�l�x��RܘF��#�<�	��z ����?��"G=�:�>�� B���嵣4�#�K�f��Sv���D�㈠_�������ӷ-yj��@z�ɨ���Yu���6ݿ���U�;3��.|�^X���bb��ߺ�R�r��Ӝx�cUǮ��VZ*��@�c)��K��M2�^���Y(�x��i.�`Q���c �%I�oc�X�B�m��R��唰��B�K��3�����m�C P��ΦƐ�w7P�@HW �ݐNK_Ș3ׅ\�;Y,�!i�/��}��i��T��>�������>6^ֹC��	1S�.����"��*K^7��^j�i/n̛�w�L���q�j����O�H
�f4/�rB���T��\M$P�̲��=	�j���MPs��מ�YɊ^�ɿ�j�l(�U��K�|��"�r+Z��P�d2�g�Q��$��\�����p{!�k�	��v���R�R֡��­�b�'�
�����$���<�^&��G`�5���Z*�<(-�|��0�[��N�b$c�z�5
XŴ�C>z v�9�����FH��-`����?F�մ�4Q�� �I�����^TIs'��2���-m�/�7����c���˞����h��?g�V�'Z=�����gu��	y\��k�:�ӝh)#5�,kH/)S���?��{^],J�����;��C 		���\KA���l�LWlK�_��U�~�V�*����v���8�gem�nN�����W
���n�UurȒ���X���z�ŧ�C=Ƹ�s@�0�UB5�]�3äߠ�'|[L/Qm��E}����4ґ��N���i�*�7�pKFq�USC�t�߅	k��K���ˊ)����	�C-\��I1���S*}�Y0=EoY��>o�Iᡃ��S�a���We���F��z�#C7��S��T�p�jţ�M)��o��L=��V޼��wɱ�4���F9�St�ثΑ^��mX�=oNpę���+;c֋��H}��6�L_����7�]��]��/v1,S�����TFߨn�>���կSĚ�Ĳ�Rv>y=l��C,������d�)���`����j8,�}\����U�,��!���[kV�%�T��ն�kp��o��B �<c��
A�m}�"��(��c�?�7��|z`��߱!��9O�O�}���Q-����^%C��:���t�	�I��?v̊�������)*�fwN�	(�L�i'���lj��c���c���PL;��o&�����xI���B �f-�]8��.ށ2�b�@5N���,f=����%��B%��lXίg�I�с�=����s�)� |� �R&d�b��1TT��+����N�馬����B��JS9�P�FK!W���A�r1�5_������#�Ϝ�׶e���Պ9�t�㌍�$���eg�D)��B�	H�bz��h2�.:��%W[I�F���p�HUDy�^��"�A��w.X��%���&\�;�+�u�*+zd��>���P8};���!���^�lJ�G�7R��]`[��1#��
�E�L���Yr>��fY<��-�؞�J�y��EGr��ю�tց���{���z�"���
�3!�@T�ـ~���e��倔�k�����gg����uڙ��z߈鋭���,� i+������P�OC���OU����ѓ&��X�%��v�ׁ�ql�^(w�S
5�$��|�-1a߼�o@q��1��TnE�on��@�*=V��c��N��ho�?������gh6��y�t���Y#W'���K��q�B��.<�w�]�q��t�݃4�����f��u��Y9QY�[�췄�����(�z�3��e1 ��#�ƾz�Z������uc�-]�@�I��w+V��V�N="=�f1cq~G�g�8~y��kS���Ӯ_�m��p�&83(o�`���t�|)�J� �[m��Ρ{�d�>�z�/�?NcMx�}�*O�<��k�¶;}A(s�ځ2{�i���oB����Ldn{G��ݼnͱ��|�U,��&�ꐔC�x�ơ���h��:j����(���d_�#D�<�`�R�Ƙ�K�Q$�����0ǟ �-q��4�O�{��K��'�"�q�-eP�U塾��;��ls.%h2���t��+�O�yۓ/ȗ�bM���u�t|���8��B���rH����r�|6���0��՝
���'̾��t�����&`�")>�x���Tit��fow�Ͱ��h �hQ�>������4���w�t$R��$'
#����<鞡]��4���8���:��j�b\
=$3s�6"��9u;�I��V��d��U�*Px�wc��mɈ>A%g%[���i�W*�M���F�����B�̍K
������H�X�T�К�ӽZ6
ިgum_w�����ݐ�fB�j�;j��_�����o�T��۽�U�>��G�%A+0c��[6��u<�(�T�y�hs'�k��9���Iݫ��Fa����&ãņ\3!&��{���n�'�!��\�9���B��i�%!
o.e��f�P�0S3�W*h��	���x�I��C���|�<%��M�l���&���3Nؓ�v����`c�v�p�(+����@	���u�Kv�,���[HʦT��mb!%?�]�Û�����c������2���ep߂=u�.������x�&����Q��-_�hx)p�FL�x���
M--��TkL�ę�mpqD�
�R��^����6����V���iCR5�K�Y�8@77j��P�����fS��0�2Q�$��kh�UfWnC�ho�T�D5�{L��t0آ}v�\Up`Qd�#Cx�#a]X��^�)�����q��A�K�jiL����i��B�ᧃ;��WV�|�~~��\P��ӹ~U�k!���ʲ�Ix^��Q{[���F�uß+�?[����K�֟��f0;����L�s��Y�A����2Ӿo���1n?c(�U/�3�_�.M��FE�k.:��"Z��T�kq��C�nXr��m���pj ��I���=�1"4�]r9S���=!��%VK���'�"H�Ã �7!�`��Sږ�1^H� j ^�%�6���������?9����Nf�4̀��������}�5�\>B��4���-�_�̰L�S[�Ս!���G[h<�y�� CX�<���}5� (�?�w���(`:�ɡ\}��a!��1"���ǣS.�xAt�;C�~��*$֚����
?@_%����s���69BAJ\�1x��@qwe�K�`�[��ݣa8#�+w�XK�m����x�I����;�����©Z��
�e�u�h�@��KIqb��W�ĞYR�����!'�_�H��6�"�W�g(Ư���8��%���Bw�>�{��4G�=��A�2�'6���7!Ϛ��Ù����r]��L@E7Ǘ���Ե�V%�7���^l��T�@m������q�O[9�Q�OAa��vP�C�)M��%��`��C"�1,y�e�s�U�3�_t�i����j�iq�d�v
�߃͖��/�6O��08RW��P[��{�5�t�t��Q�vG�� �a��A��\s���cw�|�x����Éxu�J���2�@�_�1�BeK&So�@(!ӈ&ߙ���G[+�a \��?��O��@�ux��6�~f7�Ϛ'���>6>5����_IzIz�L�f��6��G����B���+K��Z�K�YvF��=(� 1�tk��JA��b?]�i�Sr=�Q|�����e�b��R�����[�y"N��L<�5�VB3f��U�M�o2�j�nc��T)2����B�cB����xs���r�v��������Iϗ>��p��9����"-y�蟸����h?�}o��?w�B�D����צ^Ġ�t���P�#�}�N��!�Gq^�~k�C:-J%|]��`m.�-�8u�톗�������f\{e\>�T1 1�uK�C�&�U�����v���g����C���@�(i�+tl��o{�K���#��r%FP	v��X��	�a���>�k� �5V�\J4��q�E������8.l^��jO���dU��c�fG����.�����f��Ru��d簈S��͆���v���m���(���F9ҹ���K�j�Z��7P��� ��d�����m���f�o�e�������?�}T�G�m}Z�m-�(���/cg7�zc?������T��4(;�E�'�Q�)L�|L�@���q�H�[�p-,�v��T�VR��4Ӫ3I����|�9B��B@�/N�����0*2\�v�?B�����ԓy�+�]=j��gyf���\��t����k�N̐K)J~:�ʀHHE���5|�HH8��_���~U�)}�o�������ˈP麫F�Q��!p�#ǿ�NXs���f���ROJ�Q�4"����1�4�"�{����S��䅝����_R����@�l2�� m׸Y1^��AP�� N5~�/��C���%x`����qN����Q�c �O��({�W�)�\�\Ff��&(�{x�0]1���m�dJ�f(����fK��"�n��$�J*�T*���yr?捺��0\RyQ�Ys�t-���փ���3�����7�M�DB�d�s�U��(-��e���J
�����k&P�~�5��g9@�y��D܁Q$��E����0�BӾ�@���ᵐ���z`���ѧ�?�'�7uu���3���|��b��-��Vk��2�k�L�+P�3�nă��몮�kt5p�I�a�#lGGf� C���Ť� ���f�����s��[	�G?�p%��#�"�����m|i�-�zb���s�}8�[ܮ���5Y��G�6-�V�-h�O��/��aY5m�N��B�f�1B*�o�\�ڮ�c��K��b^o<��lc�uQ�c7�8��������;4��D��Jw��^��	���\���d�7����>�n"fxK��.F�s���(�#�� ��g�\n	A�U�kp*y��N	&%���7�0�*�]O���\�`����XX%�M�`��^F�Y�]�Ճ��m�`�>�NH����*�:|u�)��ru'�.F��N���^�����!�$l`dyx�p�����?"֫L���ԷP`��'����C��h$������j'n2��$��0Y~:��^��g�Q�����/e7_��E�]a�-@.��afR^V�!1�%Eb�K�Eڰ�RN��*c���F�gk�<3�<韒ϷcyJ��"%�\~���V��[@���B3�h�{���;�/אo{� �����K+cY�͸Mz${��Z��|%��U�|G�U�bw<����q4�_C0�Wt��]	�*-���7P�<���6AQH~h��w��x���-�Ցy՞�e��5�3��8�}�-ܦ"Խ��qV�_��/���a��*��6�F�_> #mV�댶tt�����F�JAx�l���vɖe����P�]���`V2Z��5�>�OM�!lᵾ+��@1�*��VoY����:��Z��D,�S���V
��b�:?���	>yg�/9lo�X)�[L`�T}�,j���F\�X4�yU�X��=�+������AX��&$���ꥫ�,���kH����~Q}
�p�5''c��B̬b�wR;�3p�ΐM���.�؍��.�	��o�U����g&oͲ�-���G�\J��3��JNMP\�_n& j@ɑ5Q�����t�\m1��͙\w�9v���JS���1vb3���-���c���4c S���M.��B�fY�����!��ǧ�冷��3Y �M=���`y��N���v�[Ա���NI/<>@`���v�	��J��}c��C[׺K��3��r��F�.�M���k!�W�vw�	d4����V�#���:����O���ɜk¦r���(�W�(s�p��m�
A&�P��U~'�	9R���W��tho[s��Ȋ�v 6P��t���ܷ�؀e��X0�>�=���.�Ұ�ͦxkJilL.����DP��MW?_���;V�:g�9~L��ru�����Qd����i%��:���\	�
r��#����ԏ���3�grLQ�K��vpn|zN>�Zy`#`���G�G~!�Ej��*�+4&����OK��������G�� 
�Q�rQ���?):Y�ݬ}�]�1"�Ύ`:�a���D��5ԅ\�Z�.�5�@�G��h'��eyO3�E���->���!9��` �5��� ����v��RX�Ɍ��j�vW/�����;�p�I����)4�n\\};j���\xG�S���;�2j���/�<��B�b`���҉�_��������[��Ҫ~�+ߝY	�x�C��,r<�s�6��)Y�&�7��!1�ZM-�[7-�̏i�)�{��8���I�$�V+_O���n�7:��ʁ�h!r	�7��th�iH�'�O��S�&5UA��Xo�{�,`��Px�ΰ�\�j��H�r���߫�OU�$�Y-x�q��1��LĤ�?3f���[3-��0V7�P�������u�f6{��A�HP˼�Z����N��Ǽ� ]��$Tr��;eD1����C\��X��ʘH��q���Դ�a���2�\=9cw���u`ﱢ V��3����N@uٯj3u5�3��X���o��7v�Xvo\����5T�}����}ʊ�B��c��@�f0���4߿���E�g�>ݙ������u�4���;�"/��^���ľY�	��Z����n �gWY���V���.��[;��Y:H{,Sq3?�ul&\-y�݂�D9��p�g�؄���Q��zz�i������m�4=`�d��LL�#xA2�O�
|+ܯ��}ĊRb�����G�����FU_X.�KY2/U��Rk��)�#��\���'z�2u�'-�,�!�4��P� J����p��L�z�Pzo�C�I����>ic��{8�~�;RW�9�x��[,I� �ƶ�J���L�;��2m���ޱ�=/n��8[��3|�}���hIP��}g���vS�)|%L��c�$M
�0QF�2B߰Xu�֗���|��W�� <���oO�c���@Q�b�s~mِ�¬��� ���i]X7���Cu���2�{��yHuVU���~xd�=����-� �=��sxf�0�����*�U+������rҿ�hm��u�N�npń�/�/$���nSӭD{����3C��������H%���95?5^�����"�*��Tu���y�h�e�=�8^�-�v��b�"|:�IZ&_>� �z	��\7�%6@��EH�7����P���k�֥�SdOK��Ei��mw��%��u4]�/�=iB�xޒ�;t6B����]j�2��8����:j��Ay��]zh� �<�s[�6�f\����o۔�	����j�??@�Y"��������Ko~����1ݢv�kЩKV��h�]N����X�5 ��� ���@��_��_ѺÆ䏍ub;�N:#��j#�6��ey�>/}7��Pv���i�_�\���q��?�x����/�s�-َ�ۦ�E|����M����ϑ|�瞁��Cs"�6�X���R�w7�h����l�0\^��N]�0)�����kF���aSJa�V���D�lR���	�ę��Ջ�Դ���|�K�e�J�E��<����'���05�虚>dd:<@0:�#��M�Ҧ��ym�j���|��4��=�Pc� ������b��SZ���Q����f3P��K0�WB�.��.{;�A�M>\g�j�ɸO���u���1^B+L��ctr�^=rh1Ӓ�M
a#�$���vQ�s��eIg�漻!y�{��Y��N��*��#5���DN��N~Iz?`�V��0�Gp*`�+�JK]G��-b���>о�k*�2�ĸ����O�,$Ȓjm�_GI�����q�����R��l�^��{�
�s�Dh�8=�?��$��s��g[y'�W���^�F����=P��$�ϥ�}w��av����>�a؜�D�� g�a�6WBݜ�|h�=)�+yF"TΜ2�o̦(!ߗ��rp@�Аi�>ΰ�����aQ������M���T���>Ը���)p��pL���Nu�Ĝ�qe��e-�AV-���[�/n\B�����cr���=���}���*�Lۄ���
B��V�ȼ�T�J�܇[����~cu�Zy �@b��[����B��o���.�t;�{.6�˓��x凂�eI�2�i�-�W�f�׌������>�c���{����YrDA�~�f�S��D;���i4���n[*����Yޣ0<Ҟ��?j4��kb/��?��pG���\�U��5�W�^
{��'op�-Y�Y� ]�9L1  ������"D����x���_��U�lI�<I"�����¸��р�>�l�'�3;��� ��%�hR;pv���Ї� �Va�ݴ3a�>ޛ�����\^�����F�:���J�͠�p_���U�O���zzQޡ�͙Tb�'R�j�]Ʉ�Tʥ6nߕ~%�Cp��}�D!���V!�����D�N\Û=Ҍ�_=1�%��/�7�69��
^�5qa���~ˢ����[N���/�Z���	H�{�Sך��FF�'�(_!�r�W�V��G�6�V�	A�-�X54�pKY���_�/���J�r�y3���̽?"��H�?Ý�\�����s��1�7�M��IP:�
���dE���_��.2U}d����q>�ˋ�`��z^z�������0Yvݜ47Q҅�F������7��7��'<��z�L����E>ykO\���T׉���Lի�L��8Ć�Hs�};�T`��D�H�0��@����-/��W��P;�8��������*-�%�IO��%�ČT�!f����A��J���%��br��e�a_����g�r���a����)̍�2.(.3�3�;�mNѾQ6Ӣ�|*lČ�[$ѷ`��9K�L�)�#	�Ž(���_�/B��)�R� Ҁ�dF��?ԏP��@7�(Ja�D��f�Ym����<���@�ǲ�`���O��)D��c|���N̩�+x�m�? �����q���VW3��:�/+�/�N����5[�u;�����$4������Y����șuK`|}1�=��K՚n�35L!(D�vv~��8�ԍ�%��W+#�CᎣ�m/�afI�r�Mx�k�y�x�~c1s���i�J�*���a�8��foź�l��%�S���h��
{#��]	Q��W�"jׁ��X�v�ӿ۔3퍆��B(s�_]�̺��~�<S��>�i{����
�P�,G����B�8�R9��[��B�w"�����|n�c�Ir�GS%�����7�3���]xnXD}�q���f���ײޣ���ߒ��d�!P��B���$�-U���W�9(��ȸ$���C�fr����Ld�M���^�F���k����nS�3���g`�����۩w���E���S
�EH�o�o/�>�/T5�����
!7/�QG��n��dH�<�͌wC�uS/���3R���B�ܡ��My��w�T� I�\�ӌ���IG�9�e���h� �E�؋�S��kJX�X�����я��FJ}P�<�LmJ�?Kew�  47���n
u��?�!Cޱ Kĕ��z���_i���\\��uwm��I9�ycW���4y�ƭ�.\���b�O�Gi�����2��bk
,�!O��E���j�����:�V�̻iⒷ�U2q2=PU����)�֌[�UĂ8��4�"�`���%��l�֓�v�+�y���&�#�����phZ�I�5��.-26Vb�C�}/�*����XWWpwRs���������<�E�����!M���&:�W�f
#8|}Gڞ������HT�Z.��%���l�4E��p��$!��ă�M_��Cw5��S���V�hh�<���Va�o�<�K�;vq������Z��ô���+az��o��
YQSIx��o;ɆE��$ܣ&=Çah����
D����p|F)�}�=v���ӈx�+i[^�����d�V�M4k�:n$ yM�v�k%�Ċ�U��&�h�Q�j�����-|\_���*�Ar�u|��6�$kT2�A�/ժtz��Pr��ݗv�M��E�c�sY<4��c#\N��摇��_q�#�{P]��_������|�K����6n�.��o�5�0?�4.0&��bLA��g����tS���;�K��t[\kj��U��@��R�{W�}�;H�9D��������$ޒ���s�����l�����@Y�X��j�6��N@DL`�M�"�i�X�L���9��[�:l�h3�#Kf�z�ք�kC ��nA����̯��LI%?%x�VI�����y 3���Y�G����f��+�*����B!ʸ���NO�&lT�~�`$�_�9U�^聗����"8�ZU�����5S�C�ݙ%���$�ހ�M�S�(����)X��܇�Ur��*��]���{\ԵD.�Q_�9z�c��Jjf<q/�ZY�
�e�Vz�y�Jb�����ƒV��T_�AL44���\��΂�K�Ua؅�����؊{dl��\Z9;%���{`.�؍^ں�$�� 󢣃(�J-�pXΙ_�Q�9w�c�=
�l� Ф�N�3�m�����r�����W������Au��}�n�>2�����}�.���ҁbx�O�<�L��&t��9,��	�U�[�DuSHvV�K�+��!���)S������� ؛���	�m*4�9�&�V1��!^���� `��hid�ɞ����ue�`�)݄�ۅQ��j+
0�,�]Ga�m�;g�r%�,j�]nN�`��S��jC.�����E�.�_�0�tx�Z�ߧ8E
	-�C/����c������gO�_\9�P~4��HP�5��Ō4ƈp�4�K#���O}a� 4vA/<��U�HY�R �^nJ7��ڤ=�t:��Y�X�O�[?L0�9D�
�}���4���p�;���<��7K/�ϦW�U���%v�fl�֨��stde!x��ԁ�\/��y����DL���S�c��;
����	�D����\��$�;òj`(���[]��gG+:��JGS"O�Ob�fG���,0)R�����~�"PEwUyR���s^S>��g��BC}k���/��_V`�nq��;�
Yi�s��.�v������	��-�N�
0��kh�����P�����go������tϺbn� ���m��QH���5���/<�*�JL�%?�	��mri�et�l΄X���N�5����\�����ɕT���_�J�g��7D��]%zL�����i�/��УS|G��ޖ��lE�O�H2zS�T�����3ߓ�o����c �]��Y�/m�Vh����b73o]ґ1�$RM;Ŕ@r���{�p�p�`H��#�)�T�Irw�,AH���@o)rk8��Ns�p�' =��Ź]}�����K#��y��bN=D̓DP;`X��SvӢ���#����bL=A�Tr������������c����a�M� \E���q�J+�g�ʣ�t�P�����R�L��ZcI
7����4�/5Z�xiCS�0H����248��@�븃 �g����Si�l�K�^U��}�>�$�����/����!����i���ED'(� �F�=��7�����w.�^����X�v�]}��\�?����e������O����B��"�p�C��8u)7z*s�Y�u�Q��/��S�,6`�h����T���C{!�Ho\$ͅ��n��l��b���\�sGO�.,��V	/�嘁�L����'�ڪ�].�O��7�,�BI�Bj;л>�C������1��S�����2-1d?���{��㞨�K�`"�������6�����6_�i2nWY��;Ie~��x�+)�.$����j���隐�$�p�7��/K���3��Ka�2�َ��M�>e^;0XM���@�¯^�ԡ����ߏN;��q3��q����!kѳA����Ҫ:D�s�*{kn����FZ�3�+59y�ˎi�y��>m7����,*�.��Z��3��\&�8G��VR�[W��ӡ�ֻ�-�=!����G�@��Au�	�R���j�D$)���ED�G�F��*�?��U'p�����Π���ivh��b��W�𕅉�6�䘐�i� �e���ʛ�r���mc`��d����2Y��q�薝�t���|7�֖C��J�9�ם��|*�Q
�M���@z���ho�����pC��kh�^�5Y����ޣ�k��@����|u