��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�R/zr�!�����-�k�w��gB�i,��==�զ��+�)q���G�]�p7j���)x�0���Y���9p��29
�a�ΐKo�m\�_*��5���� ����	?�A��S��U�(-�ߢC�ܗ�>F]n������5����?���n����I+Ii���su��E�6��i��u��-Q9��I�� ��!�B�|���������Y�,+�cN~��A����f!�r���l=
�|��Ҋ�X�Ɨ��͉��Un�qe4��\2�s�T"g7���}�Q^�������#���h�[f։�LԄ���-`��7����0��Rm�@&�-̉�Y5�ȵ�������D^����h��v;ئ���݉�m�E����A�.���S��rO꾬f	�� }�4��&w�x���{�7%rQ��=��'p1���hs�/����f�w>�?��K���Ww�>�����QT4ZT��۫1�̕s�V�?�uϢ�h ��+)��o%aS̈́$W	������U+���r1��)}�KڗA��L�e鼉�����k��	9��{+��
[���- ���Th��52�N˶K��-��ҲK�`0i�������+�_�;��E�3�L�?�@�6�܅�=�!T�d��z�@�xҷ��@���;&u^ֵr(%��3��U'���LF�'��vM슟�#��y�p	2�����1�w'�f\h�	�+2��ͳ�|<	�o'[`@�~�*:@:�����ڃ��-L>����;���靾�Oa��n��0mL�;�VS�W`J�e�r.�f��qL��D]��A�E0��)<�S��3/j.>E#��3��FH�/A.2/�"��2��-�Ь���K.se	��	DⶥU�츳?D��c�|�(��D������:5f��H6|���4����[�ʉ��*��ف����S"~�M�.6����b�G����'4�	sf"t�d~�_"9�1�����?F|��g�+�`���q������)��a��d�n�{[~����_���8���e�[�?Lq"5M��K�%��PiV�����Y�}7K���Jop�9�HW-(���[��90dט<��7n�~�i>](�)Ş��9����%a��8��D[X���Q�l�(��Ya�6�y6�;�"�
�QS\A�=���hոaf5�c��G���LE�2E�po�7�b�PТ��nه��ɭНO����<G�e����'�ŤI,غ���j6�@���p�rH�|[����>{��|Z������3�L�v���{��Ɛk���P��[T�m΍��B��wPj��[��"�5����l��7�����$ɨ"�m,�EhJ�~�Ϻv�!������p�um�`$S�<��ࠧ�_5(�4,jw���̴���u"C×�b���9OVw��DD���
s �zK�#O��@o���0�69��s@�nt�?T�N�=�� ��������Bx�NH��lb���sƛ�UA�G[$���mt��*�_�#t�auI�+mwJW�IivN[3�$\@߽oS�3$z���n�WF��%9����������;j������5�Θ"�t-T*���j��>7mꂙ����� �'� �S4�HX�$ӧ�9"�FC�����%���LpRn���D	+�ıy�%9��P����. �!T9/7+���1gK%��h����F���vs��2�.�c����J�/��W"�;�|�t�]|1B��L9{�q_K&#n�L�k-�$|���H�����v�b��"�x�q?Ɯ&���#Y>�GQ�H�g3��m>D�Պ�x���6�v��T�H�l����̬)S���}����fOH��м���\�!������q�  �b����������NƼ����-� ;Va��������,%!w��^D�aJ��-'�J�b*��W�8Yf�u3�����p�8����	XVЯ��v��]l�"Xt.��!�0�Oᡌq�l�@�o&V�
�W��97�Rwk6W��D�|���@�~9ο�ٕ��h�\���ɬ=��b	B��7�1傐�,��ؘ�%X�B Z�n��E^�@I)��'� )��k�!���b�\�1_��]&�t���Y�.D��+�`3�\}���η�1�٫]!����]��g����ګ���@?��3)ʂ�r��a���neN7��,`|B^�	���+- ܪev꾽7���o��*��HJ���m��Ifd	�EA R����ф���	�H=���4&�Lux��i�����}*�=��@΂M��Q����Z��Y$�^|�)J�yC���j7�{/	+
��j��(�h��d���ͮ�6�ԍ�&����t�43΁T}=���Ɲ����UR�'�FƯ��?7s��>p����c�n�H'���3�'{d�����(y�J�Ϛn�4�}����|H�_
���@�]5�L�T0�:"�Wu�]���%.�.*\W��w����Ơit��c4�K�{�����:�@��������������no��̸*>�����.E\��OK���E�.2������E���K�)#.�"<M��ª�jY�I-�,'�1a�Ux�f���ԯ��������x��ĹS�����24�t������SS�Ri��Q���:��h��ߎ�ʈ��>�J�iOr1C�~?7Iڄ�E�'����{��\�K�"����X�Pp�Z���_���x���}�^wyZ���e�d�Z�
[�rV�%T���g����V8���%����6)%ނ���x�c�ޢ"X�8�D1L��7�'��3�Kf\jF����s%&�$��rۢZ� �0���n�����j���F3F^0r{�h4���a ��$j�
Pu)t�.�'����5�3<3�mP�!��ݻUo� <��o�h�;E��"�|+�gdw5s.�������݌ �B��|�]Y0t�>+�W�sR&pG<Z�f�x*G�ύ��ej�6�I3y�]Yu�<�|�ATw�����w��S���̓:������@d���t�� fO?�WN����'���u���׺K�!']O�vI[P�Zu#�Vټ���9�3)(.�Zm�4¥L)���%@����zd�,��Ӧ� T����.o�^$f�P�m�f�7	<�`kړ�JM˫k}��R�ٺ��J)���+1`��ـM���X��{�'8[�Amn����)�ՑΜ&�&�n��\���f 3���śa6��?��>�� ��p����Y�w-JrW~�K��A�o�����3��VO"U�n��_��e�=z|7��k쐀��c7e	[��:��-�}�q_z�R*nr�D:��q^�>΢�m!R�Й�%A���^w�-��?a�b)xy(��~ϩ�L���֧Ò�zdT��k^\�[a��u��Io}��mӿ`���d�4��2a�� .��&�9.hLb�p!�˹bm�s���I{��W��DI��R4���o��ia��ͮ�y2��H��K0bC��O�X> �@�'�9h�ꬍ��[2w34r�� �ÖsAhЁ���y��&D゚�#v~�=/��>?�B��������d5���5J9o��0~�;ܴ����'���HQ��.�ȸ�W��"�l�����~O�}Bk�̓���J1�Rt&t,va(uˢ�/����� �&Ö�k�|r~�lb.Q�(��l_�˚Xۆ�al	�}n���v���@�\S%�FaQ��Цx�S����;�C�b�$ĝ.��!��E�?u&u�m�����cp��9�^�&���_d|Ve 3~%$���]���s�l��ކ�(��֍�f���x�x�.�4������!���YS�ԃI�n�J�D=�I�8)�뢇��Bc� ���ș@�j�v�J�Х�.����'��uC��V��;;a�=��b0�4���,ry���n���9E�%�و"ӡ�R�<Mml�C����i2K�a��P���o`�H�]���W\&V�~7���ۊ���^���{�Z<�U}pE�I������=�4��Jo�r2v��x�J�C7�t#]�~� |������sc��VC�����?���(`��ANv�଼�9��x�P=_�fF_�z����Bl�5�S��>e�F���OwzD����w�}���v%	a��8*ms��B�l�ˠ�TM��b؋��7Ht���71Ke��ڎ����.��PL;�^�i��$�lڞ&������Uu��p*Gۻᄈ'���u\=����I���b`�6Ycｘ�L57�>�"��,�#V4� ǔ��V���ԯ�C��s��4��h�_��ج���R�{�wK�Ҥh���/1p�qs���C	�b��ŏ,�\�<V�k9���D�'GoP�?��	��������v���R�oO*��+"�h�{lʅ˵�~�V�����^�O��]���	������
���vJ�,���r9_�.��:�}�o֦
���%�ɋ���=�,#�n���|�7~@'��h�sp��sD1X|4�8+�6������bj�<��!<u�<z1��4����jU��[�&vTS�Y��(F
T���k&��}|�� :E7<s���̻���.��d��-�!�x4?��V���7
Ƴ_@�
�5(��dG˛�?�;����B�o��a��W��ݸ��V�N���Ⱦ�ͣR�^�PI��i�g�W�E�E했_|��>��0���'��#ª�� $:��� 3
�@�W��4z�Xk�Ƒ���)[_yyHk�ň
��
*��1��
��>ek����
9;
�A�ц�<`�UB�9�oT����#��`_�ԨB]F^�pK���cч���,̥�F���>T��?	�����80ǌ��Ƞm&���ԧ���'	%	���KGC|��'�7iMkӜ����I�mJc�Pc��AC�&��"t�?@���>
�f��\�]�W��R��e�d��CE��$�����'Νp���"��=�TYT�R�%7�26K��2H�T�T���C�V����sd�/����z|H�(�,�K�.;O�@Y��^E�<����?���*��"-9X}bޒIw\��ܦ�f��; sdʺ��3��L�����WZ�ҝ�j]6�KS�9����mr�������i ��`���d��%e����2�kвf
z����df�hŇ��h�y��!���s`'+�2�j]���wP�u9B �	[�y���-��� �5flBƽ�Ya}�tb�ӱU&�ڒ�1��eh��A0�/� ��>y��mr݅���*�}�/�+��n�+��� �����RM��*��q|~
Tޅ�&&>G�6������_���M�;�d, +� jͨEm�DV���D,���C+W7��u�W|��RWĚ��,�۶������o�!�<�/��x~���q�e�Ґ�������x�b\\/�� �0�S���w\Y�9^� �=(��ѫޓ��jE�o-�~D'_��� +7S-BI�8oj� ��*Y���A���uC���k4V�@�Κ(Ý_6缿I*><�D�ǂ����6�xy�\��3)>D���7�}�f��N�� >ڂ1^9U��aq�� ���\JL��*�B�ZA?��/dS�Er�ki�ϩ��] V�B~�ܨ�sL	�/�ä́��)�T���rU���#�i� )�{���8���@ Uzm����a=#�t1��e��Y����g�4�µ;�2����p �H�}C���x9�v����9�s!��c�"��'i<�vp�jxQ��3�/�ߠ��W�������t�-��:�[�YB����O�U��%a�67;��