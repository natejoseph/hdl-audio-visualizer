��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]fۧ�Ɉ�A�x��6�]yJ�����L%�J���,�c(�60�g�]�t�Z^�1p�9E��B~��-��=s��{�����l�u^I�z7���h��O�:���G���R���a�d���ѱ�p$�S�)�⦺&f�C��0���R�=;�l K���� dC���"�7qyG-�(��n�|A>�%�i�����:����y#���%{p�Q�I'���YB�c�D,DRf�Wx��8m�W��2!,�_n�S�����{��um�����U��c댋�$��"�&�q���e� 1R��?�4�K���N��$��[���7����h(�ܷ#��H{���4���v��GW��G�ṿT,)(���:\w���2�	�t��D�H��Ru/K�3��x>_z|@w�d�<#Q`_N� F�n��.7��U�p������{�i��E)wZ�"so��~��g�lM	:�uA>���"X>
ͮ��PO��&��]&9�V4�+��d�.	�ʂ���ؙR�[�d���݁L�-�P<��bIEeM"�o�ݢ39؞Q�^�y�'w�fǽ��A��O+�lģ��d�0�}8�8Wp_;n�ĦOO�~�5�b1���riSu��\9�k��`�7�ղu�VǕ/�-(
���6���;��.��.����dM���ڧ2�pH�����ZӚU_�(�7�eے} �I7�'@�ͱn]�Ui���m���Ǌ��) ����?">��ӄl
)�2�͏ՠ�q,+��]?8JL��h�j YG�'|����t4t%�h��s��3Ĳ3	k��]ţ���Q� <�Y@x�̓x���o|�`6 �����G���D�O������h;�r����I��F�/�� ������U���Ȥ�.��[�bӤos#��|�	���������$�JnF�A�ӓ�7L��;��o)��ᕕ�:I��Y�-kx��Qy���E��hʞ��u�c�l��wk�\u���!��T�I�wל��i�v��a��	�7�(����Hpm����b@>�9��T�w_�|4�b�*�b�zو�B'X~����:�-���^HUW޺cщ U��=�=���Y�z(�L%��ݏ
�ڰo΋��v���3��!� &ُ7&?�I��%GECAK��6;�R`�Ot�S�]�So���p#7 �a%R�Tu	q ��V���j�?a����\�u�`l�H|h�AՄc6��ٞ�r�r<�"��t���0��9�'�EB�ۍ �>LlR��/ ����V�}vu��,=V��	/�(k�!�#����Z���V����˰@�)/
����A����[!�,HŐ�Hܖ	�A7<I����zU�tRI�);"�+|\�F��9&W��� �a91&��<b�8�����>X˪�#�d����W���
����ā�>�[稄��.:��Oq��s��=�AMM�9�F���=	 "H���W�2>6���x�M����Z�ؐ?��RM�\����� ġ���n�3LK��TZS=4��!ό�J�F�Jws�pv�6�z�	������F�e���:ο�Q�GN��U��6�ެ|������S����=P؛�����C(�MŹ�7�Jq� �/�^DBa;;���#�/%�T
c�#x�nԘ+ߓQ�W?�s7��UU�|�>%5��0!Wݝ]:{�)$P	�msZ"8[V��8Y��q�EA�4�R>�=�d5����N�C/�H�����ef"�.���/`�?��(x�>n��
��pp�3��~�-�D���CrTU9l
�?��=�n8=���U�`:������!�!���+����MKA�a�>�K��{6��@�ǟŴ����qh���\}��IG*8K��9�dP�A`́X�eO/C΍I�K\�a��ʭ��^���k��&K�
�J-�8��J�\y;�{C�#�#l@�i�bq}��~*j�5�'��W]�?�8��M�^�ޢ��G�o�U,K����hJX�3S�^�htT�V�TE�1W�e-!�s���B�e��7����!3��o�
=���.⟆��>�]k�b�x����5��,�~�F��d�U
��T(`�]��Jh��������=���5���I��pvc_������/P�_���)o��d�(,�˪�q��>p�E�!Պ�SUn�%cp�O�^E$I��}X8�m�rF�G�fs	��[RT�@;�AB����c�r1�6��|a���?���At���� "�_�!�5�����IN��6��|����s=n���8_	)7'�qd\�H(c)��E~`�>JWG�>T�Yu�D����EO��א	���'��v�ŬU�͊�	���m��W��<�g��EZ���1���+ۙT�:�iw� О%Ɗ����c�0�Z
����I�Pv��AQ~k{�(b�P��~�A��=��8�l!riE�8ⴸ�,�Y������ԣ(Z��������]0{qق#�t��1�$4I�2w�[��Ej'Yj��7EՎ�_�D�w޲�D��=tg�/&9���Ҭ�p�~spR�����Nܜa��2��3ӹJ��㏒~�J��#�K�i3�`��Q]QRs�����x�V��
��w�3�B�@��H	�����7�OY���)9KԷ�\7BbNMr��,�D��C/�������\�ÏjB�+&��b%��qXrk��`}�I��Ż�������tSh��Ȳ-g���mf�5ӹ��@L�q���Rh<���}R�����RA0�N�Y�ӊd�����gt�.�`�w��JuGt�# �ڞؓ:SB��-i�݊�g�}��"�	��qE/Y�M�²w��BB{�����Avj�֜yws�(�<�0*\ej��TN.v�X�琏�1���ث	��Ӄj$��xN��'��+,^��y?��Ch��b�,ʝ`��s��P"������C�+Ľ΋�#X�e��J�1���cqu�ŮI͇p�{��c�]�)��`G�� :���(/wL, �p2^���K�l���5`�0I X�'�����b�8��uӭٙѥ�!l�ToE�N\���鸃y9J��ڀ�N��\�?�^M�~@ּ�*�#�j����%�L�6މ �\w�7U���Ţ�*H�W�����8ەg#�<Ê���N*flZ?/�a�����U'ֱi՛�7Q��_|�U��?ykҵi��]p��묘<� ��%,y�)�vH�L���b' ��ɿ����Q��c'T�C�$�@��K��i�2�q�G"��I4����^_��3�QK/�^�CT�����>4;7S���g�Y�B�u纈k��A-s�䉾�!m�cnA��,v���;?��ܷ*ܹ��eЃSzas���|b�7��9��d�ӯ�c�$՝퉏FZ�5����F�rl7��搭C��tX�ι�:|�/ FI^}�`���箶{[�c��ٖ&E��
��6d�������~����B�K�;c��4Y�� VS���핫?ʊ���A�k�����E��r���;E��3Y8����ON����GLŧT��h�m岅�VV��j]v�K�ƛ��\��Z?LtB7��x�8ܱ�Z��ݘ-]�&�v�Qy��(.� OJ�D�ў2��3��@`
��S���a�sxL�A��ҵ[�3=������[�o�4[Xtf�@*U�;�Տ3��6.�,G+^�f�<�Ab���m��$��]���!�@sdyб^hW�/Xu�t��n8�!H�71�K��P�ʣ����s�Sf0�2l������8��U%�r��2�]|f�	 U&7��,|`�+a�cH0r��N��G;S�_i����Ν��^���:��(��^E�s	�!���*E��Q���pD=�砾hjk��s����F�ͅ(+�@��7CK�r[�	x�y�^fC��?�!�
!�*%��MޅH�<�@I�=m� <P>!���h$���үY��͹[
;c���& �{=^���,Pa�p}h��5������ H���g�yɊ>ٷ����h������:U�8ѹE�E�UE�Bg�k��uU�i8�jX��Md�t����+��;e�<���_o<�"�1Ƒ�N�":ed�uaM�� � ,Q�/�/��<�����& &���y�}��
�e���E�=Kb����B
�\X�q�u���qR+���!ˢ֯H�=��m�i3mܩ�t*d�Q��6�{���fc�\��d�.���0�D/d�<�T�唣��&_[�t� J�Ϯ��_O�P:Z8D{�F�s��1���n�� ���(����>��{3��%�]�08�;sD�;4�3l�8�ǫcy i�E�J<�X�l����^F��DH<�r��b�l%h�����
���aaO���%�	��R.�P�u䚓����ܤ����Aq���Ii���\�e�2!<�ц$-0���� ��P�{�Cщ���n]Xw�֥`r$s ����ݽ�Mb ����e�� 2_vO�� �vp�x/��O���,G��B(Bp������#�)�X�@ۤ��M�m��s�H�Z;�,�1���sѦ-�A�:�|��K��|0�+��Q=�d	��5��u��=&��(^�$��Ug��= c�����$(�����0M��`��.c�g���t7�c5eV����H�5_
�m�	B~���Q�a���dd2����V�d��?��-��6G�#$��!v{���<��`���#O�Ⴖ�n���'U��8�~s�{UZ{�B����A��ߙ3L2�b�_O���\�N0�W�lt���9�Ӹ��}��p�n��O�����U��>�a����&LWY-�X���J�����[Z�x��Wv��΁� C�YI�&n8-���wr�=��;����H;�����壏�z0�=]����r��hx����w(����a"Q�P,��_���^�o���'=�D�e"�t�~[����Du�ymH-鲃T#ފ2�!M��uS���H�m��\��5�x�����*���aﲝ����j��+=��ҭN���~���WX0f
�#����߭�M�U�V�	�S�f�w_���9_דG�J�-hV'u��?Cd{�$���ԡ�)_����Q3~c��K�ު��m�}U��-g=����;0�`�b��&�v���>�?��g�����#�ns�z��XHO��L?ޢ���.���ʃŷ@��lV��~7�?��t��)y�6#�kot<��^��6F<��ݏ���뱅0���%o�U��'��#ȯ\M���!��%|�+�ͧ���)�/�*��xC��E?ꟛ�%��b�����(���J�ˁ&�������ʿ{���R�='�%]�p�Ӂ��(����=��#|��]z�q�F[�QY��0r�E�Z?�U��ըR��璎3��
��6�
��f�^f"+�@�7��8Q�,��#)�3[���3�mW6�!����w/V�Ǌ�~�卶%@Z��PwwX�kٔ���	ƚ�#ư&�D�xHmy�AK#IЗ�}�`��]��� ���Q��NX�@惣&<�wq0����fLgm/$]X,���Z�e}Њt+�-�87`��_<+y�!`G�@��p���^�I+�[���(�������jM��&FB�%+���)j�0e�*����N��#m��T�+�/��WomE���6���L�)r��$m��<�۳&E��Գ�%�Q3aǱv�x,5������Y�KXq������S/�Qf�����-����LJP�h�h�l���MG���PZ⅙��z��L���G�t2�꽂"5#��~M���Y\c����@��;�̯�
�Π���%SD�*X�k����h�XB8)e��5�*�K�]-�_M4��J���X Se�%ϳ,��3��	J�Y<`�4X�1��0�O�iD9��H9[ 1�&�r[�t���;�|�Du��~����0�0�$(�@� T��Ǌ��6���uI�컪�����(�9̹�,�W�iՃߊ/�������0B��k0;[�����Df����d�au���V+��T��� G9�� �,F�fH�*��^V��L(�P��N���E�!�a	�P�2���:��d�v�"9��J�A�iFC�}���[���+��	�2GS�!�ڋ��ou�(fW/goe�]/ju��U���m�ҧ�x`m����������#gT�Ⱦ����HDc��ƤN�L�wz�&i���Z�w&_zl����lR~�!��3�.B'Q:��|�$ANO��:�]������_]nGs`�X��&�l��#�˞=�\�yyJA0�_XU-�'����3�e�Jm�P�q@�f�$�Tc*���ȕ�4���ӟ,:��ʜ[������^p~C�,�t�@Q�%�~�B�jІԲ8GE�k�] Z?���5�g�%ܕ��ͤn��k�)�DI"��H�U�	ͻ��fZ2[b\�F���#���"O>h����K��K]��DgƆ��&c"	O�������0��؎V�U�W]JD�j�]���g���5��PӺ26����|Hi^	q&�!U}��N�c�
Mm͝i��y���Ģ$�0;���	�VRogPܼ�+~��dYGR��m�3��$6�t�64+OB����R`0�IR\�y9`y�Ɠs� �bϠc��� ���{�����÷�$�2���_v�l'�P%9ˊ��2�����B�=�v��Dg+��+X��7%�8{�� 2t2�����e/w�JR2_�=j����J�CET���{�+xnh����K>���(�����}e�E,=�֏7�S��ݥ�7 ;�L��Q�ŉ�qȣ���������4�`�Ɋq�{Ҳ�#��)����Z�n�Z���������y��[��Զ~
܎�3ϥ�%(�,]��si��̙��b��)~���ך���50��A�,�p�5O�q���R�Ds�44�o<��>	f
=|ӏ
���/ �tr6~C����F��a�C	@�a{�0{�����+��\�'S2u�I\
@u��8j���V����8���,۰r�A��F��
���
�Z��e�`��\J�e2�F3W��x��t�X0dP�
��K*���1��t�{��� `�����(�Q�{ï������_I؃����U�b���%�����nѣ8jn�Ϛ�z ��8Cj��
zҠ�j�>���B0�=���[O_L���Q��/֮�U9�\�Bf*��[#�g���&>��/؃^M��^�\�Y��F���)��a~<\��x���-�h���N�7h{ߎ�����B7#9%7m���GO�!����qU:Q*me$�s��4$��������ٯ��Pn�s�{x��e2.�5P9�6E��1f����h�Ԉ�t!������.|� �gQB}��:dͺ�m	��\=�c$�#����+&�μ�7���AU����Gsk!�0{��c�����[��m���e�K�v@�3���N\N�Ӓ�J��v���#���Mìȩ�
,�3�KyL.hC��	�h�~�,>y����PN��1z9\�;�W�����Gqv��UЫT&��t�P�y�$�/�I&�ǐ}N���x�L�-�j���OgtNz�0�������?=;u �T�y�iF����o�6DB��-���"�	���9yCuz�YO��y�QU�Y2�����*/���N"�j�g�r��ȢB?<�<h������	p?�T@2�+����N�@�O�����p[���	� ���o�4IJ��PG����l�Bݱ %C<Z��{�U��/K�&*/��4�E�+5=1�^>9g}���VN@dr�ʶ�w����2�ڀ���>!ʿi�I�R�R�Oo���{ܧ��>�A�s/�����jX% j�˕��@�h~Un��Z��.�`�p�Hٗ sV�!Q,�M���9��7j��f#_�ڛv�$���������L7d��J��EK��P�R�6=״
|��������H�#�.�H�?�f=�~pz�6^��Kh'�9�y#��ؖ����_d���k��G2I��j1|����F�B�Cq�2�����9II�x��傈ZV�������V����{5�Q-�Ql�� �fZJ�ͷ�w��xfp*��!�]�b}ǌ�����l집��E�E��hCTG��UWF	W��[o�+��\����ݾ�Ek�Z���2�}[�+�(��e��q/���pO$0ݔpn�Y��q\��p��9a_L�Y�7؛*�d_�@�����;�b�+_�,����{�\��z��8	��ז%��r��}�|�t���\��/}���ۇ���t��ԧ��#.|,$[ڥU����hϫ06�LW��7[;�w&��LCQV:�\�Qm�
�=��F�h3�uq�ٷ��!Ȓ_��,���N����\�fq�4#i�Yzy�m�	����&^����k� AA0�u}؛y.�|��u��F��d׳�v8ߣh��ƜZ5DSjə��h#A����Q�L�5�n�K��I��>t���D�q�C�'/}^��h[&�8�	�
Q�_n���r�OZ�	�{�Jƽ2�� $�f��n(�TPZ6�;��Ĺ��ڬ�J��׌jk���1]9���v>#���~�����-Y�雵|�Qօ��w���PnO9ܫm��Q�����Fo����M5���of���2�p� ԟԬ%�=�T{�{d��E��3�XQf�qy�g���U���/�U�R�5������n>���Q�L�Q�:,�Ύ�$X�i̵�O�%��B�u�uk�IP��������F7�
ٯ�-~�E����.E�)�ÛE�B���=�����2��toZE]$'w�iI��ZH`N61^�T/���P�CԎ�-`{�����4K������jK I���ְ��5�/
����U'�n|G�!���1��X�KB����׮O[�Y��5Ķ���8�J�1��	( ���2V�~����9m
B��{��V숉��y<߿��|P����5�o�����f�bJ1�o�޲\���/삥����{ŧT�k;�!�
(<qǛ9��i�k��(f�?��^�椬n����]���/e���>$�s�Ǟ��{��m�Bb�Q����"��m����P�'=�	�<m!�/l���62IF0f�na?O��8���0v�
�c��ՑM$V���N�[1 %eTu%5�΁1.�q����͡]�D8���SMC��e�>�����qU�_2?n�;��0�3c�V3� Ù���n��ɍ���y���;��n-v�)�����Y��|V�`�f�4e'��]�y;J:�$dݜ�VU��&�5:e2vƴUFu����S�l ��&]������;��V4�oK���WC�Ҵ;q���i��;��F�I^�&s ���Fr$J�4v����H-�5v6�@����*A�m��j��SnH����*�K,��SB!T毛�3��R-�
%��6/%�w�eÙ��=�"}�%E~����Q
9ܑ���	�h���F��rs�K�_z\q_�!��^����߼&S� 5iR����f��֢��Ԙ���{�kA5j�_�>����i��W^�\��G-̮͠;��1k�q���`]C��DU�
�ߔȯ�W7;&<������଀OBE2c�k�nY�.�Bj��4("+�*nM�o�7���Qfܒ[�9w�lژ�<!K�d�sV&9���ȭ�J�((�}���B�?A�䂇��":c�0��F	�zƍ���H���V��f�b�4��»p gy&$�+��
�% ϋ8r��J��q��j�W48�aV2Ez�`��V��@��Fwq|��Qϝ�\-N'}=�d��]Y��N�b}�F�k�A�"��X����R�f�H�q}5�Y��G�cE��6Z@�b4^���ѧ��/�%�§�iD���b�ƭN�s�|���;�QD����?��!i���׏$-��uV{I��\���{�ߧ\��,Oz��/||ޢc��-RC�S� 0��	��X`.6TF2�Awp��~�k��k|���JFԧK��b|�N�M��E�A>@�Yû���"�XqJN�ŕ��M�k������βVY�\?T�ޤ��29�j�׌�oy%Pf�$�L�7iwqAXO������P.����f�N�	:���/j��Z&(�0Rk1�CD6��(�b�(}���������9Q�26-�V|�d��E���j@�ulF	�����~�N�.�[��ȩ��n�i����26ֱ6�&*���u0�v#e���Z�F_�����<e�9^O~7�{x9�4�3���H䥇64V29zKO; %����%��q����!�X�#�t�`�Iq$H]�Mb e:��a�
�!�ZF��<�VhA��� _-xF���q�ј-`{?R���hC��|��C���@��(T�����'�B��S��� u���1�D3�S���0�xz �؁}�9q��Q�Y�p�;��
b���C�~��orϧq{�#�Fx��8���skV�q���jޡ>�Ltu�}p��ñ��&��Xw�3���Ħ󾯆}���g��;I�'e��\7�@�n#�VcၪO���6wv�!+�������#�'Ij�3&�X�)b�U�Xpى�5�LZ���Q)���t�1,�иą�e������|m��8q���}���]�Ó��)B�F@���ѤY��ÿ������r)[��B5@*s���m�T�d%��4�;*n�r���٭����h������a_TW�>f��7�P�� ���	�0F�z�lI�{��HeUs�6P�B��`�B[:wdS��k�s�~`��+su�UN�5�% 4q-6��?@��fǘ�t�����V�R�zh[Gd��C�� U��	h��9� +N�e�о�����N3�<��~[1�fi�K��A3].���d\^��.�Tl�׈H��OS�+K�x�P�����b��g�7�Md5U)Pr�^*���n�d������5�ۘ�M��_�z��U����Ն{�kP����c!�l�%$�f��_v��	7����VJaws!�s%SS%d5h�*�$'I�r=�-��N�f�������l�3�;z��Uݶ%s�y+�t�
;/�@���I�_�l'������/`QMN����Y���c�ITP�vX�^a��������c��w}�'o�%)c�~�,��~#;U�",��|�/�ɇ�É���	�/�\���ΗLb"��O$��m-%�߿
���@�ʸ�k� �Uš�����7�hS�H����=^��ss龍�̧ѷ�#��m,6_�-�>n���ZwQ��L_�߳�mDm�GV6��+�s�,�K�9F�#~#
�u�"	S\����Qta�.{��۰�@g!�y�����}����ʗ�4��Ʃ�h��q|�&��fs��ȳA�x��5���6��+G���&S9��C�|�(D������*�ul�ύD3�%}������&�a��M.:ed�Ã@y�n?��g�p���?i�����%��oM	K}[�k�
��;g�SO��x,D'%a\������&�k�ZZ.�Vj0*lx�_;����wtցn�`�����eھ��a��)O�m{Π���I}'4Rƒ�]	ys�e�o���� {�
{g��L>�v�&�4>�L~�C��+�q��F�iEn$�ܛ�km� �#{pZ5��*2��X7�LX���՘��pM�?$e� ��͸�����!:h�a��D�>̠�&��l)rY��q��y��,	9��5����ƒ(8��&D�J��M!YόaP *�m���*ew�N8
�;�of▙X�e�F�At��'ҭ��D�X>�H�7���C7zy����kt���?ag8�[��ٗ��@�cdakrT��0w��kָ�iϪ��׎Z�ww���`���c����	�(,��<B�4Ӟ��m���`�h�,;5"�@��:���T)���k�#�IU�;[��=�W$b�
��Tf�M��֛��,EoÎ�b��	��&�l��I:��?@�n�u=ü��*0�K�&��V,������z�<����pq���%s�.�j)t��L����.���$v��8��E����}�X`����*�'���_�Y������}����Y$M
��=��\!ݰ̕�'ޣ���
Sԛ@��a�y�.n|p85//�Iu_R�_�Ƈ��^�4�~�j_3�s�ܛY����&��=��+������ι0\r�3 <��/�L�MXyOQ�ɨ��}�+�OV�6s���N�I����`S��[�^�z˭$�Ft�v�ZG������u@ ��>s��A�I��͹`|5�9�k�dYno�m3(�d
2Gͯ����`�[x�����h�%�?6���:~N�y��%Q��ӗ�q����G���p�)Z5:<����ZBS�7����S��$\�v�F<���D;C����S�Qzs�s�� �VQ�
�y�(��Sk��O�]��tp+�l�:�'|������AT��Am���g�XR�:B�JE�fW{g�7�5�5���-#��D�N ����g�6�����}�W]x���Å��e	#A� ���I�kZ�Y�t]�@���Qu�;������P3�BY�#l�� �ĕ�OAw3ͪY���c�L Ly<�n#�+���0aoIv��*K�{>��EkOEVj�+'΅��1�k�������&����i>�qo�\5X|���O	�۹v~�C�~�P�8�s���q����;�5�*|�j��������R��$v�)~����i���p�r�g���y�t���pڎ�DE�����U���& ��,�~��.2�cC`h���i��1�J�~�X��.�v
�6�����6�r1��a�C�bh�IU����di��z{*
"d�m�r�	��V������:z�x�gө�}� ��� 1a���e�eE��pU�1�Ï(�X�����$���6n4B�С=Lo-��K�?M���42���T�2}��ٯ��y�������֓?��KO��`6���@���*��^<�z�\:HZ�z�j�S���3HC~�'��2���{G�]��=#��BL�:�����#��c%M۠�vF�յʚ|�Tw��J�@g&�4ݠj����S#?ޠ�m"��뺅I�,J� ��+C��g-J�(��z!��ƹr�~~ٔ�e�K�ರ'��4�n��G�}�s���Ⱦ��	.R·�ꚱ��h�J��"�7\X)Y_:�tbuC^ ��`(�>�U����h�Ղ���}� N��zk�l�+��;Oda�Wۆ���c�s}b�&sڌ�`[]l)ᕂ!6�W���%�v@FC.R�L�H�"���-[C�E�^�
G��&)�Z��?b��7��F����~�Y�W٦��}���C&�\Ή�HJ�,�!�@#]Vꙿ2QL��EU�dͺ�7(3�]�����j�U�X{T�>p�j�m�lSPB�Ú��L��x�s�醎Πۤ�)KQ�t6U�<O�6��dI�T�r�Tvb;����Imw�&5��P����\����5T���ш�=�4���,4�ŀ��wn��������!4#�o����N����������#�CnV�"����m"p��B�����d�:G3�
�:n���r=s���4C���%ѧ
��/������'st/K���d-�J&�[�����UQ�.��w=ݬ��0"��n��y���(�ԃ*3��	�;u�B�Ǣ澁�i�
ֽ-�"���N��Δ�"R��wp��Q:�'����)4n��ݔ�3O��V�����w��/�a�l�g6�y�J9�iY_҈D�}�֙�WG�r~q��n���P�0%b�y*#>�(����L����'O�,��8+��\iԊCy�~��\�ǳ9���3\�g�ܪO$�A��r�قC�<z����}3��Z����M��5�
�f��xB38u2�#:�M`-����Y����	��&^:����S��������:#��b�yBM�Nh�������kÎ1a3��!�{Yy��������ŐU�i�!�Nm�є�}����?�%kn��"s3?�i� ��{��#{ׯe��s�#��W �5d�]�f?�Л,j7]5����3S�FK�͊[����@��#��ux��p`f����
�h\��A2p!�ʓ_��֏m���������EļmW)���ĔѝSQVcl����C�"��3��C�7N�r��;bA=�$/�3e0�Ev��y�q�W1y�ك|+~<�M��YZ��Ý����Ċgjt��ԏ�a< ��M1(�L���ǥ��n�o?v�����G.$U����� 6px�]�O��������#v�P=��9�TH�t�=y�Z�H���@Tz��Ѯ�6��xpi�/����>�7���{����u[?����;SYN��D��!�d��!M��2P�#5VQlF��b��Z}c~-jk	���Q� 	�y_/x���#��:X�^M!TБN5�y3S������:	%6�!a���V�cݘ�#*<��U�7���w}u/p�'�q{�٤;����B Q���?�׭��ѩ�p�� � �T��M���"��߽�jc�o��bp�<V��W�����ZȺf��M_v$g�;��O8�ki����u�������b?S8�vPsS���y��T�7��y`�UΜ�A��nLs�N�'��~�� �Bk1ID~����3���b&����U���L�iE�3���x��6齾z��ƥQ���*Ve�z���]~�6�/�~C��=�,p�ϧV=��W��w޽�����D����G��]�y��,q���,��+�~������/eW*�l�=a�δ���̵T�B:�t�RrQ ��q��qs��h>��ש�	��G�����/�qf�
`�h�[�O���!^��<)�����zLl�(=}���gUK5�5�7	�B�Z�l�2�X�E:��M�5K;��7��P���mO$Zt���Vz
�G<Mե���h�m/pi'h0>^�a6��{Y�)��!fB:3��w�P_�U�����DO�/KW+���X>u�,��p��X�~m���J�}ԇD#��l���:�(�!�0xMr�ɛ�f1�݇]����Ka�9I,T��1;��+dP���[2���,�`�5^�*%����x.T{fy�zU������r��Yv:X���w��
��Z�l�3��;t�2tf��}F�OZ�w���Y�
�2�����Z� ��Ҽ�,�D�X��1v����K	�:{��۹q칯"eVސ���+1	�1�0�i�~�C���m<Y���+|�ه�C3|F��$���%f:#<G�����(=^��X��tK:�o�N�_��ݺ}��PIh���gˈ��ʓ��^vfP��,0�g�ZE^|�GGA^q> d���.�����)��bl���{��]��ѐ^0������"����ݒ�Q�����o�<�\nhi���j�.��������-z9L���Z�`ߕ���v������p�Jx�9M[��A����=ɝN�B��4!����Ы&Y�\�8(�9z	���!��T<Z��� JO+�p����0GNQ�ן�u_ �@;W��}���?��-+�	��i�z���kX�r楥q �Ց��ԙ�|�P�W`'�0��Q��V�����A�'�f=Yv~�i�o�u��ْ����|h�NK%�о�2\fm���Vܠ(�ƅ!�1"94ֱzhw�)��P�K�an��Vg!k�"���B��T�m��eT;�}H�U���a{�,���OI$Y���N[�yOD6�H���T�X�Xb�Wrb��L�b&� ��X��0$�G>L��V�iZ⺧cN��}-�$��%����G�y�e�%U���=qi��+O�=��&x��
�J���u�����8�7c}���p櫜�,�ՙ���;�'ճ�I& �4�Z,��
d"�d���:@���A��y.T܉�����-+��rdic.�i^J^S7l�����;�i�a&��zK��%�ێI�L�s�;�1��'sII��t�E�$�WxKk��fnd�\!�$c�OmW�Ja U��A���/�#$�������dv�.'-(h��v1��P���֞| ��Z����%1��b\Qo�?�Y��*s��ٍ.��AY`T�$�Z�L"jU1���H�xc��Y,��D�x/���9o�-�JL�<B_�}����_�)J`������`*��ā�[M�'͕��D���!�T�FX;�\bz�ɼu�>��^�VmJ"��mI}�\@vv�$l0%Y*=I���$n(!���ă?����q���t���Ղ�����0|�N������{��E�������A��] қ�1��z�I���{���N��;�K�D3@���~���%��d���pq�����_K�K6�;�s_Q	�����|�"M3��g�(}gV�l�҃�	.j.�DܭXr�����۴�a�Ï�'�\4/~K�;�T�H����9;95��^�,F��`c=�/��+�>������O �ZB\������5'�g��f����F��r�/p�r.�'�]�.������L<Ԡ ��PI�|ڟ�9��SP!|[�ldX�`����T�og)E$����<��p]o�����.G��� ~�n3C������u�?ݗ��l�һ��� t������<ʻqZtx��[�7O��� n��f���^3�v��E3���:P_:4[Ƃo^=:�y�
}�0 u+����B��⚷��G�<G{�I?�y�K4$G��_��*<
��(�p뤛U"@2��?ش�Rt���"�!��2tTec����C#�����Rq�j�_�}��N�0��R������^v��9����ґ�3��#a�9՟uI�dq����E�^.�6'��gYݢ�k�5�sm��r@n��[�1/���:�B�hAn���:>8P����j���_!US.��l��̋ҠX�D��pc\�Q-[G�7K��ӛT��cOt n��&�����Y�:��'`*�,��ך`���s,��}e67.�=&r�@d�]5��{O�j����]��G���s�۶L�+��o�j�0�tS����_Jt�ΒLh�b�@�_'S�Gf��+`	���
��m1�Xf���˿w��Z�ypN������&��w#:$ �U�
�LP����>{�c-��P�bxE��k�3Lf?<XaAn��~e��{Z�01/}���ʜ�_6Dr*�oV������I3z�:��h��Q�uM�k8[�����T�Yc-R�#��oJ���-o��h@ ��	�����W�a��c�%J�E<��WQW�7�ıꦾ�	��]r�y�87N%�ݿu�&c��d�p��]�q���Gˑ�ūa�g������B۫,�f��!��L������Ywu��;! ��;a/R�U��"(����"������#�C�ߑur��y�r\��`���}]'���*KxS������c�M]����v��vm���B �	gr�q��Ȣ���*����0�6\^u�;-���jzHo���D�4�����n��t����4�J8�*�~��L[���u	��>._�m�M v��U���n�$�kw&�F�`�T��ӷ�|+^��j�I�.ٽ�)����*6YG|U�05k�=J�Jң��H�J��HE&�B�����HʣS�tFv'�[K.J�����u�#���B��6�l��Π(K�(�@������p���|�`��]
˪
k����p��:���V�Rl<u�'*C�T~9��F���f2ol�������^���RxgF����}����cd�JU��Gi�,����jTOq�#j!f6�.�|H�׏Bz�`0�)1�p��峸:�@٥t�:C�?zx�Ͼ�b���sk<U=�J��,#���\3���:�g�㥖�1�X�m��f�Guya��8�E*d��mv)b�c�p�����I�xn���n�"�������ax(~fy^�\��Ab����vA#db���v��Ѳ�U���LP7Qn�U	��`|(E}'���'�s°��,�e���guۅ�-�u���\2Jy���p��í�o�� �?��@J�7%c��GG�2���:�P��W�����h���Ɲ�/˹�<���R13Ez����n'�<fg��LGH"�ǀN�;������1�xJ��/�i1!qO]�n�t�X�DHAu+�����m�=<�����$@�c�bkX|��e�Q�L�(�v�w�&���&�p���IMa���'�y���%�����Ѕh��E0"A_T%Bn��4��\�7X+��U��aԡm���pO�.�F8���G������`u��ԁÉM�?��z&�`�-��)�~�a��R&e�T^ݞ���M�
Bz�g�s�y����t��AUc�V(ؒ�]����,TZ�����ε�G��a�`�lw���$nRo�r��TUJ*�\<��
�di;Y��`izWz�t�\��;,�re��B/k����$5*ڲ�&�=Fo��.4�<��1�P������qu5�74l��Q	��ȃ&#����*b�ly8����7�m�k�
�9!��Un8;�_��]kKDq�Q��ر���s?�.$�K����%Qe-@��	G�O	�>~bkəo��F�'�fPC4�`���R�j)K�J�R�7PW���UU�7dۄ�}b�:\]�%��`��-�<:�P�.�6��eO��!�vP�S����q����A�9�����<�G\��:������le0~����n'Bjpw�I�g������_�d���tl��c��̈�!����K�������U��C����L9H��ӽ(G�n'�,5{�w3�#9_n���*>f�	q���Te+��b2����~�eDW��xm[F-q\vC4am��]��F�[�^�?��rņr5,�c�2�(������&��!f�~m`CC�I�[��xi��5�>����6cwhf�F�PHR�����z��͑0���(�y��-�'������%5�}�	R:�J���
��a�~��@P]�Ñ�|fA���@X���k<?V>(?gQ+�28��B�[ؠ���O)hB�e/��X[P����sJ��Ɍ2���bk6+:���KT�Y��	����r�����D��6�Ea�P�P�=���z�I>�ݎGs��U���;��W��rkv����\��v05&Ɔ��b~��I��2���v��nΟ�$kX���;NZޒ�ѩd*J_�}�ǡ�ѬH!����P5�4���F򖥚�ӟG��\o�Z��rB�,!�{ׂ!��(�t�r���%Z�t�/�-��Jh�d��eHZ���?��O��W8���>��L���"~�Ł ֈ�{8������TŻ;"��:M&>өt��5���8Օg¶����E8�]�����L�:*���6"�K;n]����R���F�8k�X0Aq�x�`E!]O]R���$T��Lwf,�������J�m��L^Q��ExM �ǵ\�KX�C��9�����.9�hK$䇧��_h�y���/��;YP��B�\�}��?��D�Lb�
�X׋�&G�q"��M}
)���8�RhI&�z0T����k���*�I�CH���DH�$ �M���,�{�Lq��Y�-g�o@�;�v<��>I{�Ya ����衊���V]r5]�P�[�D^^���IpSm��$�hl�\?/h��^����-;Ks*�f�g	��/��Q;��ք����KY��Z��4LS��Ц�m���އY7@�&Xr��;�\�����bp4(��٩�o�s���^��)��}X�V6���d���6�?C7�7���֙i���99k3[J��.JE�k��C�����7��[7/X)|n�;�߯�J�ܸd|:�"��6Q�R���G�J�@v�	�kn�w��ւBEi ���g��'sr�q����l�;1t����-׈�7`�V�Y8'z��7�t�!2�,2�D]�
��M'��Nz�+&�E����3n���Z�Au��z)*]�����1���t�'~��U-�Qh똒$ϻsF$�)��~�=&����_��З=G��jEg)�K��U�9�B?qX�DV4�!�S�F�:��m�z[�ˬ,HS��[�`F�>Y�L����/�1�<1�1�w����6|�����۽j���Eͧ�����0���f�]�
̗��
I�~��G�z�c�t�Ҝ���s2$�ـn���K�1^9S�ѳZL2������"�m��nP�^�E[d��;�˾9!�	�TS1���y�drͰ&�O����vǗH{��Mj���&�r�#��d�N�?g?C�YT(�6;B[�����k�Ҷ쑊l��hi�͎�X�;Ԍp�՚�6֥�������L���ƪ/�ѧ.8����+�s~8�8n0�Bn�K�7���P�+:���&1�	�����5��|��b��8��e��!;�,W�/V���2�q��m����p�'Q���S�j�>��Ւ��fl�y"ݹn�e�cr�=n�����	���Uq�|z��Г�Y���o�? ��z2�����&���g>��=��@�,��8Q�L6�m��GrQ��	��(��� o�.��5�������W7�eӋ7H��wn��g~�OCH�*����<��Y�����Q_�s����<ِum<HEY���	A�$gj�溇�����깭���6�[�Yw���\��U^�_L?�����x��\�O�?���d���)|�^�3oG���*!M��PW��Q�
�O�Ǳ�����%��T�M�NvC�[��{�C��)��Ӏ� �X7�8Z<��d�5�� K��t�N(@c�m�+�j�70g�/K�ݼ����3����<X�'���oKR��Dc6��gwX���u[�J���XjJ�ɛ�K贇�MC��[���yjLS�"`ZR�p�+�P
�콠��p�zB�s���C�0j�<��?�8$���5F�3�i঻*`��s�Se�����kR�}N��% L��Z\1B�e�r�Y�^웳�B;!iy���������Hs��+O	�Z�?'8��c>�t
 �O/0%K,����0�K�y��H��0���d��)�BQ�Q�}�Wy7�U��&��{Ы,Q��R}idjV�kN�G��_���P>2Y��J����\����fp&�H�g_�0�s�	g=�̿%��K�4�ZQ�\�pm=I��-ޔkc4^0U;F���|�o�Ϊ.��}���t��%�3�f q1X�I�ݒb��d�-|�zF���du���� �=%t>�T�	��<�5P�����9�9�{B�����,��aJ�����w�$�{�*�B~H���S~��|�n.�7�_ "�Ɇ��:�ە����?���m�N��Ȅ6��ĥ[\|Д���*o�H���B�xj��r9SW}OG�'�S�7��$���ʶ��FC��ㅯ�qrnK]����̺�<���[�-���]����"��j!�R>����ڑ���4�ז娷�azϗ���#͋��G����O�ݍ�PS��p��c(gsL�{�	q���bv 
���=�H����	�q�� ��Ƅo�-g>���c�L=�ѯ��c�A!.�v�]�d���ms �g]��2vr*N�:cE��Jh4����?�N�ܚ�-����+6��D��מ=�>�56�^�XR����e�/���t�9�b;���r3��g��C��QLV���0m��\?�MPJ�|��[�b�����]�gE�?�8l�~�hb��K$��J��&�>��ߞhډ;�s��}����gL$7��L�:��P�c�����$�p_ү�	ȯ/�Ir��7�T�~#��'���8U�L���ף�[j	6%>Ȏp9�,�T7�B.�,-�C���v4B������a�c3a����M�`���`��xM��~;8s���t���@�d����r(ܗϛ׎U��Ҳ3)�Is;M�J[�7���k1��Q*HH��͒��XpT){�����w��ׯE�@�3���2�"4�]���!�1�=�ٽ������[�>"/r���0��E2$��(��5���C��5�j
;�zr�ä�����͢
ϴu�x��}�%���x��;\O�؀z�Sma|2�cqԙJo���F|XQ?d���GD��H�9U)��P����	A��~�rGXU<�����"9Ԥδ����T�%m,�H�k]A#7Xj.w��!�ZRq���T�H(��Q����v��U�k�h�ő�%��ѹM����ڏ+V�4���#�W�lF1+�Cw�h�m@�k�|���'.�y|<2+�D�[r95gG���L?H��'C�s����8�qK����c��W-?�;y�뭶��W~wǔ7^�p�g�<�֛�	�aDG�:�#�;?�t�,�	y<d?~������uU[��!���m� <��]�8,�_\^\��g�l�t$X(r�Ɲ\���As�(嘟�TYKJ�{�T�=�n�^�;��C��JBCN������q7��{��>�O�O���6�ՐH���P��ʩ����),���C�l i]h�5(�/��s��H��Y���ƌ�D��Rp�c[�a����#�JY�Ϸ�3�"zr��x�s�#������N���`m��wI"UR����|��z�tYz�|��˟����ł���n��M�C�1�#/�^���]\)��*��)�L�3C�Øx���Y��>�.l-�;�$�{�ʗ��FH������^��Y�N�X�ťu��:a�"� 10�%��
�	��<��/u3��oo%���K�*L��
6I�	�f�R�g�u��h��=����/O�ɕ-U����4�#:É�ˇ�	m�D���ļ_��� t1s�����1�/���8�UG�3�F7�o;ʼ�H�`٤)�X�/����^��x��7��H�F`�6v�m�����␻߹�>�59LH�\��G�p�ߚDG�7�=������+���#�@�P�OYUE���{���` -�@蝩;�Q�Q|"hl�=OG��ʰ$��Z�Q��������iN",K0EY�Ҩ6�H��t�Vt����{kn��O:�XXe���@�+���_���	��zhw�����4����������)�݀#��D��Sjaυ鸥��!%8@x���.���O��F�F=�����Rq��¹�$v�m��9�*"��u��?�6l*��#.����l����E�������k��j�������T�h�n��y��ʜ�U>{c����WF���a�dx�H�~��X,k���^��G�G���z��S�66�1��!i%kl3�-���)��So!�|���mu��A�@�t7�/yςd�zd=AC��hnɋ�x�S��~�olG��!�-дc���t��ڋ�}M}Q�lx�`�(��8�etcؓl��\w~y
�IAI�s��8�X��������x~uCj҂��%�,E���Ou�0D�δW��Hb!W-��\'�}���Db-2��x�,�m�x�t �Obd���C[c����Jr�h)!�J�O��� ��6�]qQ��e�<ߘk�
(Q�ܒ�����/-�Y�f#�Pxv3z}8�n%Y�a�kQ�(/�%~��<��q���ϩ���n��
sCg?�N|;�w!3OQ����1c���re]��6��_D��N��1�E�) D�m��)��6���W��j�� �_���_BQ�p��h@|�X$5��CvT��8�$����W��<�����ΞDX�0��X�ܗl)z:z3������V�U;���qg���wf�z�wN]t�_G�>C	����w~:�[=~C�$�N�C�"D���c��+�d�;n���ڌ�c�[��y*� `�`�a��L� n
wZ�n�3��_������m���qSZx�͹ul8����q�p�7�NB���[�/m�
#*c�C�q�$�[[��PĖ���{���iK^r
�~�����hꛞ� A)ו{����#��L��I��e]B�3��C��Ϟ'����z�,2���J81��c"��5O�r��A�X뼛\��7r\0`Җ>�T�R��'�A�J��`�@Ɲ��T"�U#=-ɼx#Q��.�X��\��ϋ(Z\:��(x2X��qW�N��j�1��M̿rm?��_H���9B�⩎Ρ�U*������jD��`2L���]��ݯF��	�0:�t-��ц, �֭�|
�� ���ɢ����^�+�(֎+���)�үE(ʹM#���v�����ӑ�{��|mO���}
��;q�5Iĸ�w�eQ�% �����Y��e�e^l2U`����~�iO		l�jZ*�-t��p�MR��;M��U���`�����YQ��%��*�i���T1����q�?����"��OR@�:p�$ן���r�0En;{�  � )#N������=�'��ddIk"&��M/��}*�jϭ��+����oע�Ҏ
7m�=���GU���87�Υ0j:���\����a������d�<���l8�u�g3η�0*��'���XI:�o��]�h1D�}���F��qRMN��C^G�-�7���'+���\��9��o�CWX�� �r�:*�# =��
r=2�B����pL��09�TyrBR}�~����"q?z�K`�>�/�d�l�dgV�7Bm�E��_�H����	�y�]5Fe�������5��^�L�+���=4%w��g]L�����ZZ;cW�,䖣��"��� �D2�7�'�\���A_�:l�[F��%��Ϣ�}B��~#}w#i�htd�	V�+���.@���6����ywV͙��5a��F��_���H�T��¶9 �c��[�w���I*�y���h�-�7�ğ�o�?�b9�p��uS��TN�ǀش�ys�� W��P E4*呖d�p�����*���q�Df�q.9�@�=d��ń_	� Q����/֩�kS)p�=���5GSN�o�xb�y�In��}�
X���EE `}%d`Vj�2{�O��&�w͔b"�w����2�j��ib�6�9��7m��]:�x��/��c��p.�e�,�̳�g����������I�F՚�;Tw=j�Z2��φ�����AU�w��F��8��N��jQ� ���~5Q��#�֝���x��?���y��D%7����*^�i�U�8j��ק��U�sQwAMX�q�(������PK���~�쌆�o �>�LB�ɱ
i`+ۈ�2���n�\|���^D4Mzζ7Kޒ#$�
o�>j�����n���I�X�X��)���K�L�σ���M] ˎ8��y�ޒ����)T�K� ����Tݬ�ӶG�Fse��|�� �wqk{8�:�L���t�Z%�w�ݸ�^���P���F�S~M���$X��%�]�Ԉhk:�|���\"�B�P�����D�c4����e��A��)��#��PdbL� (X�e�Oa���@n��/�_�W$�.{���&j��~e��D85�>[���B�1Z�Fi5d�eLT�P_��Ӆ/��N���|7�i���#I�96ތp�PUF�.n=��_b�s���`�j1���I��Mޏ������܉��trݼ,��s�O��Ɨ1��_�/�X����Z{���q'����iX��2z%$G�B����"H%��= ����E�0�~o�s+���D�Qr!8�Ƣ����s�EE��㼐��&��<O�P��\�He2���
PFʝ$���,�a���W�d�0�i.tѧ:�:��: 5P���:��8�{i����V�{����!*=F�ҳ�-����Vh���e�&�*Ć�ph���Pj;r�Qti�N.S�'�������T�Uv�TnB���m��'��m�*� %��)�g�Ao3��Y猒�����S�|$2�6�����<�O�$o����U���1Y�B�2 R&�H�;�����I^,{1��N�����%���d?�%�^Y$�V��;lf��q�O�ũ�ΥG�<^5&�'U��͵^6��������7������
B�fR�U�ʯ��,��'�����ɑPȪb�(���:+��N�9 h�� ��}4ޱ���7he����7����Y5!�.s��|�a>�BH�����J���o��Ы���8�c�s�S���lYZK{1?�Rhd\!w��9x����cO�O��I��{��.�/.���)vp���d�?V�Zf�j�ׇ*pv?S|o�Gkmr���:��q*��Z%�g-Q*!.���2~w���	�:E:hWƫ�s�n!Uy��}+~���>�� �T2Ұ�+8�(z �~b@Y- {}ת=�i.����W	+Y_�t�_Ad]G�^��Q�����~nc���eg/�?ڳUΈ���F6HH,��N~6���2�o��;gD�����ޤ�b//���g����%<˶�bC�%b��<��E��qXF�ـ�ېsYoF��Na���E�{| v�����َ��(�Ti�%.`�B�BƋL0H��Kb-��\9��@��=*!�aS��Cdٯ@6����g��9p���L�Z�j��Uo����'W3�l��+Z�؇�bô�R�jb$�3��A�ۇ�`o����15X�N���=�r���l{�� �ȁ��F��IZ�M!#sZ`ǆ��hU-i���L�-��f�'��t}D��+��e�[3D`A��P����ȩ�i�����C�xȭw�̀�k�d���Lu��ȕ�{��7��q��k}�?��/Z�1#� \��Co���+�%	I����݂*)\�X=+����m�>x�:L8ݦn2]I���r��}�9f9�d�j�L�Nd"�uY`�q�����rJ�C��%�ZJ���lF\�q7�)U4Oy8)ͷ�]C�v�{��?<�DdSZ�B����x���ǿ'�*�C���b/ ���]�x�P;&���I=hy/���F6d�����I��b!�W+����=�r����QQ݂�=�����D�g��$�$��{gԋ|�J�fr�k��,���`�A���m�}ړ&����E���!W-pH�$�ʏ�+`+~��u��'!Ц�>@���p�U��`��c����U��D�&+(�ܧ9���8�Y7�za��k�����V��&����%x�X�-�tQ0&�i-Lt�PD�Y�����kU/��uN��*"�71�jd����Zi�=]g�7�hy��ȗ𼵿bq{��S��S����9�%��P�J��%���E�c�e8ƹ�C���F����� �����8�/v�q�O>xX1��o3�m�ގ��>����p���<�hs����/c�*|"��!y"�y�̵ot��3T�0Ӄ��2�	�\�]}��7���*Դq�Ƭ�/����`N��\��<��Ҵ��:�$p����L����W�b �][��טr�=JE|�)tH`�m���,���C$Қ��AJ�Q��ҥ�sA�7�刁O}�ybWd�h����e#(���]��`	BĖ����%��
�H>-L�	�$���!�u��)K@͐��>�|E�gɲ�e6�&�%�Y�?>���Go|�'U_S��\���]���'��RcO�1L7;���/���v� ��s���F�j����TП�J8�"<�EB]�I���h�]�4�/��@����r��m�����w���Ʌӽ��\�YRӻYh���{�G����4@���n�	�
5���$r&�~6g�xX��3.��©��V�;�s��x���y���P�T]W��	
�f?s��1	]�pL�nl�/�Fk M;'_(LAӝ�%-IJfzM�F���R�8}���V|��wJxa��]���T������0���A���#R�%r��H����%��A���J=�ȏ/����&`����Y�,�ʙ�hf^����A�߱l�	q�q�<P4qgr��z)I�������D�.o�Wj�l�}�o듣�z%.�U��x!��ag�s~%�(�^c���7F��Dr'x��!b�-1Z�G�@�`�'���R��^!J���ʼ_����ֿċk-�����>�oY*jLL@8���Q4�LF�B��	A1�y����Қ�E8���竳1��aT��$��h.ĭ�y"*������!,RC7��EO�V/��T��'��o�}���؀4̭�_��C��q�!�0%���m���k* ���f����3a�]3U�}�F4C�i�f�^r0��"lV�V��V��(�P��'��ڣ��d�k&��Ʈ��
�L{�}JVx�vg
�\��0��z]�0�f&��]G��
�ױ��X���YK�R�LQF!��|v��y�J.b��e���<����~�E�� Ij�B'/Q���PH�=�f���rsh�J&Hl�HF�T�;����0g1e֔�Q�9#�����t�V��.���׀�Э�jc�e'\��k˟�5������8/Ķ����S�0��'�����Q�̦�g׈é��-w��l�FJT
���Dl�L�jBش��`k1�p�:;;��%�e=	7R#���51]�)q��S;3���3�8:"��ȵ���\A/i t� ������/����[��S�4���QXQfC�O��W���#y���뾀?��6�U"���F���RV����=J�[���7��n�xm���Hg^J��ɏV
��Ms�!f��OͽVnB�Q����l�BX5N�HUC�m�T�gl[�Lx ;��QP�m�����	�i�H@�[Uq�/����sN�.��(�$l8 I#68�{yֽ��/ǳ,û�:�(=�_�a�0�M��ѹ�bє��6�-`$�M�Pp�<v�,��D���<�)��xi�ⶡ�Z"�E�*�0��E�{�����z����M������}��7�`�C8^q�롱Ҙ�Bx���<�1���=��1 (�@�ͬ|�VJzù�����T�������sfx뭜��Ѱ{Z��2��K""���[��kx[��RS�V}���q\X�����k����8F���-����}~oI��Ӎ��!\���*+r�;�2g��|&���}t��%�%]�o���\{!b��z�Z1/\C9!7���d�t,�����\b��8�ap`^ ���A�^���rN���a?���6`Jl��U!�ϣ��}-�*?'�( ��ܡM�#�$��P*lHc�e4�W¯�e��<�X�&+�*apx#b�&��]�)�f�L���9��^l`Y�U�`D\����4ع�t�_W�\d����e~�����e:��*�B����� 0���l�Ձ��\�����9nz��ڃ.HGX��ǚ���*��$�RC��|W��i�P=��i6 ��zXD�̻v��k*���6��	�R��E���g�'�6�M�Ih|�q)�TH��{��e���"���ݑ��29���Zg~6QjN'���W�f� 0�T��j�Xf�W%���P�p�?%�L���QF��<<��[���0��b M�ԭ6Ȏ�ѓ�c���ϼ
�)}f|+g��>B��*Qfq� ��Ώ�Is���߰����L�@}��8#�U�2�1�d�5�)T�gD��_ԟg��2.���1��Y����N3J�j&��M5�Rw����� 3T}�|��ɚs���{���@YR����:�gf9�;��9�G����[��O�Ǌh�=��T��z�g
IT��c�����7;��n�����PrD�z7K�jkX�0a_��q�|A�
`H�{e͘3Ml1=�ʺ��2*z�j?�<�� ��EhI�t��'�D�@�m����^�e	O^�roauU���X/e�?L�{��I�V�O�\�&2�]4K[~�Q��}9ּ��`����S�9y�nIt�C;���[p��W1�n�����_q��FY}�n�&]���ـ�'١��ۚ�Y�~v�8*�Ð_�� �u���|�'c�����S���[왱�#�)���F믇��j�g�^m3���}bg���Wb�G@W�����%���\\V��Eo���N_�T�y�Px�TH��M!�7�	��+�Q���� �����V�<�eIϿ���}���ng�2?ioO/F��|Q!�_�ƃ�H�pt� a4"���T��5ݺ�_�N5���`�x���B��m�+�y*�dfֹE&�;Xf����FLYC����8��"�"G#��<��5"��gd�m��>w/�RƝԦ�(���4y�ɔ��hNP���ڬˠ�[�тR�q4k?]y��U
�wx���Hd�wK���E���T�'�o]�Ra&(3�M( ��;ϳ�'�תOq�"RGz)@� jm�lQSMq.���&V�f�D�uEpS�Q�c��P�)�HG�(�?����n�� >�p�`��Y�ק��K�ۻi�	!��U���B;p��� �;l�|��Wo��QR�2%t���ou?���	耖�+����.j.�gwe�b�	��r �Q%M��}�X����y�߁�
-P������A���Lf�Q���~:
�김��&l��]�J*�����[�rm��ǫ�%g����<9Fk����RѽQ��>8�}�/�R&О��e��c����
�J佇���ƺ~��Xr�<sP�����1�;Y��0#0����#���Pٗ�&e8i���@lSej��c�^�+��R��+^8���/K)��Y~~*C��`-����K���	�ۺkې��
��PJK���I��(8Y�@���
t�A�3��k̗đ�C��c!ހ'�$،ߍ��4��Ӝq?��>yS�+P#ފ5�<��:��4%��x#���c/�v��_�[y{'����%��g��ړ�;�O�9��K*������t��,upx��@A����âU�U��dL^�������=��m�f����w��ew�[�hԱ�%�$.,h�3�F�0ȏb	錾� 6�7F��6�����T��N7�vpb���9/����r|�k.����Rb��?���{�X��������Ґ=�dn9�Á�����1P]��UӾ[�`
��x8 ����+��Ӕpg�d��c'g�b9F��6W��W-�����c�"l��lZe��F����� o8G�W�F"����@��</gܡ�|ĝK�26��R7c��Wp�nj��o��%w���/��-����0�s�^���M�S�M�"m�,B&Fj�8
����v��=��p�1⣡����
_��kL(���}�jo���ڔ!��o��%�CM�&��|-���?xq�[���#���a�;���f�J�ɱ�||ڌн�s�zKx*맸�Xb��A�fv���*p~�~.vI%�g�j!�I���i�?{�W����'�̿�k@#�Q��[Q}ۥ).)c�S�@vվ�_da?���O9�P���)�����%qG��9�i*�RyUt*e	���.0<Oԇ�|�^$o.vʩ�J\O�c��C����( �Sz��ڹ��,Ō�Ra֮�;+�-������'^�C\�C�Z����b%����䩑9v�a�(��t}ګ�ĳ����xS
�o8�xq��S���U����p������v�ٶ���q���w�M����E�rd�¿�����Ľb{��$,�e� ~V�}qȏ&�K�u�
��+�6��UW�'����x�P�ck�e	9J� gؼ�(=/���k��+�U� n-)�y����"~+�y�����@�����ko�H[�.>?�ق�My��>0-�19�.Vٚ���=�.��uH��V5?8@���m ������/3���k��[�	��\!k|���5����ʆ�7��ݪ�s��X���k|e��k*�8��'����L�<4�]{7��r�6k�0C�&L������#@�����v4�ߛ���w�5BpSN8cr�1ڢ���ʋ������Un�q��D���ҝ%���}��{�*����T�YH�8n�j���a�pO�IY��T2Hރ�|�tQ�����$c}H2�Ab����]�m�@��i��7��4�UA��-c�o"���z+�RO�q� �"�����	{��®�Q>H�V���kW�P�,�{Й�cѮ_�Q=�
�9�F|�aN9���(�$�A�Md�mQ2�����qX/)���zU3�mBv����I�C�2�<)d�Z�>��ʭ�?�N\~!C-�����OA���1,�r��W��~U�!�+�z��{��f�L�;&�e���Kgu��F�6`���*���%i2ihO�HzK֯e���	Q 6�Qr�%��s��i�E7�n-NS�-��2�ꘞ�C��]	�l���2��J�F��3����.�Z�K)��1�tP�ZjB'f ����R���3��3��M�Y�l/3ӫ�w�3
[�r4�dr���,b�� �S��4d-!t4��qf= ����Sl�v����K?^�� X�tV��֩Ř���}���.�Q�a��q�Bo���T&(��s����l#@_�>e~ڗL�a+�'���݇ D\��%����,/a2����j[�q"h-�C�~�� �	����B���N�:��qp�s��l|���)u;S�h,}OP('�$Wm�~��ͽT(<��2]�W���C=>�e����/���%s�cΉLfF.T�D"��t�ZjJyL�1h/��f��z-3�Ѓ�?��dX"-uB �s��&~�N�a�7e;n� �_��ej_Z #�-0]nS�#明s��t8<�'�Q|�E�I�/�W�]�"q �&�6$Sٮ�`T��y=���E���g� ��؅�o�y|'�\�}��n�Uv��v�l�����!C���"À͕%�z�J]�����z��iߓB�ʡY���V�'+�K]$_�i���z�v�)Q{�Ñ��rh��y���Y��td�7UgAZ��4�<0���;�l3�|�eF�:}�3�_
�¢n��q�T����^&o8\r�*<F+�V�&�ڮ����Q�����Y�����`�}oh�Ģ�]3����)��.S��}�
W�`���!^28Y��A��[�ThI:�L~����[�n��#�+�Ԍk��UZp��F��^Sg;!9M����|;���#�^�I����K��+%̡�Ǎ(5j�j��'Jf�H^+��=�v�N�P��:^^bC@^�a��JMb�6�{=��N�HO����}^��~��!8�HD�(��[,�����R3ˮ	�Y��X���Q�F���?�Txa��J~�_5N��L;�۬�Gt4�N[�y�`ߝ�m�@=\�R�	�(e������2��P0}�OD���g��>b�}wq����dV�?CC�	���hW��*�z����ڋ���/(��ۗ*��eD�a�S����KU�1sR�7ZPD['M?�S&� :��TP	o�	65ť�n��k?�O����M�,�Sֱ�����g��2%,ax$�j�4GFE7�}�Y��y��\"|�C���{%l���xA��۝S����=s�<5��Ąw�6K4�������v�D��+Q$裿[^ZF�U�$��Xi�Z���?7/3C�G[5��W�q�9V��w4���ś����&ec��O���z����N��8FG��|��4#ׇ�+�6F=�����X" ��ߎ<:L%��g~v$�FeP8xf�sYda����(��IS���)]tfN,�#i��j5���cdIj���&�}��� �F�!��]kP�E"�(6}���� ������d@�׮N4<{(RFU�ߎ6�A�[�[�2�9\Ggn�Z�X�@�
����NI8���t{a�Ft	oL5���@A�Y�M��L2�2�p1#UF�F������:�Đ�Ed���^�����RG�L(L�!k@�$#�8E7�kEN�Q;�|�E _� ۟ιD�\)��vG�i��*��4��C�� YQ&`��܈��ːGz�Q|��<�Qk������3!��6�R�=&�
]3�@�(�5{���pU�$2ӹ���V?Y���ԓ����ز���?q&/.鯩��d����]�R���/CSY�F#��G��d��gܼ�����J��p��	�\.1��~ϕ��R0�b������.�1��_�3ąaZ�U(�w�|��[$e3�$/*TJ�m��9ha�uaU}���L{� s80�
}��+&gg�(���vQ�%)�J�P	�����Gb ��96�/��״:n��	�2�0�2��j�T� 
��3g�E��m{��p���X:T��ݜ����xA�C+,X���?��7�v��%˧���������M���νM4k(^?|�2��nYd����E��� �
��b�.~��lKc K���~Q�%|����  �|=��Z��MI���\�\[�h�/)&D��&uWEЌ�5\�4�1l
q�����׊��6&X�����7��{@���a�[�����)�9��f]�i�UrnoP�|p����Y�/����5H�2�j��������y��!l����XZ��}1X��n��mG���x-�,0_��0A �6*��u��W ���orͩa�w{JΚxӅ&X���.]ύU�����Ĭ �z��%0RA�V��޲Z��E�k�;�x�W/F'뛼����pS=��=:��h����Of+��l�ݦ�\�)�EIˊ��--�@#zy&��X`Q1hol-�3H�`�~	��p0�~�y�y|X'��Y���o�ј�T�����j6jN/��Da�;��;�E�E9����y��h>��&Yy��m�i����B�̃���k�!�0��͏(���,������s?,9����m+F���(�h��|g5[�-i#I<��	�Zi�)����N��e���=��XY���f��o�>쩌Qy�q)��ت�A����ew�h�����3m��9l��.u�D�^v|C�e����كr��weZ}P7�A�Q��F!d������8�C3�i����	��ү�/Yiq���#x��$�K�ݔ4G}��c�������^�,�͙�d��jp��+�uJWt��L��2E�G��6^(���a*�Vⓢ�ۛ�A'G3G�ϡ��ba*��g�+�U�F>$^��o=����nhN�+����^�^䁎��"#��ۊq������/�;*�Ն�6��� tф �<+�P#tq�P ��o�}0�o�x�:Zz�5qoٵ�MF�ere������i�v�@XcB�G@���nؠ�H�i��y�1j�$m��͠<��o�r�W��؇���(<D��	�~�zb�� ��m�?\Y��[Qpk3��-yWA��.���G$?�F�A&�u]�*��ڮ�B�;��V�}~P�)W*�Z���r�Ǆ�����u�y��e�:p�L&(����\�1�|5�i��wo�����\3{�ύ�i�k��]\�L��r՜���}�����l/��[E�Y�=���D+jeY��1;�<0����zm�QAy�r��������P��S��-�͑�X
9��
g·8��G9V$��zy)�m O��+��(��Sh�p�;�lm �����QY�L���aM�o���$n�]����ۤ���1�؁��@Y�f��G�T�4{��K�@j��>WK�[q�
,�
�^�㘖ɣ��qf��e�7h�k�B+m!{^�0�a"�[��f�*�<�#���{0xO�� �	l0�3�x)�l�y����EH�Q^o.�2��=#b0/b^d�m|L�9�j�$=��;�u@=��B�S ��<��Ox]�*���Rv�L��?���sI�rV�R�>0�q�7)ʝ��-�/�;�S�V�)�ջ�����X(�mf���a%�T���6?;�k'Jx�6�Z���3��Պ�j���]�;�m9�R���1����Ȟ�*C�*�g,2�N�Ձ�b-'�?�,�~fA'�vm�{C�-�Tu�C����}�)�dJn�+��*�M��S�l�$)#v�/A�I�>s����9�uL��9R���Y|�uF��(�Pft��}�t(a������M2���(.���]�)! v�Waq,��z�6^}�&�ءϯ�O�����x��{�?���ɨ�`�?����0�KX�5,om���;�]��*W��Ak���Y�E�<t�>��1�顱��������N�0�i_:�%�N �~�cmO
�n��=���V󷨄��\�=��%ଳ䦴�ʄ:�<��?�6��nG����HR�֋?=�C�Z��*@B!�O��ʗF)"6��Mޭ�3K9�u�4�Q^_����v*�BI�ח��d3��V_N8�R����Mǁ,�l4�SO�B���Tܶ��nE�a�v�0�}� �(mt�>���Md�,?���j��vǫ��e.��*$`
�bK{�c��b�J�bc�3����n\2��n��[�EX�H�R,�-.秐z(����ٵ(���.f����Y�+>�4����
+��	��Mh���*�g8{�X��e�(����R��qA����S�@'�$��[���&}�a<�W����3��+F����x-���5�z��L]�L����N�7�%X�0�Aj��?�f�����9���c��WC3ih�0)�fu?�$@2�:1�*Ag����u�\�����v��X�V�umi�S�2�ǋxN�γr�X���m���3C�I��2��Y$��/7M�R���|_S3Wê��<<�O�X�;a������"*�{ ſa����.��v�P����	�`m��U�Ͷy��E*�hv���)����<�/�?)���e<\בV�O0��J(�����
R%�L�����G��0c��@?B��U��g�6v��'����)���Id�^҈����5����=��{�-��+���ly4��k�U0������;$�|��NV��c_&�d��1u'crՑMa!I���$��웫Sn����%ו��PB_�<�J�:Œ
���"ρvZ�RF��]o��������~��®wQ�%�;��R�Z�Ơ��u�\6	�,����q+�
�� Į�o�Ab�J���<&j;>b��g_οL��/�u��w
�Y��ޕ��e>�E��f�=
-ِt�&�Y(��m��TIss��{۸�eD�$u��])�lAh OC���9�*'�_<��AM���4�~I��o�k_��9�r�.� �q#Ya�4)�(5�zaI	�)��2�?9����q^�x���@������R{~c^V<fWc��N�s�d��M�Ra2\�G�iGH�:�� ��'2��v6Q��{�=��mՒy���{V�`� �(54�}��.ݑr��SJ�y(ٽ�Jǫ����u�J�)*���d@���Ƙp����~-��Ԧ�pw�=p�u�z������m��w��ק`[�� M�� ���u�����F�K�L_z�?�AO('ײ�O��A$q�G���ИA^��6R�3�W� o���ޅ�J�����|�J�%�>�i��jg2�v6W�E.�{]w�𔸇�V]�t0��(1�≲�z��HӦ�)��ȋR�Q�M*��/
�PR�c���2R>i�h���#�pIzA��)�x�r;��h����l/u�����{�5?�T��E-��7��wqx	T�V%���{����~��)��f�� G�ϱuA7�9���4�0/`*)����1"
�I$a�����E!�ђ�1�l��Ʃ!�U�hzcfX�m����;�X�`���!��ȫ�^Q�K$��sB�*�1lX'�b���Y�������k*�;>q%��٠�'�Х��o�����δrh&F�b��L�řbw�q�g��]ه��Ԙ��g-mŮ��66ە]�"J���*�By�`�NOx���	�s*RQ�o7����1"���Q�C���{\j��uCe䦫�_a|�	�x˃{��M��.G���L�����`ʵ[��I�}p0�v�Q���׏r\���E�
�F�oʡ��K+1n���l��ފ�hd-�殮�kM�KA�\{�U��hc_�Z����H��:8��W���>hX�b�Ĺ
Ӻ>�����S
f�a�Z�(��~�̌,"��|��}��w���J�MD�p�ў��̫���t��l�D��-}�w��	���ԂB��C����ȥ%?x
f؍A�7'��B3�	5]@�3�7!����Ɩ)��me���[K���Q���}J
���w��Œ4��<0g9Q�D����/��\Kf��G1z��9��M�@�"m�I�?J�FS���4�������۠�$�f��ư��1[�P��4ԑJ��j�����a%�@���3�I\�\�Ε��������6Bz} �C�~��3�?�����[��{jzk�S'g�����]�"qi�	Ix��i���pN� >������t�j���/H�̜���u)��Ϩ�0�,�n���0����_6j(L8S� �t�H�p�;xS�Z���9P�0�I,��I�jS�R� ���&��"�2�Uv�E{M��*��YAmZ!%�Bh��ɟ��3���@&ݻ���Z��*�c���T��+ï��}l����u��1�`�d�o����������KN�"	y�Y���f�Y�wmlk�<��I�H��d��Q�tLN�_n��N �V�d@��a�-J(r�U�ڑ=dq�ڭ�Y+�{�C��\���cru��������(��ߞpDI^1�0ң����kAK�(�,u$q�0�(�\�Y���'�o�� �+�:n���4�&y\�a��}3��{fB���ar�}�X��ko�~K�qoPT0x�e3\��1D��X]�G).�V��Wq���Ӧ�e�B���~T
aɪ������i�ҋ��3�9&�"��z^:^����"��"�e��p�ʑČ:`���>�M��p^�|ݑϙ����D�g	Z�V��d����k􈇋:�÷�嫾�L+��/�����?Y����c0s�v�Ĭ,쮑�����|y8!���L����N>p� -��(!�q��wd��5S��F%��@��9a��C#-w�<(!�~~-�<d�f�'V�����b�+����"l�T7 ռ��H��O<��ӂ=s��C�]��@���a�o<iunlVWU��4 x&x�ix���zQ(���Np���rB��u�{Y��U�3���,�Ub�mco.�p˛�X�� �
t`۟�I<��wM���l-��9�A�7\�I/�*Yl��
Tug��M�T��p����3�|�)�G�^mq�
����ݮ ��t�jG�NsN��#Y�t��D�(&a������3S	Hs����G�*�N�x J����*V\�7����!��d����c um�`�j���_ܖ�Fmg��,���5���L�e�V��Q�&��Ζݏ�lŇ��r�����{\��"�}����=�_�$LF>%�$hە�5ƻ\����P���<�w��0�*�t�o�>(z��d��:XV��;kI�DН�Wf�s�98/!?�)�N�^*[.5�M��qp���!�k�h<�?��H�č��f�a�@y��2��ⱜ#�R�n#�`N:��A4\�OaIpμL�\��z�"_��En�T�oϨ����c$��%Z8�z�~:遼on��.���s`�/s�o��y��9����YⷵI\|�HXWW^f���U��|a�'Ƿ�c2��K+�3�t\'#}Y�p0 �$y4�9v�0dU�GI �s�f�e$~f����qbQ��[=��횊��:�"[VR���Q��G�,��V�L�)��EDoE��u� Yg達.�Ei|�1�����q��\_�����)���y�qcU���f@j���~a�[�^N��B.��I���˜=|m�k�tа˚�#X)�^�W������E���r��҂��w�U�RO�%0�G纃3�x�Gו3���e=�ſC���ZWPP���_��\;Q���o�d���ѣ��l6����^�]h	�x�`��re�G����8�"u������å�+ۼ�]�FU��P����[]uq�uw��d�[���r�=%n��c�ӌO�n�]1F8���]�''X�`0����&����t�ˌ<����Yi�7
\�3 
���$��Q�ś�w�@t�E-�mf��Q��>k8�A�uU�O,�m�� �$ہ�.ʤ��3vH5�z���2n�����/�["SfqJZ�sRv���n%q�{r��P�����,�t$�X��c�<�tP��s8���k�{�f
�.>�\�p�#���e;x����^�&�y����nl����Y��zV�09�A�	���X�N��'`�FY�wT��?��0���x�s�����gp��K�?���1���@���%��ע��U��XA�HH+�AQ߀~�*c�S\�2��N�J:u�� �����yD:�l�ì>[�D�7ׯ�}��S|��"��C��:�Wׄ�꺍�?�>iY�z�H�O0[�W�.J�#�e��2��z�D�y��a��.��h���!�joL�nwOh�󨌘2S���P�x}�t`�!�AjCdks=��%8��V#�F�*X�4%$?��m��Pt�iFȎ)��<G��K��7���|�l�w��~��TX��W �4�<�;Y�l���.��^�Ek�IԎ���R博����׌B�G�<ݚ�)�����揈���*���[�M7U/�Yh�^�!�0�ĺvK�|��V�I�]����|� ���ͮ���-/�ͼ���-wPҐ�@y�K�o8!���D�EZ���n9�k�����j�������^�yS�10��0]}@8���dn�NM[.���[Z�|B�P��ԗ������+�o�S%����x�?/(�|���P�o��X�1QA�
������Tg��w��K��� ��I=�T��l��H�*/�����{'��O�nē�^ƛ&7�f1Et�������ѓ��$�xND�Q"oK%ɇ}�>�Wa�U�+�s�l�;ȦR;˩g��+�K�|P=؍�ѯ�l����ӻ�
�iEŏ�KX��]K$V �����\�8&��"݁�;�rk�W�W�+��,�(V#w}"�m����@�Q-���  `e �x��j�Ce�D�^�3Xm�h˙�S��*˼'����P��F��qi����M�% �;�$���M#�p�}��(���^��XO�rmJ�gI�cPg��c=�E�ղ�d�c��F"�.�g+���Y}3x�1>h���i7ў&�6_`���C����v�6��0�~�����2S��9	G��A�
1&�>����ĈX �Н;��ZX�N P6%"�3R����6��ȒI�cw1K�RLB����f�|��?Ý��Y���W擞�m�d95A�Ӯ�V���[��[��/�!��ظ�/L 9����^Y�sO��/D+�|�sO#���5|A�Xs�I~V���k*�<ixV=�����7�2@������\|�D;�P�'����k�5	��DC��4P!E�HϙTR(�CS��8��F:�'���O�V���ɏ����>��D��/~��y�$@���`�e���f}:������O�a��Fg�Q	@�S�a|�2�U>i��S��-.��A�L�o��2�_ �/����L�{_�ae�7�WJ1Jj�]Դ���G��:�q����38�eyP����DJ�K
��ZO؛D� >mf����.v$>����b�z���2���Vݽ6L�D=��� d�Ө���j�z���G�Ɍ�b+��#p]Ȏ����qE@	D��=~��ڦ<l��J,��ׄba��|��&k'=�9��L,a���hp��� 0����l���߈��d�]�x��he\��P���I�8gҟ���ݏ� {�d��&]�z�������^�>#�����|˂v��~�@,�%��\���cjTѶ��w��h�JrC�o
3����RȞJ���n~�Z�CU�O�}�w��϶���0���3���h͸�}nCCj�� ��y�T��Nꊑ1������ж�!O�n�z�x�Jj����f��:*�&��?a���!���d#E���M���90�[=��h垆*I.�V{[c�Ŧ��o��
㥑GLL_������c�{�U�BvYeS �}����a/z�,s�ht�7�:#}~ߞB*����g�5�m��Ċ�NR+���7(�\J����sj�m{T�}�q�ki~�;{�)ֺ�窏6�������������C_?Ar�+Ѝ�]:UY����J����S�lTڔ�<N��|S/�spi�P*e���s���TPyY�l��r �����TW��a���|I[~s���rl%+�,��s7��D8��^F4Hs-�R���rr|Ϧ���5l�x����9����%����[v|��Z��3S���j̻��z|r�s��~��~�>06=��]�]f���6Q�b^@�!���`� ���e��.��kV.IwV`�Edy)�v�^� Y��u�YMc�6K�����ݭD�u" V:W����G�s-��� ܇��>k?�Fv����e؃�U�� 7���	v�~�q�v�:u~���\�g)���V�Q�I��ܩWf�0�U�9��5�z�Y5c�0�MuN�e�����.�4�5���y�$���ր���U��-�1xM��p�9ƯS�@��ɗ ��pd��J�Vu���:��|+���N��������.��D5�:�����+z��8M��A1�� .��M%]bڞ̈�H���kdښ��)��#cv9��J9��G�
� �eV�`dl�E
~di��瘞���]DQ��Ϯ5���ؕh����ϲ�4lJV!��8��-zYg�� �n���X�+�(d�p�͕.�� �@�t��S�G�M���踐��f�6�uD�=.���,d��2�|��9�ro-\Ϩ�lIG/��׊�PU?E��-1�N��c�h�a[���J%��of4�W��o\���ܧR�F�-Bd%����t�H��%��d��s�5؅�������F
��z�-4��{� ��~��f�,����&��!��#s	�b��}�^�dr����>X���/U�,*�y�((h�h[�٤=�Z������P���O���d/=�t%�8ȗ��!�p"��_jZ��j���ȵ�Ed�d�#��L�\�f��Zؑ�̿E#:I�y(�uPt�V �%;!CC�`�3��s,b�3�	i�)�g�4���T����e?���r4=r���=H�(�蓝�>+y��\����TY%�o�$��u��sԹ�PZ��E���)������Z	y��)�D�V0�R`� v�4f���3K�y8M�C�l\T��ٙ�V�~h���	�	I�w�L�ڙ�2���Tp�� d �&H�M��(:�*�-j�ļ���tq�0�D�)�D=/6�����;�>Gꏸ(��0r����Y;��u��p��[���}<�:��g�l��@s�rU�5����׶����4�	�	8M����{��Q��д��B�^)��d�"��I���(�6������G��ŝ��"���~a,�K���U����(���(�ξ`7���'��'��Q�pxcq�IJe�˪7��y�8
�r������V9٤�ggB�/�m��MqB��t��W+�x�˼����)��f���I�l{�[��Y�3�#�G�P��t	51C�d|���tEAB6���R�8$(^�A���h �H�y�.��j�z�O'}�XRٔV�d�+l?T&t���%�ͺ!�ܼ�l�se3ߕ;2�.�2|�KvJ�`ǈl��C��E���0��X����:q�]�0{�:ga�ӆ�ܸT�ط�Z�#%��؂��r�U8e�][����a��@�3���K��������I��jǩ=����H	��92�QP��V_I�����I�<�7G/�=AM���<�����֛��t.s��vg��}ul$�����/�U�|4м��֚[��o-�X登�b�f����ȣ�ƻ��ac�(�F�0���Tgψ:�q���� �H�2	:pmQ?
캈��ucV�+#�N��+��.�%�A�i�
��׾o.��#�Du���^m�4ID`�e\�����n�p�m���SJ���ĀcNX��1�~��@e��Z��	Oȅ�X�BG*��O��
�rVW��6ݭ���#�R�����L y�ǓnRhp�-��ʒ���q8�gx/���*���@ RLU�.��q!,ds+$ b�n1��.�<�>&#���Fש�Z�
"� ;P�7�9�m�M�L�G�ͱf��'���mS�I�P7[{����ꑴ�Ç󉉘>]��쩜+�n��Tp�Ŭ&��%o�E"�bA�ɞ#�vp�?�r��"�'�e<IJ�!��
�����Mr�����B��8�-�=|;�ᣌw�6��fq]b�T�+8y*��UU!71�.�
��'�(�ɗB���y	1m'�
:N#&��٘����T�iy:>���![Uh��e6p�qȿY'RD�b�v�B5߄\Y��"�*e����rQ�7�PR��*|1~����s�dP�6A<3����g�3�݆�Yx�8W�V2�Z5��-0^��Ѵ�3x�W��4nq� ��-��X6��z!`��*>`�ڹ"0�)#ë���%�?*�\�� ������3�x~�qkd�aS����p���w,�d�&Atp� ������F��_�N�!xP*[��j�."�?HJ${p̭�����g0͢riQp�k��.������~����#��\��6�\u�Q}D�GR���K��ҋx.k?�g����tC��.�DnC������
cD ��7?pn�%�v��U��-�����en�N���XE��
��M��9[�2����K����R�|r�ѯ��Ұ铴�[V(�['�q�z�P��^Z�̤v�p��h��WÌ|T���ec#xȪ�|Gj�|�9�	~�F�[)S}7U壣p�HQԊ��	�rT�ꕑtLt��,n��M@vMJ�?�2\�MN�o��탶�Xvc.KE��d�d�����~ˈ4z�L�o�~Q�J�֮����ĵ߂�37��!���{C�ќ $����%���� Z퉐m��a�"H�?���xt]�N�֞���=���������	{\g��Ž9���u��.y�z�N"/`�2�v�A�qg|�ľѲD����ad��y6�f����K֭�L���;Oy-	B�VɂD��i��Cƚ���۠����+=V������	�(��z5�<"���Md��y�7�L,C&�ۘ1�]�U?4�udX�O�2�I��:#������~�,1.�퇞{,k#Q�eM.�����d�r
��}�/�t�!����������+5�@fhzj�:��=a��F� ���t	���Nj�tT�����p5xy�H���ƻFj����F�9��\�%�ڎeX�[@��0����<��W���&�p��FxE��U�&�ҽx9X��_!Ja�M�&�f-oQ|ۯ���M����N�s�vM��A���AVE�i�?�s�}��$)������q�E��%�ɼ	_��b�񭏆m3u'2�׋n~��l�D"���#{׭Ew%�C��3|�n��cG�C�m��&���m�Rʐ7g�5F��h6�x6"��G.�ͻ��7̉�&��&�$1�]e^�M��pL���s�<�Z�w�S��z�����4N{"�I-��p��ͧ-4N��L�,z�!��bV觹3=�Dk���rH�.*4�q�1|�l������tA�2{!C�-�)6��ON�s޿�7#�����܄�]��gk�F���IN�ʓ/ ���Y���WY����a΃`[PĻ��]�6��� ��=K��Ԛ>�M��RգZ�ǒ��̔^�g��r��O+ՠ0�~K��Ĭ�Ќ�ڿ���x��GQh9U��g#����e�Tx�-�6]'�f�si>B��/�J��y�ײ'h]��Q:*B��*�I� ����y*F$s�����?�������	]=E���r�%�0����jk�~��򃮝�EJnU&��f�,�ꑔ�D�}Z�*�3���Ү�{���&�$��e���c^�YS�QdE�n.AZ�
��7Tᇾ���}�N�+��K���m�H�PU��T{�pSJ�����T���O5 @�ju�&=X�cO��^��b~����
]Q�2｟R.�����B��s*���a����r�V63�F�7J(��n�fͯ��a_l5� ��)뇦;�t�����i8��{�9�f�*[q���>��I]�J�0�G����qLl5��_���3�dk^of
�H! �z�D�Kq�f-JBc6h�3?���	�\�6;y���⮧���#Ytx��se��TZt���|�; $��a��$��H�v�
�����w��a��#�X<2�҃�|ʝof��������k��;t��]�j-�ZD��ݻ|F�[����<n8�����?ɖuq}�T�B�W������&X�r?�g}{e��ط�OO�(��Mr`wʃT�9�O�A�e��xU���T�aG�����5�m�]���A����{rC��z��D�n�|��GS�{��W��3�Z.!��ɵ�~���-$�ǘ��&X�1lrQg����跉��o4H�܆-�1������7��EC��[�n�S~Ȅ�#�;�A��[��vU�����-Q��u��������	f�M�}p�R�j1E���y����F/�$5��)ps	=�:�����t�;4.Hü��]]�6� �X���m����X8�FrU�}��1����E�et�%��5�?&��lµa���a��/oD��k��M׉N��j[12�h����dg�&�e�I'O�0��PR)�A�^�Bgd�?�1���ħ?��Σ�����_-Y��}~&;�@��Q�ٸ'F��$kS���O&As���[���l�ӕS�#b�X5�$�z��?�( u=v��M<��GƄ�⓴I�� �b\Z7�;��%�B�u�=t�`�1
U[)CH�3�'"R�Wc�x+�]�p�F#����3ib�)��s��.�Lh�1�q�����b(�Ϸ�G���������a���d>Ws���K�G�1s��sBh��y=�yD(78���j���/���ؚ4�6���;k��a�Ye�z:� �g��uNK�Є�����R:�u��.�w�n>i�P���dJޖ�ٟ!�tY��%�-㵇��;��������������������,yKR�@@������F^�V�刉W�M��9Ye�2"���|'~!cd`�?g�D��'Mp��A�5LA���C,�N���%�5>��б�U-��Q���'�7�]@o�)O/?�Ց��mE|H�A�Uǉ�^���ްM�KdSE�A�ɻ��	�te�u��5�O���-�J6�F�j�=Ͱ(6*�Yt������׹FG��OM/�u7�I.9y}q�OT���߬Ϭ��^��L)��tQ��?�׻vGfO��EqJT&������b4,	�,M�&����qLY�|W����~;��YBӞ��9u���M��)D7S{h���獔=xҨ��?�%qhE�x񇱢�3���c��)�.C2=���!�Zo���0�u�X�!��<:A���
+���ss��L�2�bK�n_᯵���N��f���A�pd<s��L���$��=�[e�3Hk����&V3;���#���Y�n�	�蓒���S�0ϖ�
�n�iH���z�Z|�]qc�p�����XJ����oG��P=<��%���`h:�Cʟ2 4�(T���Z�m����I�J����� ��%lV��:[w�[���({iX-��^rh!�A�e�6����s9U� ��_%�
����Q-�q�����/�T}O����=_��j�2��'޾���E���ԸE3�s�uMA��}\��q���kxg��s�/�?jǡ_��U�8���o��w-;6d���T̛^%�{�2F̍k�{�\$Ll������' #BZ���B��l�E��A����W��d���ì����de��o*�>@��	@f�u�B4 )ڡ��a�q�[bTu�����)eQu�}�)PTj1m���(7dR��N���˿���4+0*>���0��g�5�c0�9���;Ie���R��$����v��!�K$)�X��nh��D�.y�j�g>�.{0!ޒ}��DXQ���7GA-(i;����ljW�`wn�����i�^��ޤ��.��7q�������l�1bC�OLկ��y�X8��V`!���v�2�����L��#����s�c�:�6Є�e��C?R��p�g>I�Ll<���X-DvU���{��K�_t]5�-�hv�?F�@X�����Iy��v4d�;�-�M烖�M22��2�[Na��ҳ��>S4~8v�郹��;�X(��?�+��b�V]TǴa:������3�ܝ�(�&U�;�X��1�&��1�Y�<b'����ʦ�������ξ�И�"�!�@����]�CO�vw����k&wȝ�6FB��������IO��ᢉ)�æŢm��q�Sv��O������FW�}u%�U��g#� ���P����P�.��#Pl�E !�
kVo��D}$W��.P���5������G_M��YI���d��a�������0IQ?=���h,A���@�5�&��GhCV�����s;\�D�4���LSP!��]TG~G�ϛ�jr�I'�o򠠎��,�`� 2�	�Ӝ[&ã��$g��Gܵ��GP��k�3�v��J�wnJ�84�'�m��T����Q%�u�����_*�����P�fJ�ASp�~�T���]���>*/Ad��lR�N}z��������\�����.1ޞ�Cc���uA�gfjV}��/ɂ���xt]�)��oX�S�g'�w>Lթp~���'[�e��IB��Ϟ��g�̈v��go�f��y��������y@��*GՇȹ,:Udk韮��T�7x��*>�"�$_ �"�t�$x�^������g٨#ŌHq4/�et�Hـ�C�`͹R���f�@`DMȂ���|�Z;"��DQ��"�)Y�e��mñ�7��{\��Ωh%%��RI,�2~�*�2� p��~_�Y(l��d�����6�~9���xB����w��d������mw.�Q��f�*��*���f�8��\� o�C5O�
�p�6*�F!�'Hu���r��x��
��^�3�J�
U&�&�V������|0D�jYU���Yֽ��X��ܵ8�z1����f�y���qʷ�
VŶ՝����f�����jl�q)/5�:�U�7Hۂ�~ʟ�����+F�}�=OX�͹J;�PzIVˤ��zB��:��������E':�k�u���B� ��˙;�N�I��	גS��g�pSʞ�_C��e̐�$4 ������aPK�by)�0'"�k�Y��/v��US\z���I<)׻}ϰ����ElH�M�'�V���p���<B��u	�*{i�b�����kQ���_�(��NxnB��{�"��n����� ��%8�7�L�^I2;�ң׸��r�#�Z0C��k��]bj�ig����mл���Z"���fg�D^�� E�������7���@��o��c
�Ұ'��O�^�^L����Qx�G��S
����&�C�\n���ґn�O���'k�c)�V�^!4h�#�i;IS�@�	8
m�Kg����^��5L���u�����{U�1D��UF'y"r��Ө1���+��F(�=ڂ-x��er��:��'�\26����]�K7����ݧ���Y��%N�j�T�-����_�W��Z����M���%�,$)�9�������L���!�3�-���u��ဵޓG��E�8u�}<�T���n��7S����y�S�=B�8�J~ ������Ǝ����4R�}Y��R����b������h����10��a���S/9��@����ɕM�tv�߶oC�I/+ۮU�^`V=����$���Q������M������#��4ص�"�2�y���I�4��N0�h8���g��/Nޛ��UW�T����$6�,,��J�ŏ��3^jO�����5�<��������q� ������6aI �=�]�Jl�uHO�W���cvG�M�6Zde<
H��w��j��kƹۇ�-%J�ȡO��s�d"nE�K��yˍ���2��j�pP)����S�g?\�k�r�N��Vۏ~��H���~�{U�@
I�Qrj�Z8�hĹ��Ոn�*�ŅMwִwR�o�a�
uP�32<J���q�/D�{Z�@Rm_o�-:3H�v~��=�'���En�<��l��ra�cg<;-� �M=�����{�q0�ËM�4t��<a=�ֿi�3]�JGNq�}��
��u�l&�
�K7�?�\(�9{E)3���$@�Fh~�6Ѕŋ�P52S��'�6�}4��lt���ϟǈN���De5�^��мYm���/�@IY;�j=�#�-G9�LWm�)J���`{��yg&����j�,����1O�*�����T���5��D�yE�h��T�]���5�����q�$9����@f�.����f\c�#�ᠬ�bޚ�M��|u�|��U�6	7.߉���4�ק�佒����~v@��oϧ؋pq/���9�F�5����ڧ�h'���� �A�2�ʢ����������E�ֱq�� �S	�,���� ��!��(�V���ofȔ�nɟ��﫧5��]����%E�o1�!�8"]��ߟ�IK��Z�A��,Q�# q���*���jB��t�� ��t�J�z$z�*�Ғ�]�Q2���@���JSC�Uf��ڤ�K8��ey�R�`�M�Yz^�!!�?~���F����GM/�e�.�������gpA[�!
�k|��
���ƥ��%*�0�H�yIz�4P������f���*�����9�%��ym0�͂y-+��֏����*�J�ҁ����I�e+i6����ѼŁ�%x��՜݂�n̌����=�}���N�U����e�U��/���� �C$m�*(�T�.�e��cc�z$Q �cx�kS#�dII�0��N#������I�Ԃ�b�*�@
�D�J~^����R��p6���/a=?��鄱G�V�����8?E���� �a2�4L^V�-L9j�v>��F�F������Pd#w�%g���}g�+��o_����p��@Eb�G��%Kж�lFh���S<^����p#㆔>�L
��zX�_��Ȯ�V��f��ËRUUUV����c�E��c���Aƽ�U,k�f��,�A��~�F熆��?���9۾d�M��(F�7k�4�ԟ5�mo����\�Ӱ�D`�U��UQM$IF6w���eb���7צ�� Η�K�����"�J�
xQ����a�W�K�� �s�����Z�fsJ$������=���~p�G�dDΉ#�A�%��b�P�'
�,?�8;�
K���
��aR�l��o�i��)����^.�k��0j�5����S��|�u�m�8�G�f&��r�x0�_z���[�>k���m�E?�.vC��BF8�7E�(p
*!��w�䔣-�����)�~(4����9���Ic��[���h�C07� cs�lUD5~�}N��,^ͧ���#����`d	T_Z�+oV��! ��>���C�M����)Ny���=�|D�jW	��!9��W!B�IYe�=��O7㜙�6�vt��7��nj�vV� ��1���Ԩ�Ƹ4���Y�.& 9n�4� �ė�O���S�������Z�k��HQ�?Z���d�魼l�,
�V���/k���:[R���fy�xf�����ւ�#%v���Gh��0u�/\���T栩��jZ]"�y즑ɗi���i���wd��}U<��]�n�)����E���J�Ӯ:�b�~��Z㢦��iYu��_����P�"Lx�q����TE|��@���ؾ c���ʾ���L&"d��}�8R>Z�a֥"��Ǐ��oi�X���:�v9^2�`�x��_���锓�Q�x�Y}��xm�k5ϔ��� �x�e��rB�Q&���IL�� ��?�x�h#��J���7"B'�����v��ؠ��^��G;���WI�%i|� /I�r�6k�I@U%���~]�C�E$0<���_$�t�۶�DcFy���/SJZen^d\����&F�Q��?�ږ2�]�����B)�~�1����;P���)��Em��t�g1NcD�_��:�����F�f�Vr���ŕC�FDF��7=�����%�\��	�e=Y�i�0_��'U��b=\��ƞxp�f���6�~p��o�)�"���YkEw>>����6��Lk٩��Է�Ir=�e��P�h���o�R����acZI�;����\	_��,-gk㞃�[m�l5Rh��>��z�=���N�S�31��`�<3�T��"/}����`u���.·W�wOKR=��������|k�n����%���㬏dїi��.7�wG��z���x�s�e`$v4�:�tx���I���}��ɧF���pp�s`�c�.���˥���m�����|l�-��w&D[��ǘ%���K��J[���0_��$;qMO
_���v������V)h{���.����E�*� ހ;B��i�-V��S�k��
y�������D	��3��"�6O,�`ȈڹF1~8�V�C�P��ӿ���_<�P�+jl�qT����]���hIA[�@�1!ttn��j���p�i�x.��T��4%H�h��J�Pv���.5���>�(R�x�/�@j�4	/�V֐�s2'����>��*Xt:�)�?X�,z����AEZ�������B�PQ:d��뤙��жˍ{�0Zİjm�ħW@�N֫$�)1V�l�G��d쮃���.�J0�����Pc)5��ڠ77G��uCo����OE����������I��ȲnX��;�e�.�k�`�8"'D�.�>��7��(;����`�d릲���,9��Jas�o,�v��ڍZ?�,�UD��P����{b�كgbn���C�WỆ���y�Mv�R}fM]<�� vYO�Htpu��d��N+N(�n�$��j_GN�";4_D0��m��F��P��8r�"r����dT�j��m*QA2�$���}�G����Q4�ռ	)�n��X�C�$���#p=Q8\�p hVS�f�!�>�	��?�1ᇞ��,bD���O���W�����k5�I�Dj���X�Gt���s�y�z���-Dy���|hR�{�4�Q/�����\!���s]��4w�����H��CF�ܬ�"K�	�����]"���ܦ<��@0!�~��ҹ�D�(O?����;h`�͜��V� �}�Q��Q��P2�M�HiF����{��ײ��e+�Ddp���)�l4c��4�� �h	
,H�8*��v]�^�$�h ���ʡ�8KH4�`8<����䨉����I�lؼ�i��au�梞p�
��r�\0�b�}��r{9�ƁcU�r����}3ζ��o� ߈���@�@4	�拳�U&C�0�7��4Vn$Qy5[�	�Fݤ%�� �^E�k�����\������"�R[�UQ�K��x��ݔ����ۂS�bK��O4,��>!�l�A�P�+��Ns�Ab-@��G�=Ecc�~W޴Pv�
�1'V�.�^6��ߴE��<��2�y�����E��_��m��� 6�Y��0�}�����Z����O������G��)p��.����ְt���nm�s�UqC��#k�)�6W�� ��G���]�_���=���1(��^��R1�N�ŵ��:*��p��GD���B��߆1��@����9�u�Țo�ť�����m�Jbb��T�i�8X�<��M�.I?򥈊E���S��*�Z�N�S�* P�_���Kn��
���M�ͱ��	5 4c�����e62��k��
q2����T^H��`s�-��BБh��^�_Pj ����r	K�8$w��P�wBKu��RB�"+[{Ԭ� �(}�Go_���C���k�zU���*M�ܳw{X�[��s���?���(~�v�푯��6A��G �6���Xk���I��3�0�1�^��K[�,C't3����&�ׁ>���!d9��=@{I���$�h�`���K�a/�萍9M�	p�� ̙x��v:�} �MFN�����ԩ�*@�w=�n�k�O�:U�#������Te�f)�t���Wp3�)�K$s�=Y,7�S`%8�A�t��e|�j���Q`���;�P����sj����O���*��"�i�����#Y�N��r��3��yq���xw�XA���k����-�l..�0����1vZ������7k��/)[���6P�+�G1�vS��\g,���c��N-np���t�3�ģIZډHktn���F�ӿU���f/�����u�� �̿�;��է���8l�AJ�y��(�&"a�~[4�.�Gb{���&��s�giG%uzr�o�Y���t 1e^E^��>n%�"�p*���94��;�s���7�!�GA<�Ǹ�uR=гr�>IW*�wQ����d.,�u��g�=ub�E�Pl���q�#y�m=c�$����Q�Q�K%�Ezb�l��4��\h����\�@�L��_���W���J"���G��
�Z���p%��]�(�m:0}�p����Cܥi�o��t&KN��ț�>K0~ ����6�'닛_�'�Q�6hd$0VS�3)������	mV�ֵ"�e,���*B!�3!�~?���4��}w��!6_�k���b\��:h0L�;�	�R���� �!>���hI�}q9� @�r�Q�!@&]�����,�|`�M�����*���*��l�$���Ea��d/��R���l�����(Κ��!�llSq��K}�H|�;�����k����Fp�(ے��	�P��7g�&R�����Ӿ8W��&e��p��q�����w�r��:X��f�)�_�°-w����_(W��"��R�6ͻɐ�`��@u���̕��s�;s_n Q�j�����`�� q�Z�u.L�3��Vi��DH���+�1YSڄn����d��yu�g��^�!���{����V���i���B�����,֔�5��Z��l^�@O�x���W�9{J#��JD��|cܬ�t^��L��6cW;�B�A�&8���-V�!�".뮂����%z	[`�����A��	�/HM~��
����4�8��WU<����3�cXoO���(�ݸ@g�f�P��k�c�&���4"������>�R�5^ݮ%Y�i��m� �Sa"S������RѲ�����^"9[���� ��y^V]��g)Kl�f���e���aj	Gk��8��	,/�8�}2�m0抻���*���bQ�B�pL���a5����`i"GL���;�Pp�z�����M-(G^�q����9Mg��s.��6��S�윻�r��	Ϻ�h��:d��+C)��֫�z{ۆ
S��@� l7Tl� �$�o��b�(\Ɏit�ȷ�v�Fل3����b<)�zz=�F���=	��/��� ���G~�D���)��[s�J�u%�S��@-�7��rT�M.��9�7Ęw�d�`��o���SԽG��hp��ͪ�
f
^%��#��F%D��}Jӛ~��|5ÊR�	�߼���R�ڎ�8�����EJ������n;����6"t��^a����Xm�����(5S�����("pF�&Y]�qF<vV�:�O(ND�k*�!�L�9��'�h�/kM��+�ک���(�$�U$R����?E�����M>���3}���M�K�X�hJ�6qa^kGIx*uR��Ȩ�����}z�B�x�'���j��b�Rw��!��hj�a2Y�?�;�f�i�2��*K�P�5R����8���9/@j�-��u f���\T�׮zT�S�m�/�����"0���#���(\--�H���'eQ�~��tV4K�nE�U�s�8��F�� �U��iGD�+62�`���1GL��9�ޑc�qZ�_J����r�"ƶ�w[5�q27EBM�u3l�1�hՅ��-f,��m�7�ʭj�+�F�+��--o<2%N��)H��lK�[[Ql)YG�����A����]�-��U9tm����{)�X ���������́(��aƉj�T�����1��y �$���9���P�yyh���[	�����4�����а���Pn��5���H��?*F��ʆ'h�/� FZ+�hB�����
����GvO�������)��W���uDt-���.�A�0$��R'�:�
C�A#��?�e���,"��ȏ��ą*����bO��kj��`��27��u�,i���anz ��&���L��YQ�!H�N��x�x�u+��W���
ŢMG.��ו�B���.2�l�a��k�f\�[��D��߁��3�X �������w�7o\?S�����;@��p���͇ޙ'���uΘB���CN3)֣���H,AV7�Fq
��Lƭ[���} ~�_��y U�>�J6�kº����1#�7l����T����q�55�P�#RP;rRQa����1�t�BP�Z_�]'��lE�u�D�u
�x���!��A��"	jn���΀Z1�<�͆]p$	~&��J�Ρ2i3\o�p(�9���݅��g���]����*TEK���/��|�����h�W�/�5�|��jy�K���k����F���L�y��=�x����i��k.ԭ��q�$O���}"Nt�)1����af��(�lUA�G���)ߤ�Y��/�Z ��6�A!���/��U�2��B�W�����m�߰W`4��J��Y�H?]|��3�v!�s��W�]W��~LG�L�m��a�K��p���][���r���b�����f�..��\���?%�>K~�Sl ��Q5�����;'��f�P���E �����gp��OJ+��#xF�X�=H��:��+\��ǁ��P� S=�SK��v�,Q`���"�����٘kV�iT+�׽�%w*PuS+��wl��EFf�^D9b��3��Z�mz�s�S�`��}�>Z�t�r��yJF,�S	�t�����}�OyK��3���T����N��#��^�$��A�J�Ŧ}��k����z��O���S��n�����[��o[�d\�YZ\��1����ݠ��Q��-��G��|�%65�\��# E�r�*8���d���y���^�.|Pʒ��0��G+"�O���w�C��0��Z,����FF�m�2�d�|�4���W�3���6���b�X�xQz��1��"d��Ia'D�v����Eo�g�qL���8KD�)W��t$&}4�����0�o��x����tJO{nʹ�C#;�fJ�?!����\��w ��y�{��>��s�b��P�+ޡctR��Y'ŷ�T�o�j��}z�?���%�dLЅ���#čx��q$�󙽈ڙ�C݂����w�����&��Tf�}�2�~9>�b����o�#MH������Ig8Ѝ	�ȧ�|��y���l���xI��Wf����3"u�H�zuF!�A9T�"l�xΖP�� �r���K�cK���Bwܴ���:̨���m&>1�(���E��i(=^M�T\�V���Ɋ)�J����GQv�L�.�e���?�a�Y��)�X�m���%�^��(^�_���EU=��ή���2^c��չ=B���.��h{����s��;�}\�E����������>�<eEҝ��FSJ׌�H���6ܕ�S�Iw�Q6�%���dI�I^}��E�:�K^��5�mL))�s�=�ҏ�~M�~>�!^�w��@���V�������<�"��-�����A����	/v"XIe�#��$H��ω1�ȗW��s&��
�󊪻"u�=�l��d\����$ލ4�9(���O�Tjy\uw�c\���\	|�iX������j�/�6�ӆ��x��rh�f�mF3h
�6IL��I_DF%��n�նVu
(DG���I]Ѿ����)��� }� ����03�4�x���ݫ@c�%,vX�aQg(�����>���E��R�Xi�1���ȼ��M %�4W=Ԥщ<�Nx��K���'ф�ۉ:l��ϕ����	�UoxlG*��ڍ�@nr9u�瀘Ɏp��Q]1>p%W'��Bac���Qb�^�4�����nb9h5����%�����U��	�c7���Z��A�s��_g�$��"�q�r�>����#X�8p�=���5�`�����F%�9�!�`T�C�Q�3�!�?it���a�3��,�TQs\��٧j�D�m�5����[�t5����!�ݤ�3fk��BM��z��]
=X?RNP��u���J6�qZ�����
�'��8�H�L���f]P��(k��&��'�V2Aghq~7�B��#�S*�ָߛ�J���`��Q���8�*�RF"��7@1�b��M���g�����1}~f�-D���1�76{��$�{.�q]�'Ud�J!��~\}��)eE���C��nH�������B(���N2T��"&�+�/ ɣ�[�@f�
uʦ7t.�2sNi�'����
?��(���S����,��U��j_`}���la�RS������s�����FZ$>tY��<�����G0E����8�q�����9kH�Y�Wg)a��X�o(�	���0"���~�L:�z�I>��T�8���?�n�8gu�c<Q^�Å�ˌF �2�({�޴@�Ta�h�,�+J��w�x�a�����#�~uW����uR����p'���W�n>s�_�d�;��=����,h���!�WQ[�c=r�JOݡ������nA0@���Q��=���*�g����0!c 
�/+��js�_8u�m^�`��I1ZDoNg����z<�6�E��۬X�
a'�'u�=&�[��@�9��XX��Dm��>G��TVd8^R��� �8��Anګ: 4W��	�g޴���(	�1��jZ�5��{������Pp��_Oz��fB��9��Uذ� �_�뙇���0��\5��k���.[��AQ�+�ۡ{�:p��@�%�������sr�'�6dD���y$_Qִ��fW@}!�a�ޯ�RE�OR�@�U���=��K���槉�r��a�Y��QHe��:#� D���\;����)�q�p�Sz�Ra�0���v���P&��u͵zX�1*���&����E�jm�4�<V���%��˙ޑ0⽚��:�d�49�H����f�"���V�V$���V�Vh�wA˨2�@�K9R��0�露���j��+��}0Jt���|c�e(
1����	�@fn�U5a��I��=B���:�C0 ���FG���aYoGP$%R�D�oILo�F����ӂ&�Q����y�#b}��E!5�78�=�}\�F-��S�L��Y��	/�|$ԋ���p"�o��{R�З��{����
��a��}
"�,�r��ß��+����]s�®��c�9�P�H�^��k�z)p��E�D����cHc��d~뜙v�E+���k��a�`?#�7�.�.�ඃ�ݏO��(�I,�m&�n.�S �~w�߱~\j�d�lޞ߅�;g�?c�=����mt.��b��å�>JӂZcE-LT!#x���f�(�>�nX�ܾ�N��"��m~��4!�6B�;?\����%�
G>\�k[?>��|ٲY:�/��|�?C(��O��I���Rx���%���Ӫ?��\�*!�D�:#"@JP'\ŋ�XҘ��'�C|��ڮ:+$��@�9l�����Jig���=�/[S2�c��Q2���f��I����z)�mV~l�je�Ӗ��m�M(�	׋5�� �M�v?�mS��itC>����	D6�r6>͊؊I�y��b0;?��S��+�ێ�fqYO��[#������𐓆�1K��L{���5kXaЛw��߹4�Z]��ZA�tT-ٛ�E~6XY��x(.9ɂ]=��g��^B�>�o�(>Ҕ����D�9 BJ�#� ��:�Wt\["� o+����Ius�V+'=�0��Ć�S%�-�����
V�(o/�|����A ��{
:�͔}k�G�4�S���mCw�mk)t�n�s�>��Ak��؉	�ng	}��
W]ΐ���{�za4�����|- �v�`�0Ha3(xk���Gh ����Sp��3�ώ�t���lP!|��3O�:6�h��5��P1��sh�*T��ak	A��IjޜZ��(��B���G�������q������.�˙�^�
Y��Pb@υeІJ� -[�ss��7�%��������m���f����_;f� 1R�i
}��B+F~O+֣>AR��A�$��-i��M��ʸJ{F�p���g��U'����'KQ��'��o�\t��dz��4�E��F5�*�2;7��>�8wЕzW��
�½S�� ����o?���p�?U
���� g/�+5Rp%�A�F��Ğ	��c�\�y֞k��b�o�l�/�L�ݰ�>��[��8��-��2Nn��SW����맠�G)v��5]C���f�ʐ��u��w��2�4��f��8��h�xO=?�뭷�p�B�D��f͸�:��.pB-u�A^�����M�Ӎiִ�O�]c���C��M���rv3w��F��	:o9+	�*9Y��y�A�{����X�Ok\F�彰��yj�C@HD7�������Z�r�媝� �>��:D�������d�����?S�K�&��['�i����VnP1k2�ܡUh٫�=�Av�j�����],�ǋ���|� ��3O=�ä��j��<_���ֹ+N�#�֠T���Ĩ`x�PIŷz�5֫`3�nkHm&fR��s�Ǐ�֩��h޲������
��0��/Ó���e[����/lJJ�rvAC愄K�&�/<��V1������i�]�^���`p��^���U���`#/h��;�pW�6:�6�?�nO�ޗ>����<�f;ܶ���?�Z��t#�J�Q�38��q���/�aJu�N@��)��ŹZM�mA����_v����|��{f�qk0xQ�kMG-7���a>�����:g��m�[�Q,�e�7�|:'�ɼ;�怞�Hg�����T�]���z�"�l9�WP�D���ׄ�p=ӴeIg0�O�df�>D��ϵP�c�W�0&#l�"���!�#�s3���f�6�(���|{p�� ��L}^gb�DJx߳QE��7����ё�N�8�slla��b�(_����ˌl���F7�^^�4<�#Mq3�S�,��5Hdkz����{�����M�B���m��D!:g|j:Qyu�P���aC��N��}�bU�m��~gR��<\γ�b��t3gS/�h���x�;^#��eO�����8c 1�{���]��0؀��jCz��3�j]	�Q�8j�o� ��>��x�����ڱ�_���.�SE��둾>(����"t. �1���-G�,������\#ˉ��OʳԵ���	�KTL��� ���d���C^�mAbGzCf�8d�Q9�4���L�Lq3`�a�S[��
Y[(�@攩ŭi�����l��j��;&��i6`˟���yN�K ��f[���)5'X�Y�KG�^�ǉ��Ǿ��(EP/��x"��Ǹ���D�0��d�|GK���+�N8������z�o�{'��$t�Q�۽K�>�UQ)Rg'�9�
}.���� ��4X�ne���5��L5g��d|1#i�'������XB�9��>��7�C�Rn�����ucd�k�k����/��8 �����H!�/�P���[�]��,v� &�("j6j����K�]��I�'s$��@H��b���E ����L��Β���&�s��|S�g�+o����C��.�!iA�� �6M��r��oH���>��@�yY���PX���ua�G�E٩�'r��jz�K�_2��Z�ʟ#�zɡ��g7�n���Gg�v1"�����$������W���k˽q?S��,��+v=>�x��5l�&�1px��aR��z�.rXu��-?��YIԃ}[� �w��o�+R�|R�	���{�2���v��(�I�IP����bJ�Y�SV�7G��k��(��q���Epe4��KG�d�/����q���m`�DE�)=�[�~��tǬ�z,�N7rU�$�c<��ݵ�GuSއT�ᆅ�Np☶��p݇�*�5�_y��kZ�*������������~���ȸ�����= +��+���R�˽�)>-Iup��M�o,5á=?6����2�`c�8�\!�����	��T<��ciW!���/eGY%��}��gV).\H��n��U(1�ߩ ��t�`?,P�N��ŕ��ޏ�9B�yboD	��q"א"ōX�h�'� ���ţ�E=1_��4 �+6!�)�^�Џ�3o�*	Y1)E^�^���r�(܍�@�mfs�}�a#�no_����bMSݧե�	�0��Ö*����ڌp���:��ɽ�Ң�'c��=�f2�!�mcQ�:�����q�w��.�2yV�aS(f����Z��|v��� xF_
p��$q�V�a�T.�K'*L�+c��:��܏~/~l�P4(˺�j���h#\���D��d�_����6v�øX��A1;~����ʭF_�sKÕ�R�MU��P=��D՟Pm�?��;��|� k�oJ)���E���^��j�@x�C��K��_,�
���ߛ�gސQ4��)?�$�O�Z���(�=�|Y:��9�~D����/��fme~4��Ŷ��^��Rxy��g�SiCb�E�tA߼^�4\�_4'��ȯq�6+cr��b��/��1�1I���mWwt�� ���y��"ĸ�N2��.�uÑoP����J�� �h\��}|���K�z�pT�_彶��n��;�x��0�Q����7+OG� ���,埆�>��fJZN51p^d2]�5}���H�	���"p'�"_���Wn���4d���%�֤ҊX9�6���l�
G��6�qWN�ץZ"���J"w�G�P���5R���c���ț辩pM��Q�h��~����re�f�NN�*F�cDiQ�5X�%@�?n��#�`�BugN���mN+Yڋ�J�1��P>w2q�Nl4�SV���>%|C�w�=�]�jl��CB��[P��s�>��4=YÀG�&�18Xr)JלN���!�V����N%3����>R@��6���@�լa&s�D$�2��,��LHKJ[t�V���1n��S�������-,6���G��'���f�a��K��iI��$<A�AO�]�J�dh4E*ӽ�g�?Ǡ�z�@!c_�x�{{�p�r�D�`�^c
6'O�0�D�DS��bɰ�P^;�].�~��Ś{i��|aJ�˖�F�1��-W#�v^��?*j:K`�-W��p�;6���?t ���}ݵUx������iq���p3�2���2؞��(���Q��<C���fy){��y���_g=_ɇ7?J��K�1K�!.��:s��ŷ�B���a� 6J�+"�P���(�X�;H'��U�� Z��\�pn#�r��O��Q϶���V�ҝ�LN�_Mq�i�\ȢL�n�o�ٱ]����}��3�\�:Ó�ǟ����*:LN�$��:�}�ǚ/�=:s;�i��v6rLd'$�����J��ˉnvʆ�Hz+!:#��� �8��[�c��J���s������@̌Xdn�w�㽊\M��K��퉳�I=�=��>mOcp��I���9�s�ﶬ_��rK�?&{)c�бL���Z�x1��:���"+ԛ��J ~���C��H�P{��㵝P�>U���d�+z�����$�D���N�j�y44�$�J)�x�\~ �#�߉8Ӄ����j�7-���V������s-{���]/Ŀ���grސq~��g�1��*��֩����b.v�=��ZN&�K��a�]�Ȫ#�P�X�0۪�&�9���n���ث��+ �Yw�y��aQ�S7�:`��N�����pf	��0��� �-��q���E�/*�;a��*�:ݏ�o�ٯ�͉�H��fu����%&�$A�gp�ׄT&aB�^f�����#=4)J|q�2ɒ�iL��lN~�����YPw�͐�xmP�/wS|�'�G$}�n��V��1�$�jAA�2i���7���ʃ5oU̡��X��5�P�fd��=f%�Q���*R�E�(���' �T��A�,���6A�N��A����<ca|&�y˷�N=��V�T�&Y?�@$ԧ��q���3��K����
��7B��H��Ll6wzk5B\�{iy���],q�~eM1�����o:���pc:�m%6�vQ��G�3.�zm��V��0e܃"�5�_>mf}q9Br��pOR𿓚��/�����gu�&����!�>3� /�?`g6�Ǝ3�p��MJ�|KjGE�d�E�S�"�����۶���1����k�{${�A��fʢ�����p<T��\��% :(^�N锖�BV�MP<��V���#`�A)�݉�50���bVe�^�w��"��SQ��;ӏ���g�Q���X���"��U�8j}gލŰ;˅��b�N��zx?3h֋�z�$X?����7!�PU�)�"
17 �xf�u*]��W��,|กH������,cb�L�/`?��Sa�Ej��(�X��CЎ�a���.0���v�	1z�K�A�٢��X4{q�CD��W��qʙǲp�PP<)��m��:]Y/��S�
{8��Yd|�ш�����N�7�$�D�	Ȍ�~��J���(�2|w<<��60cW��zv2�ee��=��Dg��v��H�M񄥏E�S�-&�_p.��́KW*�<_u ��ae��h��áG�:]���h�'y�@Yo��u�$�s���I'v����뫠��t#h����,����a'K(.�JLU&����Z(0E'�!����@�}f.y�-Լ�P)�h
@�,�Yص�{MAI�Ҕ�H���@}n�����v	c~E���5�:��{W���?>��Y�5`�,*oT��Z�?yf�P<S�a���5u�6+Z�x����L�C ��Mӝ0d�?7 5���ɵ�;����J�0�J9��ID��8��dZ1j�([��R�-T	X��ڬ����@�:�$?P�����/֟(��K��*�,�л?��ǁ��Tr�eK	����8�7�?
p\��vL��R(D\����?h�`�R�I�wS5Qxi�!�sV�C���+z�Jo�&�^�,�B�{)Z�7�{���p�_�2U���/�|Q��\����	��>q�E��S�;��D�J��fy\�m�
x�
��������ė�Yɑ�̘���(��G���]�:�Q8o=�]o��� "���1Fm5:��sn�)8!A�{4&��=�/��"G���<E���,�H�{���w��.�:��>O\��������mQ�S�E#nl0��n�,�\����KY��\s�����r�Kϲ6vl��N�38H�^@)T���4�{���IA��.\Q
�J�į��P<6�;]ƫ�����hEKZ��bf��ˤQ܊���Ŷ)4�Yr��p�##� Ja��� Rm�fE�ja�w�8
/�ɺ�H�'G�Υ��'ڞ��"��xx*�72� f����<m��u'���c�p@,%�{�;�e�x+�o5`�4��x��m+� �8��,�Oh�d=�U6�bu1���eY��hh��G �dW���<�"����;���=(g�݈�w��qÆBк� �;�ʒ2=7���KlP*>-8��9������$To,����V@��锩2��h�`��a���0��ta����l�O6��� y}�(fg���ǩvk��BCU}����Jv���F�Q�wxM�4h�O���m�#7r����^u�~<B2���H�ې\��'�~=��g�
�4�m@&��~P��4x��dyo�)�fţ�n���� a�҂��x�"�w�1.ġA}�M&p0ԣ���>@tn&�F���������� 5Xob���I�[�g���_LO����eOp�h�ɢ�Ŧ��*�{��B����a6���]1r��o�z3�ս|����)�)7�K�����	Բ�V�ĮK3󜓰�i0]�bfW슆)g>���'��X�/�Y}�&�����S>�dN9��e\��T@I�Al@�H����r��&��O�#cb������#�7O���m^�:Ō�F��kxYlC�8A��5�D���+�^����Ye��x�#WZM�û<�͹�Lm���ܠaU����8j������`�>&>���8���p�/�.U��J#�>�h�;�S���h����tWq6IMns���K@a���
v�އh�;�ɗ ;���(�W��iΕ��}����?d�S���ՇXI����x$�2Y�W�q�Ӕ6���;{�A�m�gLY��v����K{k�ƛ4���[ƪ��������\��z⡤NI��T0ܾ&.�����L2>޽����c7�F�`~��3>���*N���FRt�H&0���ד��;�����A��#�)&�"�W�(�O�95�h�2܃�����$��?����N��"$�'F�XH����r�S{nl��Zוˊ>��hDs��h�I!3+I2��̄�53����T�0�� ,N���"��ڄ,>5���J��f���|�<-��ܖ|�m�+��+&��1SܠJ����x��0�D5��L{��Su�r�7f$-�9�	$� \h.mւ�
�fZS&�����t!�K[��>�8>�C��tA��T�����|�NFg�9����w��{�7�0l��7Аd�+`�������'00���._�g��#��t�2c��?�]�,�Qe"?��,mwD��z,�I��#�+MK��H�����Қ�¼�ݢO�g�7�k�WCvWƋ�+w�)�kDji3W���DN#��3xMؚ
�L�'�y�i=Sj����Oq����M-0��ʞ�Y���C���uX�e���a=�6{Q��U�Uan?���`�.!��讯D���Ud�F��jy�}?'ns��b��a"�"i��Ȼ�ǚ9&�����i޽��W���M�бk�Z,����P�?�,a�874�32�鍘u_lz�lf:��.3�.��8S.U��}DJ"mqI$y�I�{O^���^��[1�腨S��Г�Ԓ�ɗg��	�������5zw؉��E&2$(째TW��ɛ�l�#�Θ�-�d�e1�1��.��U�Uf��~�&�#.|b����U=#�gt~���d}�'�3P���P4�Z��P��5���hi�޵.+dQ{_ݾ/��pU5�Y�(����q�tR�`t���S�`\�]��Sz���0�5���X�}2�m�6�eM�����z����(a�h������5���)�:"8�WS$������QC:�V��%�p3A�|O7�|���	� +�'H:����G�z��/�N��i��2��J��_���Ʋ?�T���!Z�#�ҥ"?j��X@a9=�[�U�y�vq�@٭P�>b^�Ťe\��;�3n��Pi�O>�{"���ӏ���Y���)1���{�e�l���/�'�~�j���t��ݤy)�떔�;.L�w$����	P�WP'����Y��u6mV���;@-�"��Q6~i�)��9�\��6)��s�޷3��^尀�kWMuN� �ZG�}�$�AtY���CJ�Ôh[oM�M��o�B��.��L�zت���|bz��&&�ryp��_]�M�A�޷+�=w��E�Z�xp��H�ItUo��D�Y!}��ր�]�ٞ^�]�8�fzޮ����b���z��(����|��Sz�x�
�<�o���_l��/V�v�	
�Lӂ�����k�����Wj�^��*��\@�)�EJ�؄Ǿ���n>l�)�V��7����Ic��jx�5�痐�`-��ϔ�U(�0I����iLx������vV�ɉ��Qy�Q,dH)��F�	�6Z�>�q�J�K2EB��<%�͓�r�#����b��1��r}+�u�C���<���;+�	ȗ�OJ�m���Ui�Gm�w����\���A�����-�t���|�L�4��}L���E��ML�o�����b9!B?��%BkQ9��؇���g�3jG$:�R�re[�� �rj�%�*�I[�%$o9��g�j�ar3��_6]��x�o#\�H_��L��i9���b��M�< �5܈z���8�?v��\��GT�8pF�4G���US�����DQ&ƙ�r��ÎT4v@/�do��-�4�;H9t@,�A:E������m�4���+7�=kB�+�t�xi�T:���'r�l.������ ^Q��}+�ޙC�-���<�lK�j��۟uCK
�V+@�f�n�]Up6��R��,���J�ތ�3 ���Q�v!11 ��.
3V��D>�7Zq�O�E<iI���q�'�jX�"#Y3�
rI�a�au���a�(/�Q���8�I[�ļHoʻO{����O)�5|�"�O��<���5�U�U��ں�EVm ���T$�+�96"��(^gďC_E��a� `�J�8�P
OF���4p���r��p6<b>2�t����i������Ţp�'��X��	c�qX�I�> '��q���b<����cv6؇�o����$�8��-g����d��a���5��u�]�N^�/U#d;��/�*���Zp`��X��"��B�s1�ъ��
 ��j�d��H����	��]E�����<~�Eb������C�p[���ȸFE�����NRI��*Pd��<��R����]�*��t�����7�GV�?��F��Σ ���������`�>�=<޻Aj�Z Ap�֩3Q�f\�U�f�TU$����ɤ弃�� �!y�Ș�˂��i	{�XI\,����}���X5R��'N@���
%�*⡂N��@��E�S�n�`9�lb(,cI��t/<��-ߦ��&M�:&���p�"o*��E�s]IpĂ��B��'�qBg�#ef^5I
b�q��n�#�m�k��<��6m��̡N ]��@�t��FkwƉ���3���LD��h���w�ߕk�\2E����q�4�L-Ĉ��B��d�C�P+UЛm�E�KR�T6����8��<�Z0{�0*Z�G�@�\oBԅ�3��z?؋*i�ӳ�h$D��	�V��q:w��5��[V^jloﯔ��ǝ�<�R�]��w�ީ�Ts����a�Q���K7}J�Cͱ![|�ۄ��Y��tܚ@G�<�+����^��4���H�/w:�������p��,(���c�:�U�;�j�2� "@�����6`��1 S2mu0>G��H%r�)x+�C��Q�<Bxچ�_`���Q|Y5'�O�8����qӶM��`k��t���AHQ�`�is��-K;K�4��]���� �;^a�K����B�$Z�#�W���|F��~� ��D� ֫�n*r������CC���5��v���h8�߽x�Skw�;�-5t��P���
�u���W�����ec��o�%Q��xb��ΰp�h�]4ʵ����t&p��M�#�^85 ����{�nl��vN��w�0n~�k7"F����D/�W�`V���r,]� ����V:#��ܷ	6�H�ƅ��[�bw/�Jtm�����w�a��9�_sxm�&�E��nX���^�O✅�<}!�	a��Ŕ^_9��\����ui��)9�@o��/���ъ8"�%�бI��!!�����]����q��ǃ+��l�M(������������OԪ�z�~��v�^�/1���D��Q��������&�?.����T��	uқWV����������t���I��6�V(US1��z����lR���kT%�&��MB�!l��+�8"A�	O(N��K�jJ����9պ`P5Q���{�;W�X7E����D�~l�=�p�����]
�W��(���ggCbQ��y�t� ���_v�S�J�?�	�L�<L�7"�� |�s#�6uKS_5��ժ���#��.3�*2X��;�f	1��vV"\��Ǳ��,h�~+]g�Q<�a�A2
�C��ɥ�ێ�|�����6���$|�D�O�7��8�HV�t��&a2c���"��*7�*�zw'c'�v�Y��<�%�Ī �! ��5Fc��7�\����4��zz�+UM/�Kb�Ӹv/��e`��{�V��w5���Y#Ǡf��a]���|.�r������N5���R�IR`T�c�j:��u���^�HĘpЕ;��~��?�ͬ]I��1�̂r6I/��_����(C���z!��*��Sm
8_KD+�S�Z]<'|�ɕr�U�5�^Z8���8���'��LT��x,<� R�'>�$s�K?U���������myk��n��*e��d�I���rA)��<ԗ�A�-�_,$�-ӊ����q�]u��龜>tz�_6D�~���3+�xn�ौH<l�ן�-E�z[c�u�e`Ǿ{a6͟Z��֢��V��pŞAɌ�v19En�I�>�>�z�6Nɻտ�汞�/�ןw��R�X�, ^��x��
����Wf0s؉�A�>�2�/�Ώ��I?fc����耓�����)H�)L;����t�-�[|���TW����A�l��L#��kn��6	���+�ݸ��~��m\�+� ���D���#`��4a��ੋ"�/mO]%����ơL%����om�%�R�6J���SD.+�.P1��YM�>�j��lN�hZN�e�y�qOQF�Y�?��CWI�ri�k!����d�LM!ן玫9��ᗋ��Ƨuf�p��Y�v~o�˗�U���Ds��^��id5��Nf�&F4��S��?n�������w�P�/��.˘��'w�/xF7���>����leR���IwA�.yT�l!WO'���5r����I�PY���+S)��h*���M���c�1��2�|(�u�}�������g��>���q��(d~�oo{}7�~�,C'#�"��L�R�I�8����9)���N΃�ֻX����S1��8'� E���S��U{��֦|�����~�JrvfL�0��^x��A��nQ��)��:��)�x�m8���p'9��GB�z$�)������
[~x7g�[�h��f�v}�O�:�UpN�o�з��>n#~���6��N��Q1 S��,-<Bq:��� �+�|������?��ژBǽ�1�\z�E��eB�{2�D�Hr��0Lu#�Ӑ*p���95�ʆ�cE$������Q��m���Dä߱���MA|�$�-�
��;�Z�����fÅl��	����xi�*6�$�i�b'�|	��DR�_F����0��S�ݪ^��&#��ǩ���H��8`:"Ԁ=�m�vz�z��{�~ӓ3-�k��lS?�W�:���%r&Ԩ٫��G6F�7��*���qY�¡L��c���;��v��g"I4���1';Nq5�{Ӯ���<C����>睖�$�� F�G��e�}�d /��i��4�Z�>]�>�7��;��|�l�����!�`���ݻښ����"ƠW���+ȋ8��5q���~�υR��/�d�F�_����SE����4<�E�#E�����c������ȏ�X�>�H)b�g�-�{�1N� ր'�v-A}Tq
�����7�%�G˲<��&��#0u�&��.��܎/|�$PK���㛂8$o$D�ADk�(=u��/<�e w�"�25��~	痿&��tl0�eH�e�Sh�� ����< aYq���_�����b?���R{��Ƈ�hdy^�-�k���4�@�����S,��T�6t�θ�%RzU�El?�Ʌ� ;�E�w������_�`���z��̸�=��Ǚ���34�_jGS����M���_���>�G$����Zے���Q�(��q<DO��h��A"�F#c�ڂp����<��F�T����A����M^|��9��-��T�T���>�SE�2Q�`y�����ɨ�ʞ�u�))��~���ٮG�뒀�H3�FJW,�2�!>��}��>��T⃺wV~�5��İ����裁�U%9�"�Z��f6��;ޞ^���)0#M��Vd�#}r�n��
0�C*r��䵟�ݍ�͌���[:8��a@ZiģFEW' 8Q�Ey�q
�=���t4�?ũF7Rã��C�~s��A����®���v	�7�:�����XB��>�{�"u�kwi�������57:�4N��dڠ|�j�)	Ye"�7�� ohU6��ĳe6x&�s�b�f��`�D7���u�Ր��А�η�b�z�v΂�s߉�6��<�����5����+Ym�9�����e� �BA��`���rF��ce挅~�2w���D��vCt���+.DĿS-]�c�=��M�g�,�4��Gŗ�C�3�~�p(�.Ұ����_U9���_��`|�ǳ�g�q��z�/O�N��mD!`Uxj�dҎ��Z �R�,,�����{�̸ Һ2������	�Yj��hM�b���aM���D�5?��C
�G��$�i��s�ҕג��{�d�s
�x�O����6�������vX)�a��"��l�1{�	�zw����äF���W�1]ٺ~���O|?�� Rs��}����D�-�A�� �IT#�j�Ԝ�����ݣ�b��z0�M�(��8��o�����!�!S�EV���*bW{�.�M'Һ�(?� ̏]}�$`O����{e�/;��8E�V��ƥx�$��G����a,y���$U@�B^v���μu�B`��վ������G�F=�Mگ�����g(	N�c�!���������+я�vXx���`��^e����P,�+���,�ך����k)��������#Ϟ�`��IE�'��kw�K�~���E�ke�� IB�+g�/*�z@Ӌ̃B����^�m��`9ʹ�N-�d=�$?�v�$v��Zmv��ш����*]nm��u$Y�ei�Í�(� ��O<�����C���{��)��.�fr��[�=���. ��
-<���j�/����d�ɋ-���gxo8Xy��qM;aWu?9ۅ?(������5���P_�<�FW���^*�~ �L����	�E� fF��'j�'�@2��d3>�S,�D���J":�^��af��f��X�]��+U�|9�h�e@͗sj�9AvG���Σֻ�A�àXn��_���3>��L�}5��Ŧ� �S���8���E�;|a֣��+�Z�_�t{�t��]��m�ɼ��E_#xtE;ƙ�f�t4fV��F�j�����ф4�dY�!�F!�R	*�$���#a\�u��CYB �㲵�!������Z?�>!�"8a`#��<Y��ȹRr��q ɨ�<����y���?Y��J�Չ\��(	��z���7���"ެ�W��aӑ�,>+���Y��B3�&h��M[D3.7�sLX.9���%y�*�� �"����� �<u��b���ѣ���N���n.FAO��9�"��E�RJ���~:�ayd�v�F�/e����0K�9!p9 ߌn��K��q��������N�����b�	3�f0�B�?D����a����lEUN�b�r���u58���!\!����� �S���Ic{��ˤ֘�!!��3.:��,Q��V9\D���� �ݿ����N��6D6�Q��3���U�����s`�8�+� ��4��C�+�']J�x��WՍK|&�A<^̅3��$>�^��$ O��SސG+S�W����Ӟ��[�{И��y~^���=���0 �FZ⨙Ď��T�8� +ˢ�!H&�S�S����KFԿ2����Q=�l ���k82G���#��P����Nń�P:g���6Z^�ڇ���D��N��]��U9~�H�w��"��e!���- ��0N�p�9/��%�X��` {?� �11=��]�d�ad��J(���t��*^���ͦ����ք}Zw���U���?-�*Y��/��vzL��Q���TJk�J>z/�}��sWI]�Q���:���7�E�/^���q��h�vG���;��C���jJM�<L�=��	�ZB�V�B#$n�*��𳤮�_U:�{��o��08�d�#���[�zrD�uh�enU�^�s�1P�7�����|$;(�� �W7�`�7���C�ꁘ���D3-	|�:�F&Ԕ�-3t�O�2���|��b}`�>m׻��)X摗�zYs O!T��܊Fe�1�Q�a�<�x�}�a$
C����qec�0�P��hl�������Ԣ���GK�!��[�M�yM^�o����lԍ�|H�X�� ��o��GXJ��.9RM!�v#��r{�Y��T�ɶ.�`M�0mЪ�8}�ݢY����%jD՛�Sz����A5y�-�(�o�쳚�7ѫ���=������$�<�q8��]H�/"�YD��D���%~�tN�p�z�D��#F�X'�[1����W�v�u��o@~=:JrD��º�N������lBI���Ԕ2��1�x�_�m�����#�,����׳}�c�C�ֽg�S���K�&j+ZOy�2w��J�C(�d�����A#�;V�c	�wY�]�+����A�z�y�-��hhq2����b���9�x��a�쩝jh��tU�:	�v�n�vˡ�Ӳ�R�v�U��=Z��̢�<��I)fx6��7�',Գ������Jȅzv��qx?�+B{������w�"�,��'�]O�'����9��������n��N�	�a�O�M A^��P�J �G�(��}�Y��d�51t�����2�QӮ!�ڨ	��Bd�04��cY�Z��q��U�E�ӱ�����h�*i^e����z�$�G1mm���JG�yNG�쐙��5W*(;��k�K<��3��c�a�M�o:G�+f��˹zk�)��� 5��a@��XmS������އL��,Z�ON0J��F�%�p=��5Kzˍ��d	�]p�����q��5�e�ڂ&�hٵ�������x8� �Qr�����ƠeL��j��%y�D��-�%,1��9n�7uV���R��a��M�Ԇ)`� �{,�+_2ŎD�c�y��<Na/�Cn��$Ê���Kb܍Mv̹`�]���t�:��ʼ�ڥК;�W�Ѿ��Z?ܝ����x��o�N�"���
brz�_=}5� �=S�QoM������֏9he�Cb�A��n}���JA;к�;'�E��s8�y�_�s����!Ϳ�s��n��5i�	�O��4���������Y�V",0K��/�ϋ<�����W_�����*�1b�'$T��tF"�60l'g��� �V�� �fB�2�������9L:��<v�w$�l���y�n��6��t�������o&*��k�1[��,"�����78kL�g$��n� ��
��B��2k�x'Ȏ#�� �k�L{̖e��K�V<I"Lax����z�΂�"����}�y��v#�΂����ُہ�o��6"к�*+�g�8e-�$�W
5��y�laO�V$?�6��Q�<�΍jW�!hœ��!�検6�`h[�>�)�i�6�$�+�O�M�ֲ~�����p\��ep�76{�`�{mdlI�����0`��6v9��#�.3��'���C[&1���Kʺ��g��Z�ܤ���_F8)�,���4x��5O�m�����ߤ��Kp�'8@I�w"�jUR�������1kOѯ�c�!·����Zܤ�Îou��u������yZ|�+6�اSKf|�~�ӛd�F�k7�z�P�iC��դxC���~������ҢpGm��q��T# �[A��T�O�&�?�r_S#Ra��RC#f8�O/�40<��'P�+��<���QF��v��6r� Hu���m�QI�m,�{�� �K���9NH�?��^;�����i$5�󳟢��"+�h8GVz�DN��U	�{�)�����K�'���m��&L�w�ϋvKAc�0���64����m�L�[�塞4��+{h�\���^���PV��G`qSY�#vy\ԉ0E� W�ot�D�Ο���P�� �ott��Q>,f�`B��U��Q��I�/W\Ml�#c^���M'�X��4���!2���Ϧ�Z��5���1S�~P���;4~,�iߗ��<�e��4�^���/3)�{��������p3;5Gt��vfG�؊<���g0	�rp���K���)H=��F}j:�ӱ���q����'�՛�yJz,'�,��t����$�
8{$���}�(w�G��u �G<*3y��~�n��49�%�� ���i�֕���QdiB�
���g������O�x�N:�{��&�l⁋5�	`Fb�Gr�9�z���hp���+9��op��X�sZ�#M�����n/��b>�������w�ռ��9�@L�P�+�As�:�-W6u��n��F[��zq�T7���d6��Ɇ����(P&��7���Zsz�)+������5L�e�B�Ϛ�@jR3ԬW�x���%�Y��3��ZC���*��S������JY�������{47R9^�m�P�X�+��Hu%%�;>�8h����@ޏ.��d���$��U��c�qZh�+XM.��Xl� ��q�� }�e�4�G�om���x¨��ӎHs�@���/���M�N�75_pk���t}v��-�]]Qf�l��rɋj>R�vW�fjv˯L�jTku'��O�x=���[hHM�����K��|���r<�I���^<(`,N�v`��q��oy�n\b{e�Þ�!�sG�Ꝛ��U�QOtp��#���R���rv_0�G�j��:r���p�J����j�C,�M���v��b�J�-����hG-�d�5��ju䞴���Y�1��fr�a/����˥�V<tԡ�8�/�b���[�V|mWЅ�����{�HC7?�A�H���n�r\�����N�O��\���Fh�5��������p��5����
��rc�����R��f���t�K��� �*"����Vzï�6S	o)���!g�HP����e��"h¯�=L�s�n����B��V��Y
Z%
Ο������ ��kЋ�8�;�sĮy^�ʩ���c��n�>f[��o�H?k�t=I99�`
�0�����uIj��=�Pb�'D�ڊC�R��D��f�c���64���rB���_bL�*��f�w��/-q��ą4ҔtV�-$��.���i�㍇����G�>��K~�0Y�w�"��)̤�e��1�m_�����T���g��%���f& �V�MQ�f�3����!l���~t�	O�9���1M���ؠ �#Py�w%TA^���gnm�@��ynoW�}�2�J�5]�M�>S��.��5�d��$����W�u�װ�:Y�׷.d]1�y�9�6?(,�wV &N�1::�Ϝj�ŽI^����Z,�~�-�6粓!������ٿ_zl9HF���[Xz�}m9d,�sN5���+�U��9lw;������ҭۻ�쒠4�n^&1��eh���06�u?ᾒB�4�r^��c��ߚH+#skB�ڨ��(�^	�����[6zf��tY6gM��9�7�w�	h�sL�>�P��`���o0�N�߂�(0Ƴ�S6DT�uU��%?�F�=~O�O���{�3�A�N�^e 4�g(O����H��hd|�g��>�Nr�߿q#�� `�?�Y�9éX�5a�9(M��5E���k�|=a�v�wi��A�򽊼��j��5�0����=��3�='�#f()Δ�;&g��X[DV
ቻ��,�]%Ϲ�b܈|}����z0"�>�:�1��	�Q�bB�}���gV^�5��ؠ��;ao��zG�
���z����� ������XDY��^�����R�+C_�������(��}wRǈ8Ys�������I��R��6e��N�uQ�kk���6J~�^�a+זT�E)#ԦM����,H�;���SW
��I�j�����@����������3��.�<��f�����d��_k6��;W��v"��?�6�����}��Y"Fþ��I�|��<3�lyn�w��#�v
S�)@��w$��d}�t��%�V�+ټ�2�(ֻ�G�S˱�.����Y$!&1������E	v����2���U��e��@�ǟJ�~�6����@�E���<�ʬ&Wz��,���5�S��rt>��S���%��8�eoF��R�9�Os��Im˟Z��3��xe�����NA�W���U���ֆ� �J��Y�t�Q0��S�O�V[����}�㥆����&�n�ف/�;�f8v�N܅��%V��.��˜���!����=S�ؒmDJ fvZ�D%	����|�.U��e���ژ��%o�~��^�����|/[�Z�=6���@>�iџ+85�����FR�)g���JY���r�@��p�/�}VcA��Ҳ�0���{�Y�DOa&X�Ј�t�i��	��1�&K���5�G�c�D��|Co�҂�)��A4?g�U�mQ���!�{�S90��j�$V�R����PD%��d�D�ZW���g/�+�kپ��,�s�0�hA���s/hrg~�c�H��X�����%0�ˤf*cS١�'o�,a����ڮ��3<�	�G T�
�^�F�f�?�ݕ���;z�����.��x-;1���-�ٕ�6;/5�Oߕ�M�S7&;�ʈ�	��>4�R_����7��Qa4A�G�t(��_�f�L��!@��J�FS��'y��m��<\U�S��.�l��op'�T06	B3����/��=���:�ԉ���1v�d��e���2p ƍǅ�H�y��E��[n�y��� �F��rz���-*'"�H�~�UT&wȵ��*�D�x
q�  �v��ހ�mHB�x'�5����ީ�F���0~m��Cs�j�c�Jn�㏎�~^���o�W��&����ʖ��k�=�/�p�I.��2?S�����=���lOl����?y*|�u���=�s5��=9�)y�e"(_�6kc�d����^�"v0$8������˚�ś�Ӷ��93�x[̷�ן(�$;�f�$���J��޵7�z���c��mm�n��\-֫���E�1�:x\���5�J����1^����"���
7��^?:ܮ���`pZ��V�ipsN����E:���D8i�uFz9b�\�N�;�A����m%��
����f!���#S��Q��*r0γ��#�Ȣ�έ%��C���!�� br9�$n>�S?�����+1���m�)�?����M}����y��*e���Z�i9=/���Fp�`շ�����t=
�
��R�N���m@k<���0��%H�_��_:�$ &�<y�=�r�}(;�w��)7^��$��&���J�q��]6���JI�Pq!�1�|��B����|��B�i�K�q�lH���b�K��|��ҁ���J@��!̜q�����p w»���}^I�F�J�GA=S�i'r�����ȡ q�_���}���Rt��Q����+o_}��K̆u���K4���({{��X�i��ô�2'3�dT7�5�';wb ��O�];��O���\4-j�v�%�9��Z�ˈmp+��q;0�^5*
x�
��k�"�7i�!�/���)3J<l���y�4�PA�Vj~3P��f����+��
j�e-֭��8!;��=r��=��x�g�2����]���D�8�%�(�L�EC��H�a��� �5�������@���Ov���G���)�ɭ��n[U鹣�- &!�7|ɧ ���10�	�X���lu�u�4�VK���\l��l�/7V���K��-m���mLFk��^GϤ�א]�[���X9�LG`̈�V�6�������oq}@V���5}z�e�f�jt�̸:�7����Q"w���|�c��Z�:nY���݋�ݦt���>0-|�� )Q����#�Lu����(��{�&�����Y�<���Q� )��b9��տ��X\<i$|��J�Ak*��!өg!6�Z���
���KM�]�ȩ^�: {{�ļ'��P�0'RI��K=����|\�ݙ:If>�b���29s���-�8�#���qM��+��J�H'j�z���Iᄨ�����h�-��	������s� ����WV�_�x?M��=ֵXSp@��Uy��D��vX�D���+p�Έ�Qr`H�+挓���!�覇wB�x �h���ڗ��2������I��0�V�
3 �P��V>��yj�kQp�P8~��&���عY��}R��M�t���y����W�}��[8 !Ȉ2�́o�]ڔF��<����A|���?�DVx|�]�H���c���Dq���o�x�w]<�z 5(�J��Z�[ۺU7)�H�K�ͨF-yL�X��C-83.�C��N�z�W�O�U�0�׻Z�
(�!��iz[�!����\9�+�w2G���¥e�۠�F��GY�^��.�@�C�Q�฀YA���*)��	�Рi[Jbn7>Wˡ��<99�_7�촳��2��$�<c����?)s�[��c���y849}�� �í�H#q������#-���Y �MD��d������d��:�e��xq�2�i����g��R}x�z��,G@K�5H,�.&��_�B��V����c����Ŏ�}\쯤��c�"�Κ�CY���d���:K}@�Y1�V\��ʞG�����������eg��z�8dl�D��f��@;��qu����d�P��9�k2O���Ȑ�Co%�+��u�F�<.x�
� )��7i����K����=iQ`J��s��~x�a4Qw�YZr!n����Am�U��"=��#�2�F��Euw�a����N��)<��^)v:�KT�:����|��ʎ��|MW�P�df�\X O�ꢑ�aY�*�B���������YȊ+�Hj���.��g�g�^��$�^|�%�S���,��b`���˿�4�_��i����Di% � ���W���Z��"����QT����V�f_^'�j_r"�����+5�a&��\P"����'��:�z�'�q'�Kw)�,�����Wۿ��MC$���n6�剝�,?D��I2���QT�)(��ռ�F�y%��H�,��)�M��>�����m[���׵R�rQ�Gao,9brc4	
���ם�&�c��/1�|$}Y]��~T[�g�����6�ܥ^k���sFBk�~�gƸlSS}�%ଢ଼�Ӱ�ܖ��{Ϭ��H��V�#��k�����4��B�� YdU�����8$M�Y��eVH���aӥH�ӭe��Z�~0�K��\4�_c��4D�x�u!� yz�R��bso�F:�Zn��*�*��8e�z�����kFry5g2/��|����~�_.?�UuO�8���~I3q��rpu�5t4:�Q�:n₤+}=Il�ե��`�r��wRf�;&�]de
�QF�)������[�����4){udUn���&Į�WhM�O��<��!κ�H0"̤�L������G��H�9�#aT3�R{�CQ�R�Q"��쟎n<=� 9!�3����MQ�ZBK1���'��[�2),���_jtOZ92�^f{���W�g\���k{3�W�!oHq\ue�����O0�����i�qyB>p�>ݭL�&'�FϚ�RO8/��r�?���D�g�e!�ۺ�Q�c!����9�N)G�"w�����D�m�P�"��GT�6�LE�C��xuF�R�
"A��Tr��J��8~BH<}���^Ʈ������&7���9�W:P��e򹒺�Z�`	!>f>��K^����s�ϕ:%g�rn"��� Ҟ�,�@cb����kr���~~�d�� pGv���-W����E@���L%T�S��y޾m#?�s��|7/�l1q8�X�Fn���tO����|�:�~u�w!.���Y
��G��A�R��a�#�ODi(����d�������_�s� ���F��m]�9L�
�wqQEBu|���·!�LV��D���K�a�[�f��.`�2����0�~�a���;{ ��,m�n4T��s��H�8��hg-I�Ƿ�Em��]OO��<P�?i�����).�u{l�ڔk9�k5�7�>@�'Es0P��+$��%��n�s�
�f��@���E\(����*@����H�b��`L���u�O>�M��
E����"� �.r�]`�rIÇJϣ�	?�g^�g���yQ�(PB��qǃ�oɵ�5��KaJ�H�����	�Z�,�?��2|���T��>rm�pd�Gx��T󀫻I�E��I�����bM�_"��AWA���k֛Opu�)���H��X� ��,%y��-"����Vv�1��Þ^&�^#�SAm^����\;�V�	�Ӈ���0�� R�:�b젊/a�F������#���B͗�	X �����Bd�J9�������hԕ��x��Z�>��ρt�ڹh�\ɋ��[4��M[mP'gW<r"���"`6M=�^d�}�$�=N($�%5 ��LU�=K������x�bH�|�\IJ��'4/B�Ef�����S}I�H������Mc�F^G���s�БpG�PC��Z�'������r�w�����W><�[��z�#JnWôL�%s�Ih�7I(���M���G�,�luDϛ��7v}��x~Ǝ�y�;�^�B�8(pKm++��ɒ]����J�C��I;\��隦��ts�D�9��
ιN\d8A,ֳ&mC�S-�7\�T�N���/"v��"�q~�ʪ���Az��?���0P���1��:���t�9,U[����vN]����@����LY�����LIDȓZ��b�x�~E�L�	Yy�PҭS��2����r�����ި|xD����D��爢�
��\�pt�o�mf�.�035Q��-��'��vb��e�w�'�0d�h\f.�V�R���F��C+�K2�y(���J�Ԫo4F6��s{��
�=�D��(:�BR�nʹ{�< �L�xyqX�N@��AÞ?v*� {��x?�Q�ݠ���&Y�DQ�|P}4R{ai%g��(DtY��	���O[w?�����iK�"u%@�5��u�/�i���$rq��oY�sߢ|#$I>I�	�q�z{3(IW���&�~���~_5�-cϺA�ǔ�`$���IVe���H�)���	�����V����8�i,'�B@�E�4:? N�s����c��d�9<M�y��a�����Tʃe��� e{�wDOUև�=�k�VtA�{�&�����9/3ǋH@ �7G�7�d�8��N��~��6�Rʘo���l>�7x�,Xv���qНpod�'�XS�:����>���y�q���lB��	v��/����)$LƧm_��V_o�`�tYe-��a�� ��d!��s�^�ͯ����n`��x:��ዣ��O:�m�p��e
�wZ���#
�<��U�� 
g_󲭪f��Ռ�*ҟ
��@�(�zK�1����Q$��g�p6�FBW��LCi��y�P��@�oۭ�����5c�]��;f��YS��b��#J�T X2�������F�Q�Sc7X)��?&���(�Aw�څ��TNM�>V�%�C���K�"?D����JMW8�~�,f�?���5�c�2އ�}��XoT��c��}r7 J�w�[�'��� ��9��/�4�jJ�����|���#��+{�����P��J��sep<�<��C?�'�#c�q��Y����m�m�R�\��m���V!hb��g�;����6�D��v$�� ��s�������Z$����m;���y�� �#����l�-cb��P��ݹ�k�R]�|��⩘��S���I��H<r�o���1���h1�O�=8��/�?��+4��z�K�ő��C[7�N��ZƳ�ʶ��5ZѧQ2���������=��w*F����5;�r6�8�ͧk�:^�D�)\N�A?����=sC�L ����˯�
�G\��O�n[DCڕkE7�g.�TbԋLL�ś���l���eJ6���o�r)�tz����P"5��]C��|�ՠ�"���~�It�(�X&��8~���{������O.��.D9�$L��%r]Q�6��-�	�t��hJ������4�A0��*��7��;���W������jf���ܜ��o+j:��.���1A��DI�o�0䬰���j�_K�v�A۵JԷӷ�J�L��Jl�3|��3�V=,���'Ju�%i8�?���rn���c�։����p����a��Z�(䛨C��T����,Kg'�ni"ٟ#�ū�3�� _�(�83��p0�A�<-�+�UN2P�G_K��a���Ĩ*�Ӧ>ؤ��6�L��=[O=�iS��x�Ce���Qޙ ����pŻ pR�DOG���V�.OV�נ�Z@��gH{�ԅ��VV3���#V����y2���fw���cPy��V�ks$�	*���[���w�)c:S�\N�j�-#H��ixƺ�n��kt�6^��攽78l˽�>�3aA���cd��<���,L�qO��edf�;�VԜQ�D��[�]�w�)Ȓ���iT}+�jo{e�Eq���0�K0�C�(�ś}Jz藙�S���u]�W�/$�zG���(�˩���K�!E�U�8 �������8 �����٩�rH�[�p����cJ `��������K���Ao�C��՗����_T��n��S�M���"�[x��a�*$���ןE�!xjX�l�i�R��	Wv{�T6 /�@WσN2�^"�h&���^�|�8J{��}�x��	J�OίB��x~�ڃ`�s.91��\�j��K��X��Ӓ�Vi��T32�D�'#��$L`�&@d�GM~0��~��}s`�B�ᑧS����hm���iQm<wqcR� ��1�c"R�/���a�H2�]U�d�>�|����^ŽD��1��F@	U?$[�[VF:dG�V�Z2��m�q;7ˆ�k����p�`�gQ;&;	��0�"`���}q���Q�*��� ;?N����vZ-4��R8q|A�ɩ/Qe3P���X〰%_�b���&���+R"n����6�T�O,p�'��n��%�� F�1x�c��#x.@�J�Y
�ߡʥ�t�̤%[�=$�in �V�Y��~�等~�mX�n�xz#%C�薛k�2e�y��^oq����%�ko)�pH�R�@%Nt�|���[���h+��E0ٓo�k��A3���g%b�x<�^�՞����B���[
�0�`�f�:#e�B��z�gR=�ۆ���m��/l�)'l5�)χ���y���f�WuebW>�sTm�W!tq�V��H Q{�����B<�;׬��S����YL#�1���a�X�l�뇱�B3��a4ҷ�t��N�v���/��X+Rq�� ^�:��������-/	��BA�VCJ��gVڹ��ö:����¶��Z|篏?�av�
p�����y