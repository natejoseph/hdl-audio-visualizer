��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��TdO����g�!\/�lmH&���� �G䳺�ʏ43�4�g����]���3p}�����ow�U�����,��m��U7lS������C�7�f}�qx��j6z�|��ɱI�U����z!�LXC>e�����Y&s�?�/��!Z�I[T���Ud}4��e���$h�_������Aϫ�޷k/S@���&���i翈���� �T���J�̉�5��n���f\K�rF��Rlg�*'�fJVQ[�Zf�*{w�~����r�{��m�@ճ7qk5�RP�טP7��`�����P^a��&­�,6�����`ߤڈ X��ODAv�X��6�g�d:GB����DB��5�d����NV ���J�&Bs�%~"��7���H�C������k�&e�D�J�?����ž�����dł��T�T��)�ܭ� bU�1ݼK�<���z�FR�忥��A���џ1UIc�0:�byue��Z6/��BUO�^#!�, �)�Z�f��Rz�r�B�&|��g���f�C"�A�;0�b~��'Z��L:v���[)j��5��~�SE��C��(k�`�w�E@�νN��؊$S.���u�h@Q(�-9�*�,��i\�+=��7:Λ=�8QB�ga�Ԙ��	G%EĖ��8��&�T��[&RG1]3O{uS�4����c�(d�a�\>����~#�oN�[�vâ W?��T�뺁�M#\gq �� ��ux%�3���VJpkz\&�m�_FQ�!H��Pǁ6S�)�|��rD�)��"������W\h�!{ÿ7�9v�_4���O=YLFIt�7��3�x�&�t5���Fo`>+_(� �/E�TKk\��6��._#g(�88o��~Nnp��.�����Qb�T�Re��ɳq[E��c��f�=9n��c�7��.��U}�`�Y>҃Á�W|7ԧT��1
쪳�Qb��rx�G��Ƴ���AQ��!>5�������$����0�Lo.��Z��_�3[�\t 
.���Sar������k�Q�-�3lі�R�nm�y�A�����L�����ͳ�U'}�er��ab��A$���<����en���R���o�Q	� t�w��|�����pl
=��"�k6�{0n��6�	�B_�Nb��MG-p�R�N���N����v(yX��6]-���U6�<I��cyF+���N��h{�~��Y���Kx�м�X�@D�u�`�� L�_�N�u,3/߻�y/�Q�ӨqSsY�cWՇ3���z���0rK� }t�[Rw_���
�΃�9�)���T%�����dN�TtWh�UV��9�٢��q��r��Q'ҁ�=�x�(� �I9�3|%�NP�,#�dP��Q���H�����X	����KY5�@+�Z���#�s2�7���X�Yn� x��7�#۟<n���k�:�v��3ȑ�l/
w���S�c:\'�
���������O���Pb���<�Nv$�}�s��ݡN��[0���h�]h7���eD��)N2<���	)X}mC�y#JG�#�!"��3y�?��V{A�w���,�(l@N��@�W���Zڂ���K��隃�]C�\�_RQ�2x�e�. ���#�$��KM�u]&}SI�l��Ӹ�/�����ن��6p��`e�ĝ�6=L�l�@=��dQ�ݨ!��V6�ZvZ� t��["J���9 ��UA7��tګY�d�Í~��bߵ���_�K۵�o6:�`ׁ�Q�Vlm(r��gA�����P�P �ח�������"���1��/nf�l@�\�����b�Q�1>��Qܦ�ܝ�^��! �����}��n��&Q�2�l�S_�y��e�f	�!���;�'����O*�١�ۧg쫒l�'ɕ���Ym�f�]�� D�0eu#`��J�W�)ʚ������I����K��5�x4�|�WB:ʬ�糸��uG���#�ӯ�i��h�I�~>��Q]�B�( f��Wvp�mlʨ,�Ⱦ�6�V�%��S���"�*Ƨ �� r��g�=&IB�H�T��h����6#;�-�l��7K�w�����q�/��R�� ��ݾث�D�[H���� XA�1=�p��l���z���	0'Ūx"�5���HJXa�?	6wc9��ڄ�ڬ�*ݰܭC6'��}k`zrD�ď��j���/`1���*�[PP�V3�ܮ�پ�鲂w��r)�x��S`��Lg5���������Y:v\��G���$d��	��ѥsx�GFΪČ � *N4�=�r���% ��.y��3������M�C=�P�u��F���$Di��AGB�%�.c�O�+]��.ձ�3=q	��,��l��f�7�D�A5�+��b�ܚp!��γ�(s��;��qM^��@"��,.g���� 5�P���I��0ɜ���c!��"�S���I�$ᱴ%᷀��r싮�.YˆK�|ڨ}�g�8�W�w��h��ϸ]�K���ߗ�DkpY�n�fz;������2�/}R���Qi���X+�r�,]D�%�V���$}�oΕ͛\�y�IN
��Dk��hi�h�Ŵ~g��ً�@J��D.W��a�F+H�D):�[58K�J�mlm�<~�]צ^f�Z�@�3Sc���F��FӮ��J2Dg7{��ϯ97�QI���	 �����$c'�eTP�H��!@2�GW���q1L�ܵI�ث���B�fP��� �o�� ��g���d� �/������������?��֚ޡH�a�)
���ʄ'�sZ���`H1?�E����zjYk�qJS~�
r"Z��Wgu�� ��Z���x�ª�xѕR��T*n��W4aQ�����N�+έ-�_�m�/l~��5<n���LRѥ��o��0��>���M JK����F"Yolo�v0;ao�+_cƩ .9|��6jB�b3�򁖓1�I�M�d�a���G���8y���i@��n��=)�����3��UDVnbBf�J]2k5O۱�MZ�I��) rI�1�ٙ�3��1�X��R�C�N�B�.,&
%z���1]�ƶ�A_Z�F>�R�0Л�~��imxMKUX ��`b��횇�Y}
�7�3�Ӵ��\#�+�P�JW.>�ϟ�L�;�jQ�2x^Y�ee؀ �ص��ɟ�`B�͉ׄ�J��F��Ej^	��+�i
�Ι�~U�d��N\'j�G� Z�7���iĭ�RpĨ�B
�N���C%�U� !��jA���f��,���^�1�zA�_�B+p܀/2x�7����P�OITΣ���
{�SG�����x�F���T�u��)(����d%��/��m1a0�n��Cmή���ʭS�w�r���8�|
4F}�Rڻ͹h�X,I6�~�0d<�.��W����*��xM�u�T�b#�p�p�S�5�כ)\5H��$B��6�rIY|�`� ���o�0����m���_PX3��@��6iåEf�w����ˬ<�fL!f�<���9�|i��ذ��/M>�s��U�J�(Tx��l���h���f��<�q�݈e��*����0�Y�R�;��f����4Ʃk���ҸA\�\���OK��e��z~��-�I�)nb
�g$V_,kzh!��t�V���Y��\����cQ�gΒ�Da@07L�ٗ$��u�pU֋��2ЦI^���+�D��=��{�[�X���������'�>B����e���������F�����GP�Z������1%ʽ,�=��y1����x#;Y��¯�;H!4>�i`򫾭�fBb,˅�)���O���x�j��G�=��d����8��>�K���k��ێ&�;����{+�tV��j�x�,B�t�ע�����
�J�N� �!��h�W�ӏ��0��y@$������R;��Vtb�����By+��̔ �-jjl!ʈ��5�DVs�`�y��v�Xv�~n{�.�IQHi��v7�L�Q��^��2�A��_��/�lKW�:|
M��4�Y.����,،@G+ϗ���>�!>3v�u�0�T��n�>K&Z���LK�W�8�]q�]7��>Z�����;#q;P���ki	8T��q�D8�m5YX��/��K��Ͱ�U*&d��x�������6)���^���ڜ�s��p�fV��N���p����	N{r����C��l�|XV���Ցƴ�^o]��%�)w�ᢁ�映���ԼB�aA>_�8��j9��=�uÍ�y�j��	�#�?)�a���\�`<<�ʷ�m���%#��*����xG9囉��#�PE5H�{��^�F����p�GMvn]�̬�l���Z�ENp�i���g�O�{`���E�$����wh��{�x�˝郳 �g8=9�6�A�tf��P�YX���R.����紁�G��<[@�9�r1�$�V{!F|�+#W�T���P����۫�8�)������-��KSx�3��xVZ���j9M��(�����
��>�n �h�ކ�K��<~��IkJ�M�$�k�:>r� T�'�Y��5��.����i.�����u���=R�C��m~�z�Sa@�4�r�o��v/�H׭�j�C@�QjOS6@�<��qy�����"U��ʒ�Ls�9�N���nd)��H@�*?�v���d ���s.��	���#?�S��V�6��&_Z���	u᩠U.��\�_Y��֤t��Kh'�o�|
x0_�c�7���6.k��'���n'o��r`=צ��p�y�ōAwi��]y1���]�y���؉ɶ]�o�;��?�'/�R�>��J�:�����?���V̐��Pq���c\��2ьQq��"�G�S���o�"�^IUl�ɠ���u�FR�lsޛ�Ql��:� Sx�>�>�6"o]rb���/���ÿ0�>�_p�>����]ͱ 'Rֽ�˾O����R��˺�'ELd��.�'60V�j��4	m�u��G/~e�C�~֏��