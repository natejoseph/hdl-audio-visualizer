��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X�-�����2�Aѐ��6���X�
P �2��@-+g�$�FQf��-,�.�lq�r�D��uәz��F�k�`���8W���k#�#3�׿'�4R��K�%�s��3�S�	��-� A����wުz��j6��]E�Y�Lhl�͔d��̈́�!���6�tT����$�d�g���}��F��x�o\��LN/���x��	��+�gvN��Mhor�`Z�P��*�:��U��ыΫ�;�j�Nf�`dϡ�lp���_�s~��a�ɮ�RG����v�QX��C4�}8���۞���Y�4�{X���^�VQ�MN��B���m�aڮ���,ñҾi%�v说�l���9��e��p4~���b˘v�p�=r� ��Ù<)�3��	[���M�Q�ą�dΌ�L���S��3�xAQcr��WYy�f<xN7u�@S����%z<��z^)Y'�d��1��a���e"�Ah"�n����Wf٢����d��6���{�	��[���֌1k���w#��	���� ׵�s3�e6��ny�Z��["9E�A��Âz	V����x�X��(�b�,e�Yy����Q`�whQ�I� }Lw��:�`��p�dl^4l6ݬ�>�o@�%m��۴>������춑jN`� �qz1m+�&Z?$�M�a�-��V/J}���~&��'�6��l�JJ(w�s�r���5���A�V>�r�Fs��˾�Y�*ӱY1��N���]X>|VÚI��ۛ����S3�c:T��"E� !�b���P$��cZ[��[cm�VZ���#��RxC/��`���T�ת�Pp�4��zGwB����J���3��y.�)���O~U�
2mܲ Â@�4���ٟ)!��A�m�Wk�m��M�+�Ǎ����(c�M�I����瀆�r���	Dd�t��Beҥʧ�L��N=@���ջM	z��р��>l����㐳ؼf��^TA��L���U���DE���K[��a~���I�ȭ��ʉ�w,�匸_<�aS�E���4 ?0��wM��3r���^=�������+SAU2q�x�Lt���㊧:< z4�l��c=��L�%̫�����VpN�p]w�����wZ�U� 8�!/>gO�l6��!c�sGML��؍���ƈ��{�[��@��{�Q7_����i�ؚf���A�U����K�L����4g����9\㮐��cg�����- ��1��q�9�I�/�s1�}��]�ߖ> H�Z�oH�L��ɓ4�T��#FTol�v	<kȇ2�,C}I{���o�E)�~�1Hə����@�B�H���v&�.�D�3���c>�m4�t����c��m�5G���вq�l�f�D�Yvz��,һ�Ӓ-�,^%��E�l���O[��"T�y�2�AQ�����?�l��k�����g�0�Mx�2�����WT�̋��3ʞC7���Δ�5��٤�`���.�����g�BUs�D�N'�ޔ>Qh��qh+���x�81��Ba�3��T��C� ����Jf�qRtFCS�ˍ�������75�d�����mx��`�Ԃ��d@� �遜 ˇ� �β.��UmSA�q��G�.�L�Ga9e�uu��ӷ!��eR��b
�=�
�ZԓU��"ϤdU���#$��{\K��;����A|<6�Ȍ1D �5������q�f,�w&D�ϱ�o�G쯍� ��TlH!bңN Qw|������{hQ������碣x�Ԣ?��F��Ȗ��a���Cd+��릁Jp�W~���K�����'�S(���f�H('[U}:�`�B�l4Z�f�g_�wi�?�q`�.;�_��	���{W(��O������Ihl��H����b&����8w%a��w���hNR���	M#�77A)Z��Mf;T����΁o�c��"�)�����X^$y�L�p��c�}0�H��e2���O:$���ғ�$� !�bf�n8��Z;�z��=�:w�2*�9y-<�'��ZR��=8O�t�o�9ac��J���E-NV��}&�T�p���ӓӠ"`���i�l�А�*]�- ��*Bũ,�Z�@" ��>_�'�:^)�L�{C��T�-�.gGG5_��80� <�W�%���G _;�d���dnѿT�w�b�z^�s�u����/��_�� �)�R�k��]��GTJ���߯�i����dS�h�ʓ�	Y���OI'���`&��7l�±?��ρލԝ:�F�k��͔��
��w�*�W��#׽��y���n��O��j7��
O��x�����x�����n�+'ZV�{�n�2<#/�	}v�V�tf��tzB��{����m�L߁T��{c�cY�6ѱ��Ŕ��s�$�x�#k6`ߒ�m�=[J�~���+w��94l��-Kyֶ�-Y�j�Mۓ����z^GL����.W��.�u�����1������^�@w���[u����(7Ea��DW�����%��"�O�7�	4z�"�9ڼ�)����8��ێb&k��hKS�Fy��h�{�h�.=�����|�o
dUq՟�t�fGE��K!ޡ:��Rp4��y�X�|��$>O��	FH9����2�5�~aM�#9����.���M59�AG��>{�~q�ӭ"_қ'�ݓ����L-@Z��yB��xZYc� } �Z�熚���I�.���Ito����QO�����d�;y-����vyD��Ha��8�����1�����H6(h���[z_���q�}�B��Q�o���!u�sV���a*ͨ&_;�e!Q�S��0���zT�X�J ���,�Da���&�& 	đ�<*�n2�b����CG%�x�p&����o�tx))$E(����3.T-��)Q��o�%1,*�hU���$R�[��5Ҩ��V^t~b��|�Eђ���4X�WS"��"�[��~3r���hS;�ʷŲτ���x�ѕ���T����,�=��#�ˠ�'�ʦq����gU} 2E��D��ņ�&dž��i��j--ms��4�ڕ9у���)K[�bϧ�R4���:���:�ɹR�z����L�� �z�V�k0�f&�nASQ�C:����O��1��/�(B���O��1ǤC�l�<��+�X=���O�F5����*Πcz��h}L�7)��3���K�)r���^!|�C�H"��g}�Q�Q�Bt��(��q,�����L��i���%+l^��'ƾ���=z،ƭﱦ�����^�����)�sb�M�O�3"+�����b�J2�D����0��2NV�N�(&�-I��t)��$�Q�"��=�D�_=������a0A��=���h�V�lx�F�̘b�Ѷw.���)Ľ�:?X��7��Z�R烯:���]��vBr����	Q:)��Y`o쬯��M�n�+��Z_���R��Zf&�����Ov�>�N=� ��+1�S�c� @���9	YD����?l�5ķL�E�1#�#Vٔ��7ÀN��	�|	�w��<.p�,Zp�F�J��X���&���/	����"QF��3���ʙ��q's��q'�ToNF����O���Ծ�ݚG*h�Kh
��{��nx)Gg(�@�"$l����Fޑ��~r�S!��;�%N�4���"W���Y*z�ь[��`��'��]b���d�!�"6f�.ڵ s�ݏ�����&Җ���Ԅ�\X{�o���q��G��C/q�O��1X�� ��z��n��f�:h�Lq����A�o�UϔńuY $ܚc{�/�9��p��9Z�)&�C
�y��SZH%���s�VwV�>�.�zFC�l��<���̓XF#O����� �z�t�yuZQ��i��9M
�|�,����O���2�]ȡI��5�4�OD�c�+��,vlH���-m����r�t�5|������ �
���z�fJgc���ԗ��^�!	A�(i�F�oG6���A�Ԡ|�3�8V8����na ��}��jo�qX�x�;f�=�[�K�� ��L�/,L��
��~�X����^P -�a����������-�����<���*��[��f�a��A��M��4x���1/Omla