��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�YO{��|+T����� ��9�jk>Q�5������3�+���Wv�X��u.�������|�[�}�QMvTB�űB�t+�%�B�����$�;�-Wŭ�L�R/�c��cu���jh�����Ѭ���_�<�@H{0��]iG,X����4S���$!�b1���B�ZE�i�\N�;6>@����j��L%�O����XVN ;���u�e{�P� R>�hi	��"��(cR�����R:�2-������u��(�3n�q'p���O��5٣U��&��w�1�E�;�(hi�$��V9ʒT
�i�KLx�ӡ:��9I�����+�U-��?�t�Wn�S;W���}O���s`�q@"�D߿�o����须�����n���[~�H�ȴh�^C����F3��U�t��/z��v��~ ��ĺ��)�-����u���j�'o�l�k�H��e�U����Lʚ����9%��h��}�z��:����Ο�$�d��b�4e�3�x1n�_�̄����#v��y���Y�ө���#0�=�'=��o�n�h)�8��IM�4�FͶ����M�3Ț���?Wa���-%�t#�p/7$�ؕ�����M�q�=�h2�9��Bڣ�%d���گ��Ò�rxK�qR۽�p�s���V�ӵէ�&�8�	�F#��i�ط5kc�:����O�՛��R��C�#��#v�kJ�3��d�C_:�t%�+�����P��G �pǤ�\��i��2�Ü�6!�l�݉���q��.�7���bb�����X�?OO�
�X$�WӔ�����i�!��.)xH*7 �ǯh�,tL�5�mZ��~�i��p^A\�5�l�ΐ�%;�맞N&���@xO��Z�[�(�WT�:ܸ6�!��X�?��Q2�u�f胘P-/V�����?����^�܀Z�'0�Fs�ׁ�L�i��L;�b-��ʤ���y�u���\��*dB͚��Wo����)�UZ��u�����K:u�1�"r&C��t5١[ʙ`�_G��t�*����M�lL����(M��S��h$�A4`L�c��Y���D�Qn�a�����`���)��q��xI <���:����?����璧��ֳ�%9~Y�a�ن�~��A�p�_@���v�5W�c�#�I��ӽ055y���KU:1��pdx�E���:і�1$h�����W<�ةd��Ì��	'��!������O �ѯw�Z
����l����H�d�����|�_F�.�9!&����N���J�5���gJ.,������eә1����o�W?��M�Lc�bZ�t`"Q֯���jh����}���x�&�u{@V�zML:7��G������!b�I�6I��z�T8����L�/5�S����D����N��4��L����g�ߊ�{����V{�^��i�W/�_)�Y?�W�6�B��,�?��Y�W.�ҿL��I�^�%����7Bu�D)iD���]NH�}�BX:,h�V4�n�6Όsm:b�3��h�+��/���M�� �H��L�FX�LZ��V������Z��,�w���N ��+)@�����U���-�1泈c��}8j�<��~u���l624���#����|��n�xWPŹI���d���y
3�Q���$R:����{T
�Pk�H�n݆t������r�Q��'�u��)���!� �?.�'i�mL+���j�:���vwo��Lu�O�Y���O���ì#��fd��M�U��J��􀥋�7�V���G�	Ǖ����s���Q V�\�d�<Y�*�d���L!��]{7�M�$�Q���m���`=f�1+�>�<-U�����.�;��g�Z�3�}�?ޒCU���"y��ح�������R4�N�i;��F�U�j��$>t�_�#౪j%�Z�hy���oT�/����y+�7+ ?���e<���I[����X�?%���U���b5���C�3�ג����h!�k��
��O
��}X�4�R�Ժ�����Iyd(���TO�Bw&Eq鋮�񝇥ނ����:��g;�XV�8��Ua[�_�3�
�-�~.�L�o[;\Ć�]���K��aapb�)�~
�C������	d���^��\�
���/�����'�["͘ ����R���jeW��z�@���@��q9"-�nx�f��R���4����N�����C�ɸ0�I9��iiI���d" �� �S �Nk���=�QR\�~��m?�S^� aD����>���3�rmÁ`l�7���˙Ę�6x�{�O��\��{/���ӄ'ǲ��ԍ�535�:r�ZGR=�-]���ӸJ�/IQܵs�O;Lˡْ�^'<��<���� ���PG����xi'������
ª�yWF�j1-`�+
A����6qJ�E����g��S����+`��J�/�WB�`���(�V��#��r>��n5@�fe@(p$���LIK�YU��,nM'aq�'�p7o�%}�:��I �<��<	���dQT.��8�ƨs�x��j�Ig
�~��
%s�QS��0X�bϓ&�/dy$Y��p
F��r`��c�B����<����4�1SrQ��:������)�N�X��u^���-4�p�e۳増���E��U�1�l"��-���-�m�۹���iE�&r�:<�+���r�m��4��,����9�7��K8���߹7�3<xL�����+$�v
��LP�)�;��� ��<O�p���~x�қ:Q���?��ȟUX�ϊ�~e������$���C���?��H�
�s'f)t�WSΩ"N��C�M�/��F�n�`,�w�C��\jF8�	lW5��U���ձqy�����=��C�S5�D#'n���"µ+��bd��B��I�'YG#w9�u_��)���igQ�Mqr>�����N��/1m��/!w�O<T(����^������>�<D�ɱK^��oJOj���Bk�����ߝ?�[P¯'�a��}�Q���n�2��� ��#R <�I�0>=w�&-�n�g�t*Is�5�c�$2+���ʚ��.G+]7���"2c_�����'y�dV�B�?LQQ��pl�����9p5��6B�ZҖ��9�����{tMN�_y	^����zq��%!c��@���H����}2���a���^�Sx������]�|d*d_��.��z�4�7��Z�|fǓ���jy,�*��ӥ� ��k�慺�2�)ZB=�`n)�AA~���0�ʆ�m���󆈮P��b�ҝ�<���oH�I��Ii�����	�������V> ��Ȏ����W��p���_��}���8��&���Z�� �4������`8��{�l�,�f;8M4z��F�q��U
��Iz0�+<'�J���k���#�9$��`��aâ"�*�zv2w�d?2��t�g)/�l�V
v`|�իN�.O���t�6����r��3�.��,hW}���tϘ��=��{��҄ �q���c/��/T�n#�%A�Ӽ�p���@�I��q+�~�<��!��D5U���1�/o���Ki�D\�Զ'įZ�=T�n)�8+�M����x��]b�jK9f7O�u�����
��~&GpZeڽ�Mı�P������Rk��J)�W�@I�U�t��p{�kCh1a��b�U�?ͫ�z\�� JEjaET�:�?=MVX� ���<H"f�e��	]?wU����\ݴ���
Oޟ.'N6�w��~��ˎqe��C���f��ҡ��5�9�De�l���7����^�����[����үvI�0����x���b���ʗ����TU����_��c8�Q��7���\qR���X�r����|j$�9�m�~F��,�� &�'x;���'}su��G�<R�pr$\�_�B�@v�}+���+�3Vk�A�|6dZ�Oҙ�47g�/`�;Ѧ<���	(sI�m/�����E�( �4�4#cH�
Sv�m���T�@~ۉ*����<̎���i"�����2��po�I�C�|c^��*��w5;��~�G�ĵ�)u_,9PWȳ��}�+��J�����`��1�P[���i�ҝ }��g}���3��G4�[D��ŵr�s͝Ӛ�6