��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N�����d纼��[�p��)I������_� �Ř�ͻ|I����#A$Z���W슥���'O��� 
�>E�y7��h�sR/1�m��dI�
!Gk�� ��?���c?�\UѲ�݁}�tN��9.��k�K*~�xRZMVZ�s��������s��^�/堀����t���v���k�h@!�cBb))υ�4�HV�0�3S��,4��FϋQ<iڷb�L�iČ�35Q�{2.*ݔ\�Z�-����'�J1�p�%V��Ʈ���L��!�C��Pd%�ӈq�Q|�gl-�]�dv�H����.}QEI|�A�&��ɟ�޳�a�zee���u�!eNp�<��W/��?����K蒦��CÕj�w��o��.v�g�[(KSU�������ƶ�E�VPwb�
Wi,�ؐ�6x�=e&Δz/���MT\g�7��ܿ���>T�EQ��/��x\9�;�8��8v�'�����ޏD�[�82��1�@����D�ށ\|���bw��BJD'�.��ARN�����<��{����<�6����a���t�1�a�����\`0I}����\B\��aCa��v1I�
�q���eTSE��_WAѩ���`Ɗr���9������/����a٬3*��?��q��>���� �K>m�7�%����YP��Ň~ȏ
]:�⊍���[ʦiE���t�ߓ2����hBiry���)������`�U���$D��B^�U��ߒ,[ݡH�B��c�Y9[��N2A��H	ٶI<�[�J��d^i�ƺ&bt�W.����\Xz]���[/�8)]�B�n�$�l)��	#.)�}j���|��N��o��I���:�蘔fl^ ��G#r��"��%2N�,T�3���=6�s[��vY�:�k�=&Aߎ�ĺ�^B"w�>3[$ݡ���f��@��W)� H��̥�����`%�̐�_���s�P?��gI�Ij�j3Vs� ��o�!|�}`z���?7^x�5;<��}d�J��KJa������_^&�?i��y�FGtC(F��J�l�!8	|O�#Ɠ!�a�˅�'.�M-��p`�gt� �6��x�?�׼����(���p�0�OF�Cu��p%�2)p$>��z�(	+���-�� �t�a�Cđ� �(h���w���&��C��'I��< I�Fc��'���6��Edm@��ik�8��[� 1������~p���z�'�.��L�ᄧ��i��&|1�e�CzX`�Έ���ƈ���x5�V���}�U�������r;�U���^*������b���AK6b{�N��;�9�c�V���d�O-��|$��K��w��@h�a���4�Z����l��f��k]b�k�a�"٣�+��v�rD�1,�w����4E>��GxW��*;�}WCZ��[M���(�J���j�������b��$6CEMlxyb��Z������z@8ǡ'=�~~Rn��\сE3�|M@��.�t�����K�|(@�7�O� �9�^ԁ��\cYc�d~N��F��E�*�&�;np�S׃�8�+l�oD����j/��)]Db�
����o���k,�ϔ GM)<0P��3�{ KNV����)1�MS�?ئ��}@�-�٭G�7���zP.Qq$��߁BQ���
�ba�l����rd0\}]�SC�j��� W��A�=c@���$�V�?��,�����k�5`PAz^5��
[�48��ܘL"/�)<h��Oux�8����e�Ȩ��s=/x�/��_��^s���X�m�ޕa ]�U�q�;p�f2�i�Řv�\���#^;������p�Ρ�8�.Ʒ\�M�J��e��Ҽ��d��,�L��`V�e�,����d>��"��C�6tp���ݕ�������e��'b�>�Nh
V����#H�:PK�Z�����:i�܂�/���c�F�P��'e*�z)�W�ؾʏ%0�j�3�F~�L��;a�g1h�%R������ɻ�"��s�[���5L
8���vaM2%���h_Y{����P�<��HɅ��H�e_�O��j:�o{��.G� ,�}�5�/��t=�1�������z"�������AL�Z\���,�@2c����z�:u�޻H����������w����_KG��*��W���$Y��כ���6f�5���D�q�d0�BqB���?����	���d�r�^�jdڔ���׾���sOǈ��Q۔ÒE���u�X�.�����ͣwrr���T�A�z��TQ<��;��2�maIb_!���ydɱ�q�l16�������w9��bU�R�[�Bc#0s�ܸ4=9�l�h2~��)-�u��i�M(���x#H�D�h�3R�n׻[��3��4ɼX�9t�&U`Dyޱ�*�$�Y-��L��?�ZO�����\q�f���F;��8_�Q)���lz!ݏ���f���N��� q+nȺ��/�.�ث��I�;�Dz7H8%��5�.�#JCS9��ŗ(pp�'Nˠ*�|L��5vʚ�ZQ}��6��G]�mP���쑾bI����}�Z��,���Yr�=���]���T�������Ě�K���S���o���C������(]y���m���&dig�OR\X�"}��Dc�U��uH��_�uE
�U�F��9 �4!�Ğ��o����)��V�����c��P.�+���:�^8XK�&M�@N^\� %�����i늟�7�^�D���=2%������g�fB�-�-=�:�lM$�e@ɓ�����8d؃���Y����?�|���VG�;7�D������I)�g���?��+Rr����&<e�t�V�Ƿ*[�@.��更��T��VDv�y���&px�1������[��p<�c+�DrQP���O�R���J��g0�q��ȣpki2e�8��^��8iЭ�͘O�/ޟ�E\x}�������A	�L��B�Y�--�Ez�l��"�	2����o���^����G�|iux��� �U>W�=U�������aŏ��Ea놬��R��o�I_��\q�l�W���P�Њ��%�:D�O�e��1�Z��eep����
#m�տt ʋwM'Ir�ON�4L<]��Xm�m�D���CR�A����;���N��7���Oڧ;"�J�8�H�z :z-�������h��P�-u���V�}l3��#���{q�0�J�<�e���g��-�ێ���v-*/g���Br�TD�q�G)���!�L������S-ԟ�'*��m&����������>U��d�)@��G�u9Zt�3���5�U �Z��	e�Iyýey�Dw���u��K�a��-�!��os�E�b	�L�J�ު{~˷\mu���<>_u��{c��M��O �כ['+5�CI/w}��:��Z`k]��-�J�>E���v��@�?u�`b�"���X�J��6��=����̽P!�Q�����-�w�ǐ�W�G�p�Z�+o���PP��Vc�')\w�p��S?�p=:�]Q)��<Q��5��È��F��5��J�Sc�.���w����(���(�����U�#��l>}IR�#+<8
z���,%rm�BPi�|$��'f/�ö�rǌC�(�4rG���;����]}�0�ڎ�iܢD��`N�����9�������R@�.q\mse�nh���Jw.rD���pp+�Ґ�_RP��ˤz.����|0�'��J�J�(����� S�?�0��'�G"�|5/,��^�h�2�����{5�t�:A�yq|�׭lu.��{`3w�'y�����\ O�t�	�\_b=�n��� �~�H}+�9BC�����x�����P�m��(���ܪz��@� +wq�*<J4�\/��ls��K�5Y�u��Oɟ5\Vg�s�ʟ�t.}���Ւ}�b(AI��3y_�������Ak�J�@���r�(O����#�O������#�M���c<8��U�rͪ)���$O^r������)��L'P��i&Z8t4�}n0�f���'�2�O%ʦ.�_�zX"sL��+��}��c�3�H??��J��+u"�*~P���co6���/�ى f�('\&w���D��.F�G�Oq���{c�f���|�&��U%�OnA���tQt)�/`ۚ�O��\4��|"�o�^���Tx��u0�3?-����R����`OWF�4w��a�T뻭X�kUO��7^fn�B�(6��^'���c��7Ed�=�l0M	�)z>��6Ad�;*=��֫a��(��Ϸi�aO���P��`�L�|Qk���"�R؂�q�|�ב��+���Ϧ�\���[��FΟ��˿�8$�N���b ���*�؂��D�Z�Ͷ�#��zTp�Y�����)9��O��Qă.��8��I��_7XU8!��F���^q_Mr?%�|6:��̑�5�N^-lY��Vq�;�ФEF[cREGx�pT�n��PC�
�]���C�|�
]u�C�f"��[���r�r:�V�9p,Vm�vEN���樱���"�`8?K�__��D�!�����X�-�;�A��9e�p��ȵG�L��Z��Nq��:j�լl��4�Gf=D���,z6!.(޾xv������{Ϟ�N�/�	�<��	"��<��$
"͕57������E�+c}Ca�O���.�%��:F�y�����!������hLm��z����?�7��*wR�.���w�_L�E:"2�w�G,�0��N��X-a��@ܳt|t��1 \5d��mB����A:*�b �ɵ�T�Iy����jd@����������e��(aE��o��H�����
��|�4\T�ޒop�B/#�"��Qd�Δ���?Z�Ѥ���cO��:v����u�^�b㜥	�e*�hI��.͍SR&�~��}M�f����fyx	�1�39�,V�������nD������«��Y�3Ӵr��)<E�y쫍}��O�G�%���դbXLg�������m?P�+s�^����Ww7 ��g�>f �/P�	�Ƙ@�/��!�t�GJ�C+w�MW©�Zo0���䄜�qy����k���q��l\�R!�s.�~��_F���_rK'?r[�5s��JeRC�#A6�����m�m �Ĳdk+�z7y��}MƄ��`��Ps�we`���N�۫�LƗfz�A��M����и]�m0O�Ă�OZq�r��[�9h�@�T{�;CV�gT࿋o�L����cpaZ�z�Tj�A���c�o=Mj]y�1�#]�?s�YX��HV�,�%T҆��[bJ��M�1ɋlG���V*�)�����6�Cn�ɀz/b��Ex�ϢlHI��:�^l�`�"#��WT��-K�,@��#��-`;����MY�?�c&VҴ�u��}NF���"t�;W<ֻ�_W�� ^Ɩ�MJ�ey�	'�a����}LF�j�ֳ��a(��b�su�ق����E���}q�-7�����ઝ��Z����:��[&34ux�Ȱv�?ؗ7��#Y�us��b�I�BXҩ��v�IY���~4=�g����\=w� �*cw�~8�W������|8�����Lm�&��^!|�(ioi��oe|��WǺ�,/������Kym:,e1:21���7>ȍ
z���w�'~7����4��Hutz׈�G�:��tB��T�UG��Z��fUSS�-@���杔��w6��8�k�GS�W:�Xdُ��Ȱ��o@��j�Q	V@���-vO��(��d;�Ȭ}b�kK�+VH�C����Pa�*霖Pl�q��Ax�����!@�;�~٥�3w�pz�J���f9�ͯ2K��xۡ���s��NU0���7ppx���Gv�BY�ɵ�+\�U�v�!?��!��]7��S���������"de��ƅ�U�(���j��1q���~}/N���"Co"�#?B͒zm�j�LV���i�^��j�L1Ȱ��Y� �el@]5�K��:�墌��vq���!����t�
���nC
xއ���)��"Q��@��
u��t�%v}g�'���x�?��:���d���ײjё�'���%����CG-�a#㗂�'�J=Lޠ)�6�d���i�,L����ܤW�E�Ƚ�����.\��NF�뙧�>�H|�གྷlѺKg�H� ѾoL4F85�����@#�T��� Uܰ���7ފrXH|^��I*�y��w��4�D�=#p������HXz����&�r4�Y3��O���Pb�9�&�1�gag��o�o*���i{�R	�}�Cpo�Z��^XĨ����
,�p�q"�J�^kQ����^����\�7����@׼s]&��ҏN/��d�u�bBF��z4,�*��m�=��1�?�d��/��S����h�qۇ�4��	��.$�����,��sp(/�M#������)��F&��l=&�3��@���EkI� �Z{���w�URR@�T�.���W����6K��RY4��c�[�g�+|�"r#��==p�%���&��V4��4?�.����������Y�98z�u"$�I�ǫ'Z�խ9q���A�3H�w�6�(E�� �}��w��n�}j��_�wC��\�xDϪ�;u�B�&F-=^ 7��`vC��`�NQnI/95����`e˹+=���r�6��U!H��F`���E-�Ŵ����'�e~Uԇ�-�B�1�R����!�uf5{�?���n/N�d'�?�-p��u�tH
���j��O]��>��'5���X�k�b�
%i�*�G��.�;>�g���7�K�ʵmJ���"0eǛ�Hq�b�ݖ6���Jƚ1�s��e
H�{�,<ܪ|{G��@T�'��O�l���j��V/�3U���]w���$��F
�e~��g8� h��:�T4s^bK��K.��38�ԉ[��vތ-�3E�x��$*��wnF|0� g�,L���%�����ٴU�E�AOp,���<�d�\*�r�)�{p��ec�� ���o� �n�������&���8��<9�q��Zʦq���m0�3������PJC��x�4!�t���z��w��#5�\T;i�[�M�*�Zq�N����Q��� �h fr�KL��I3��v�J#��9�0C�+��C���K�����N�a����yB�s���U=S�j�џӑZ0N_NF�+�wz�{�p#��㾨!w䡃����̈���V �x]3>��.�S�UH_��ʨ����+���R��0�XX�{/�����;�+Z��ӕ������ܴ��#���x��8��mf�!Zbw��7��4��h��lm�_��!{��ȲjF6�o��H%�]�	+�e��R�Wݡg���E��H�'�s1��Y���g ����tDH����;Ͽ!���l>n�ļ(�����t#�}���G��h�|DoUy4�9 ��x�g,@��^��6S��x��[�N�:�uleVmM�턮44�ݼs�K�u�V�0�YV7�%1�6ߡ���\�1���΢����.��3Pꃴy��~��(˱.zC�n�F�N��.D��]S�z25�)���D�,���7����.�0�>�:E�pVͶ�\y��Iˣu.�JB��������I�{W  �����u�ӨK��XGr�����O]�5�ͳt�BC�~��&L� ��Z�VT���{p�Y�A����Q�at�K�?���J��I���"b� /oļ̱�!.��R&�h��/�|���$�$�!1�|�֍�V�����Wԝ��[9��Vְ�b�|Pb�G��ԏ�vEl:z�q�(�|��G�p&(28\P��c*'8�`1<�*�v��qի�x���~2�U���A�4�QSm|��z��ങ�bD�]�js��\��P��k���v���0u�LV�Sl!4����u�> C���x�
ҝMx�X��� ��1Z���H`�0έ'm�����NP�\@��Ҽt���XTF��3�����d��{%��d�y�^�KA�I�?��L�h�I�R���W��'!V����=�����X����,׈��?�X��у���ھ�@CJxXކ���K�P�(��Mմ�J�4+�J~�v����<w�尤ì!���_qW���TN�ǡD��\H�H���2#�2�?�a^B���X�M! ݐoFV~+)V����|�?�V�:�Nl�Q�|���g}��������R�O!����u�L��=\�n�o�`E�Jy�Y��0t�xYe׌L��)��7	���|smr�<{��-����$k������]i�9W�!y���U�wTW�G��$����i�`zw��gA:�l�&#3����/�T����=AB�J��p	��z,����g���/���Ǳ��Mf�M� _�ھK O�`�=�YmZ�=�K�� �|ð�I�sIi-O����g�kL���ߧ��\����S�ZN�)v�� 1�CݑHo�/{�=�I״WP�9��!�~�[쩐��r&Ol/�]t��c��g��p7ӡ���nW�v�nW��ht'��0|�#*�I3��$�e�<'��ݤ��b�e����p�Ş,����4$���7�ˢ#%�M�����W�K��C@�UIF�\o���6�W�4
ӯ�<���p�n� ѐ�yB�U�������x;����5�&H�cT��FV�А<إA�)ۅ(��]> ɥ^�m���}��p�L���W�ϔx`�>����I`
�,�$��K�i���N���SY�m;<XCO�Q�j�oAG|W�ѻ�-v���� ����t�q�)D@����U\����|�kB,�� �b�����Ouj����0f|;��|r�$���'�����vY��$e�-7;�5:DB]�����Mnngӡ�l�*�R����;d��T4�o!q�@_v6ZT���2{��������k�`噬�d��l�sl�&M�����@]mF��ZTz�O⃘5�P�셪S�&�䧎t�;‿Yu�sm[*0�s�H�a ���׫B��K�X�@����S�˾iv��Bx�!b�*�-S_���-3��ѥ�:�_͆G�,·j �[�����I���;��6k��-{��iF}�W(tZeVsxp��&�(�`;��s{+��_���"Dȝkئ�B����5��
N�̼��i����ӵ�(�V��۪MC0R��'��[�B�&<\�N����C>6A������g&����F[(Fc�e_H�K�Z� `�hL��0U/�/�b�_%q�o���9��ɐ���Q�!��+$���Z�GG�H��/�!�.�5[z�GI�ܿ����9��s���̠����A�?3���s���
��}!b<����a��3_#��dy(�b�tX�ޣ�!�êd��M2m76 �7X��I'�0/��Y*�7�������$(��80+џۯ���]2(��LL?g�p���EɊ�^,��~�tl��'����1<���R?L�8��Y��	�9�;(Yh)�*	H�h/d�����JM;���؁�Ej%X%d���}[}�^�Y۞�ʋ!��g(�vKS%�}|�Ouqp��6L�aD�/�)IyT^�^�7A�/29bT櫙�ջ�?gD�{"{��9N�Ā3 ��B�42xUN_�g����F�\�jB����6�Ą'-A,t~���f��K��K��i�::P�2GvX��~Oj;^W$H;�d����Nqd��S�\�ե񳂟-	��pmSq��<�ߢ�Sie�_�$��݃J��W^�6�62��m�B�����ߤO���Y�y<
���rw��G&_ᬻ�M�����KW�"�!��w��&G��j���3Q��)�r���uV�����@��!@GŒ�X�=k�_���ύ����E�~$�e[��%k�jғa���� �䓤1�z��n�/.R_��S͞�4$V~3d� n��F��^�@�<�n�C���c�j��x���X�z�W��T�J�S����2��g'&�?�N�?2���;�����an���+�cl/^��ltl�`7��s�hp�����������s䑭��{%*$<n�ewbc��L�a�4��O�OH�pk�z>�*eSS����%5'�^(v�M�'��3��eV+Gʹ�,��jf�� ���W��:`f)ϋ$G��ܹ <�3V�䞹�~���l������:|]�/�U�Y�j3��*�ĥ:�`�R�����N�kzÂc��x�Sh�ڶ0�s�Rځ)�B���䴵p
,T9��~!�&o���+���)��������`?�c��h1��}_�r�Q��HR��}��Ս��E,�"����[����x����'�0��z��jϏ�%�L�����P�Ք�w�����wi���T���`���w�Ov���v
y�|v�����7OT=�t%�T�_�C+}�L�C]T����$5�ٯ�����.nѣ��J���B�U�[��f����^�c�$
�LmIS}+m����hn�(4�O9�.lC�00��s$w79Õ	�����|��c{ykA�F��	���Y2����s�J���#Ӈ���N�s�")""A2�BC ������OD�\�v��ZY�!�7��7�#"���'��1�q˛�2�$h0Tv'F���)䊺;������Ǩj��=�� �ؗ=s�<'�:�M�7�@{���m�w�1�T�@ZX���[,�R��;��B+���{,�W	ώ�G�<%�u+��YA�W%���e��F�o_��&��=)�;;1by�!��d���W�v�͆���&����W^�㔭KXޒH���$h�$1D������^��8$��͟���ך6�|>?n��$��H1^~c��i�H۪����D�Z��^��op���<��o����L�T��F����D��n���5H�اV�ӏX�DZ?ຢ�J{r��n�[��f��D�!V[ŗ��S�c�:&9�Q'�1D�l��'�[���(��E_�^�`s��u�����Mq��E���y -��<��K��n@����h�6ֻw�� �?ͯ�w+ j�N��E�(��g�pP;�ť�<*Bt��Ø��'_��
m�D��C��-4A����;Wy
���w���|g�ۯ���Ea��ɻ�uh֍��h�k�I��16���
l�_[qT��2��o��qp��i,_x�������.������s��xj*�}\"�1����'0�Dq��ha�dZ\�)mҹ(�=�hi��v0��F��H=$���s�0+�m��]B��}�Z�x���X0���S㝄���;�!c�|%7cf�#L��:��� s|=�RW/Tn���Ѯ�h��[	B$[^��_M���;�BS�ˏ;0�4\����XTyY��]Ez��U~��|�������v�x`�m
�X�^����q{aێ���w(Fc���� ְ��6/��G�KR�X�@��g�n{��ؘ��*�	��r<��H�C�\�59��,�.��Y����5�s��!����'��u�s���UKj��sg\����*��6n|�I����O]+z��O7H��Ģ�2;��s�)�$���� $��G$>�TV!�=_9gyn�X����غz���k�w�y�v�r/a�ў+f����*+x�6����ɿ%{ֆZ��x �MÑ����]ۡ��o=:���tk��R�+� �l��CQJ���-�@�x���n�l��Ԓ�����[�+iK�,�'�Pm�sQ$�v`M�J_h^�Gi���O5��Iٜ�~L��C �60O��'�Aåu����$P#	��5js��h���{􌷬\��J�[�O
��L@Q��̳�|Gn�J�<�ゟ�������F%���G������,"X���5���ж�!ц�?��!�Q�t勊��7m0��)ʨk&�\��nހ���~w�&�\+l"�!gMI ��sa��<3��������l�xL�w��%`b{���-DVY�ǒb��J���KM1!G�paI�M����c�~&̈�#u!�UU��߉���R� +�i����y�W	�*W��3�c8��8�3�$˗̌HƇ�&g�%o��AU<���"qEً��(yu[0���ɦ��j��	&T�ɫ�a���n�$X����!��B���1{fi��{2���NZ�ap0.�Ԃ��{5̼�_���3ʓ�}�<�,Ș�G���԰��eN�=�Q�a��`��C_�o���c�O��|$�q�o5�`����z6XY�^>��ov'�xG�0�NZ���J1C]�2u�&��}5i ��M�����d}o�����WZ��[ ��̠%FX�7���=�}^���J����30���ml�B5��t�	b}�nF��V�ŋ�ʫR�B+�[�oG;�帳�Kb������\�����\��嬹�D�cc����:�IDJb働�����B��mn���?y$��K�m}N���炋w�#�����Au�b8��3���(Lb���Z�FY��q�Ɵ�D��Y1����M��[D݄����e����W�t�h�uR�6�m���R�9��9�(1il�A�P�N�`�Ze�Ng*�5dy�l�����ۥ��K�1g1�y�'�x$��� c}35f��
T����c\��"��z���b�[����&72�����e�rw�1�MS��������0:�	��.D | 4˻Mj����g�V���2��s�K 9�F�L��������#�5��rAW��w��~��-�Q�2@9�7�>��QcH�4��z*4ܴy�u�/V�]L|��Q��o��Ө��n�^��,�=��N��-���AO($�qл:����P����CT�~}�[qg8ޏ��<ʑ$p�t�lV�����K��� �)˹KK%����v9i�E_	L�B;P��'1=+�"F��"e�uW;�Tz.�̟&��;��E� O�	mE�����J3|���{��]BQp�.>I	��i�Rz�S	|�����"ҋ�>�@�ճ�L�!���o���.ߍ��F��3�V�Ey;A�a�EP��D�9\^&\�t=\�N8�=S�1��0��ʣ��1u5��ȇfG!/Zt;?I�J*�⨻�-�R{�	�t� ;U?��P�ĩv|!Ka�ͪ��"̆E�r�Y�n�RP��� *�����X��ՙ4�D[=�q'�g�z���F9.w�=b�"�/�{d�{�>K	�'�qr�t�D[e�����8L�y��M�����v���j���EߌhV�>v���LJ����T��$t�M]e���Md�z�zz�u��}>
�]؏IwA� 63��M
"��0�W�u��k&cӿ�����i=��
��v-�<�8��������`:����%��|���Wz���'�=��O�,mt�V|�ɯ=�B���]W��Jq\ ��m ��0�q�k �-p�C��|^��� ���K��a�Ix������X5�:z�݂H��B�����f�����o�>��,h�����5�{\���]� �M�v�$+^�ɐ��R���/�W M���	��Z~>�4��&����V҅P�.\��R�W��xJ�J��k�̲ը��,L/��Ϸ`��EsI;�rc��m���F�D%�=׫��k�Sq)���Ad��Ñ���ϗ2�y6��1��C�	�+)��?'E˛Y�3��OW8v���1?��. e7�A�c�nLGi?#t����y3�t|~P�����@K�<U��´ḛ�D���g啕2IR���=��`�["����,/���(�j䇑2�\}P�q�;e�tmR=(��_E�.X�n[�}(�N\g�K�8�]�q_��M�֪W��YN��U���'"ŔYl�T'���}�`��\�L��R���3�w�46`��s.xU��n/8���*nko���.���R�뼚�n�a� {`Q�>�>���V��_���ۂ�]+��x����G�*�VNS��8�6�@��B�8���J(B�"�ԋ ��������0Ue�O�ȑ��zyqK"ěTTS��6�F?�q�Z��+:���2E#?�����ov��CQ¶�st�~Ŋ�iUAۘ����V��K�.�;+{���S~�.���u�ԍ��7�o�V����+&��=���F�+,G6LsTtF��Q�,��d�~��g��H5���w����F[���o�J�	�;�i��S���%ƼgM�:PCM��A�N����Z����>�̀�7V�6�H�_��J@���~�-�`�y'J�A)
��{͜�ʓ�2K3sD�_4�<���N�L���'�;��F�&;,�sy��z�Y�@�4���H�Sr��C�V��	�E��x���B?uu���@���J�w��+�F�2u���P�/���-m��E_��)��P�G�J;�^��uCo�#�~HFk[�*���_��ܵ�r-qq���)��c)*T a�_�5x��z9��\%/���¸���hQ�yȖ �	ȩܴ���mJ�D���m�����֐���$\b����M� �!J]�G�r�I!���[^k�C:z���ݷ�H|l��u@�����C��U)��]4%~VE�h\�V��j���:��c�w۟h�řD����e�*�<8������S�$F،��|��rY� bs�����yڦ�i���$\�wŪ@�Z!��&8IX&C?\�����%�8̆�^g������q~�߮I�H�tN�����qQ�H�� -KV9Ϻu�ed����\e��2_̠V���=����,�8��f������V�j-ׁ����K��\���	Wf�1y몜n�����Ti:ΐ���Ompؔ�t@����7'�J����P���dU���̓���@ijQ�fYE�9 �r��&J�r�A�&�T�K��H���u_�B�+��dx��n}�QId�ͳ���r ��v�}.;�\����e5<)���O>r��Pi0��]W�nU(q��()�R^d�i+8Zx2�s �����>xv�Ę@�j-�!f���a��ew�|�q#\ڥ2�zavN�7�#:��;�����e�������9�e���Oa����]�2�>y�wg��E��k�қ�;`����6$-��!b��{��4�X�$zG�t��e��sT�_�"݌["p53-ǰ�i༯ H.guC��}����`��@�8��r��L����̞D�\a��Z�ZתZ�c�����Sm�����Gd#ԡ�y���(z|��	T6�4dm�d�]Y�s�w��J�AF0s�n�N�!	�*\d��/3]��& ��[b��ǲ�i��#��	����-%�@g�������8S¡�6�$��{����0��S�*���󄨪�D��ɓO�����6x=U����ZiJ�$�0�6utt����M�>a�bߡ�TcYT�i�Zhu��0���2�k�(]�IzH����y6�>��_�RG���uZ�w+b�A��3�Vk��h�C�ᖾ� �_6J{2H��~�>��X�e7~>�h2�k=�N��%��-Y���ϜnS��V.jBz��7͎H��T��a���3g��l`����0��E�ķ���UA��&	����q�欙���s]������ u	�lTGEs�N�(�2`M?����l�J:Q~]�M�62�o����M�
���\��i5�[Z�7�^ŋW7'���KN�Y> `T�Ԕj}�R��� �<��5�{�nc7R��2��-����1WV��L#��(�Mĳ�����REyI7��4j������Ķ�C.
��oPH>�z�F[�!s��{�Q��9��O�"g��ؼ�n���=�I|�ܑ��8��,����[�m�'���q}�)Xm\R��k�n���~�
C+#�Ƨ,�|��[^�l���i��;�)��e%�4����_9`;4�i�H=9}(!Ò)��]1��WyW���^H�I9�2n����-&
�ՔcGhLyu{N�>@I��浏I2"%�L2�
����j���9֊a��g���_���e�Uy��%�x�ۻ%%���g��r���%]�e�E���/��Ïoi��Ō�� p�"�����aߋo��~Gi�}�*pd�"��Z�3II���� Y�|��q' �֌H��[.q�m�6O-����/�0�֨ز���G��]���J9 �r�j&�	���S�]�5R[�Ț�I#4h��@;u9Xw�����_ߧ�5
t0�Q�J<�϶8^�.�j�H�UV�r�wV���ӄk~�w�m���X���=�jb��w��k�� �-�
�OF5��{`����5xBk���]����`M�_=\C-i8���x("�#:^�6O����lsiGm�U(�~5�fk�{1,]s�I���WhD�ڬ� h����I���,#r{��~���,
�L(�T�����'�g�C#��`��ϡt�w�rFD�������Y�S����.5bȘ9���LӸ��FQ0	�����i�ܟ���yZ�L�=�t7�(�f�XM���X{�O�Q�)h2&�!)�B2'��]]��D���/�yL�A`��^�J�A��tJW�������U}�@��t���p����T^���}ko�F]�xF�"x͕��M��n�Y�Ь���˳� 's�w�n�(�ӴK��"T�~�_W��K��X��)�����b��+d�>y/�0���0{��0��o��( 渠GP`�`�}]ɓI���5�̴p��<�Y�8��vf��\�?h+�3����2pN�]������� � ~"|�J���0m@q(�;���*�e����������/�8�gd�y�6 e����09-!��X?�ަ8�R��Z�:i*��I�c�a�5w����&��}!��gbsm8*�*D"�̧�]�ӊ��S_N�F��b�G�����0=ײ�}g7�w��Mq�^ed��r�`�b����� ��������5-�Q]ώ.��l���0BߗD�hA�R�?+��t!��Z��s,���o�xxO�Y?6霿Ԑ1+Hh��9�!
5�6n�L�*^��3
����+ɻ*������� '�~����H�Øk��J`Ns-V7\���(JmRv��K�Y���A��)����o		h�O�	xek�a����5�y�?'?B��G��q��~t�Ѣ��V=*���'���X^l�哅��-����7 ���C������7W�b��Oz}��RiIđ%r>,5a�UA(�h�'�S��:��
�^ �lحpv}:4����!��(�|yܰ/�V��z.D=_�=e6t�o���
+jXWl�cL�I�é<
���#ݼLAM賨{�NjV��C8�TG��6,|A��W�P(��_�
Mc,LF��%쌲��6�ݔڈw�3��z3���@����?5
W��KmS>��S��z0�i��S��=�!���yHAc�=�d&i�;�ЀS��.i����Zq�Z�3�οg7V�-���i��u�MC��p�ӄ\��-|Β>R�A@H�v1�{m\��F	�\�¢��<p%�#0���g;������,���6���0R|�d���q�!:�0N�y���Ot+�}�&��5y�d�8�9-ϡ9Y�j�^��k��}����N���ʈI�Әv��.,O-���J�Ѻ� O��_}��J�eU��ki>����&_�t4�%�p�g[;����ͣ���~$�/�M�.�dP����+p��]�J�t!���CiI�GC&��D4�m�1�L�ad��& Y�T??�uB��D�e1|9��js���8�dFH�f���g�tL�QP/�mBZ�o�r�M%�hl��;�BJpkׄ��5r>`��G���yi5�cE 4��7�֒n�:��(- 7w��^�@�<�lTo��9����s��{�����w�|�	;.�m!�9|�����d��I=��yK�qJ�r��zaC���Sq��Cy�X���t�e��\|7��WH� �V�O�ݭL]�!f��q�U����u� ���������fǭٖ��M����/�20��u~���9
��:��蝊�(�U�J�^��ө�B�A�JJ"����g=D.����3��B�"l������Ps��5A���Wv�8ɘ�)�AaM�8���B�������x�1N�p 	~o9@���^��@�������R'���F.�&��nCOV�8�|7$%0˓-z$�?B$P��b�}�a�*LpTÉ|j��l%04�;�Y���ىD�7���O7C�5�U�;Qhm�j���Ge����-^(���3i�1�l*�tѲ�$����Hlw����*]C�>�R�Z��T��j-�&�]�sKՋS%��Ef�"C�b�� ��,Ksp����wH��Z��ߊ�؃mb��������~~���ի�n�=DR��B�o��W	��3GJJ�{z�2°v/����zP%2�C+�x��Wc(�O�!������m�ek�y *7(M
X0H3��$�ȡ��q�:�C���u7xܤF%��';���N)'�ľ{�ST}�N��&�G�W����ta�Q�.1Ü9��АT�@������q�̗�\���@���矡�X-�:6k��HJI��٬��-��XJ+6��C��V
vn����O�"E��z;+�'�b�W�&�Z(/r�Y�I��t̉a�\�9*J��$��"7:2��cEn���hdK��Yр���R�|�]��)q�g�N�je*��������`�R�#��/�b�{�O4��&�ދ���B�{�DT�����_�Q�'P���T���#G�Xd��-��ȤԘ�A�-�mgq�d?�[��w�,1RW14���ܻ`��eA.4"�9���
�F��jq鋹��`X��ѫ�	1b����x�5j0i1y�43���g��mz����K�R[�����n����Íj���ɤ$����Y?}�uhF�|�Z�d�z:ȧO2��dk���T�������
C� 2�5.���! {���U}���(�M֔8�"���UYbk�,�w����y��ôB0�\y�u��;��s�A�8��	����7^-�b��=�:,x'Vh7���r��
w�J���U��0�ǡYR� G�չ==�7�����*J��09kif��"��3�i��MLH�e�-����s���� ��WwV������tw2��蠼��z��5u�x��(�磅X�S���Z��C��/@�j�#�N'RxI�Q���"<u�0�0�����>�&��2I�<���*�o�_��\8^�:���p�aI�ķM���Tǵ M,n�$f���.���赚�	 ���T��*c>r���giE��XӅ��3�Uu�WY�Y�,\R�����K�B�_(^,t�z���3�n�\}�OA�p%=��}`ڜ�B/�ǐ�kϛSh�Kڷ��=�-9rC�	�<G3��hB��Q{鈫J��r0M�"}����I��4C;;����"x�v&��c,|��9�m�5yn�I=�*��jʣ��*���J2��ǁ�O�r(�A��o�DO^��-e����}�_���������R��8��dإ�0�@�ǥ���;��a'tNF�Gt�.�lpo��N�)���ߡ���5�� �]`�JT�F���+����R��[�O$n��;�>*ͺ��ݽ[S�3	��$�d�u�.�)���iq@r���޾SR�v|� :�A����!��M��U|�ͱ������G	��FVUE�(h;�YYV�z�א��h�p"�,0v��	��g-;v.���D�\��H�0R!����?�)-���'A@f TUy@��[����)Cr"��ԃ�*,�K����0z���}2+��7�΀�Ș��4-3Ӟ�W��|a�"L�Ѽ��<zh�h	J�����ќQsP�%�i�c-,I�8o��f�M��O�)�d����m~�6����1�-Zt���bnqӤ$�H�8+Ώ�Х�*(_�b�p�^�?��B�m�-���B�]�X�e
y[�TV���k6���0�Yv"Ɖ��(�ˊ���J��Y�o#��Vl/K����<�q�!"�X Hc���-�w�^Ç��������ī0�fO"#*�œ�K�C�O��u*l^	X�
����y�
�e,V"��m��1����9=J�x�İ�8P�u,�U ���}���j�3����P�b�lt�*3�.O��,Qԩ�v"�8Ȑ�^pt�y%Z���ic�_�AW�`��[D�d��w��cj{ip�^N���?��"qk]n"@���η���}�������O�on��?�im���`Ƅ1��+�oC�$���N�-������a% ����kFʹʱҚZH�;��V�i�������3M�G���75�HS�}@���)-'���6)A����>��M)-�χ�\.�9t�s��;9�|��O X��@��'�L���+~~ G9O*]� )��	�0��۶M�fd,āC𞵚2K�@	�)[۔H����vȯ���0f�Oc1˂��wR�=/I�'��D�/�J,�H�NR�ѷW�r���������͑ ���ܡ��Ms��o^}#�b�(�	����A��rK1�v�߄F��_��6S���K��p$H	�Ӱ�v�Ow�ʸ~&D|���$�X-��b�<�QUu���� Qу�Qk�����v�:�����<��[�r/�LR�_�LUk0���`̒� l������U�Ӎ���q�r%�^� ��@�s�H[@���$��%� ��s���]g)�D=�U�Zq�	0����X�=;2p{<��.�G��՛��z�i��n!=�U����8P��Rޑ:ŉ��	��>,�a�CE0W�*����Ӭ�}�zRh$4��aF��cH���G�r��A��z0���ST�V3u��;�i��p��Ѩ����[���=��%}�B~K��e�V%:�I�k�N���!MJ_�쟰��8Ea�z���i
k�$�*'(
٧�q�Gx&K�lJ!S~�x���%�ʖ��G��\�5����[���,Wi�Y} "c,���0\��w���"��zF��,hu^ r�e=�+rp���OF 
����`���_�m4s�W�4�T�G����;���M�>:!�<��b�|n͡L�i�%��*���ҌL���=�Tm������M�	�W�xdEJ�ņ5/�D�:	-5���~k;0@����N�S8?͜�OZ	��E�;n)�\5�xX)o.@�h�"C�s�jf=d�b�.�x�a�¹zK�渧J�[2O�!���Z#�%S�ȧ�7	c��v1��(��b��Q;�9�R0�1��iD�l�$3W�3����2��-NT�����%�F\
�4��s���_��M�?(Y���oC�<�~��՛c*���� ��;YO�cg��
�Ry{?t�����	��;�,���I�����H៳X�x��C/	�%8m�D7�*@��4��}Y~/xy�񤹘��g�*�}���L�Ӑ��TFVd��T7��{�P�A��X�}g y���t��Ǽ�ء����I��.�{Ӯ���h\ɕ���"���c�v�o'<�=)�u�Í�����XF.����BLu����B��QK�ƺǞx�4m�I�Lϝ! EG�J�\h}Ij�жq��>wO�\5��on�=�d��;�L�!�{W��� ���`��kGP^ʂu����Y��*�o�P���G܄;��O �~�wVhR��H�Ҡ,�z��-w��N����-+BF9����O�謾���Fc؆�Lr���M��E�}Өn�l��*|����◊��x`�>(9��}�訛�lK'��߀*�8HS+��x��B�T�.�p 3}U&�g{	XW�8�Xxɲ��z��+C��>��b�v���I�=�T�P�����DhЏw���9���v�#U{��El��k&
1�7i7�f�E|�|A��p�T��aJQf�?<J�<��S���T\�p���Tuq��W]�{s:N�Ya �B<��^-c�2���w�ь��Fb�ߥ���LjWf���ő�~]�"tS{7��E�PImP��mǵ�w��]���sq��*��K�0gv	�˨-��Y������'��0���r�7�R�6�S�ԁl��R}hI�[� ����w�%yv��}�Q����$b����^7qA̩L��P��s������5�P���s{Ԁ}X����4��o���P�e��t`βm�)�W�_�K��D]u%;�3}6U�8���7W�$Su�
�/$!;�Apޅm�>��"3 �[�8��m���a�n.�jS�J��a�
=�� A0t�ͅ{��
�Ƹ;�y� ͥ�O���-��!AO�ۑ�34�M��ZO�é/-�EI�/�˒b`FG��  �>h�B�y�/#��pJ�VW�g��~c��1+d5�`�V������.P��Rt�GL�j����R׻Օ=�9@�31B�)�L�s���j�����
`Kls 6b�y���t���<M�E	��~�d�i���`6�͈T����*���槨Kvy���}'\��)���k--�'B� ��w��aAq+mXr�������-[�B�_�2o��~��u)�t��I��T�N�3�l�d#)��+����4�wBw�L�^�v^�;����|�L��� \�����7�˹��ߏ���v��+-�B�O���(l $���%�֚�a��cm�[=qy1�Y�����S��#f�����x��7�E[B}Y��5d���ы*.Q ���*(��G0ƵD���o��y���Χ0�#� HuA�I�`����"��e�c���J�c��^�Q����bC���[|��3�,}�#Z�$�蓮�|T3�3�H��������8Ր����|`=��������C�L��Q[�	v�{��˶���K�c
��N<H'j&�Fl�F%>�y����p�FE�'+���Q:nAV�?����������Pe�@�%ΰE�# ��1����CK��O�Y����j ���@�f4�;{˴����+	�'�x#	 
���`J��Ht��v���w�%<�A�h����&x�I���M��`�=��T֦����wmt"	�.�v��GA�}�G�V�dODA\�a!0���k� �w ��������dP6ƛd$�OS��ƴ�Y��1�o����uIk*J��$E�,�e,o�$OFB�?�=���
��4�fi+:���HC��=Mq!�mҢO��	�V��pt|����SAs����3�N0U�y2�S���b����a/;�v�7h��LҴ�Tj�N�a�@Lg��e9_M""z��1�QOo�� ���<������o��r5y��TÙ$|�G�uBh
�*8�����=�s�:|�Y�a-��ùh_K~�nd=&�+�_����pM���LDV<_n1�駑���F�����Uc�e���!�����.�*
w��m�6�"���vP0�ڤB�8?Q?�JZ��B|�_����*I4������6x`@�b�mmL��K��Wg/,��XN���_��@C�B˭P��æ�5B������.:���Tm��9PL��ƛ<��G{��SH�����E1���?�Aݖ�S��<��	i�˄��B����>�e�$��7~�~����vg5hڬ¢z��|��WT8J�|
,���9�?E�g^V7!ǭ�$JO��\�S�c�2��T<2�5���}���J���啕2#��F�f�(`���S��nc�axg�'�e��.𻵚7��ļ���X��i��0�p�i�k�緩��_P��Ѧ&��M�F��+�!�����& WT�)z���3DOS�BEy�z�Xƿ*�r X�� ��S���ͥf"h\�s��2�؄�#�`4T.f��ߤ/�������u:ĥoڙ��Zh� ��j�T��"��o9I��˝\S�o3�M���!�V��8o��|l��z�,�t�9��k(`Ccj;�F,f�3mݷ�p��M��dO�}�
\���r'�(����%����ߴQlܚ.�_���YM�.�e�j1���#�������>���;�+Y�ēLG��:�`��NQ�Ȁ�{�o�qܩ�rƌ�z���5����1e�22��S��q�8oZ����*�hci��Pa�^���gf4�!u:�O��;?-�G�u��L���ΐm(��82��3/ĩ���(c�܎�pRL�T���g���\���|R�e�6�G$M�%�3}��ӏ���1�wd�5E��w�.٣�Uç]�s�\�c*�~�������m^Jp�'��@$MBIE�p/6�C�D��A$���;��U��V�N�9A?k�zQk�ҢNEh���5 ����a"x�^4��vH��±�)�'�_iN:)۟XO
��Q"
���c턟���FY���Њ���V���t[Z��GC{��k�u�	+���{ڑ��n=[5�}=�g4�Ye�Nu=Ρ�V�hba�r��mIn/9�^m����"C�4�qRL]g��޷��&l���DF�����#MQR#;	����N�`���V.SaB^�0���~�ڸ���ګ��C�������",�$��mSGAo}���Κ��S�jgK�V�[*���5I�$7����6I�����B�z��g�3�Zrg�n.ͧ�T}��[�D~:`(�eYBX]�3��d�� ��O���~W��:%�e6����i��ƣ����9'
��Pua�;+X����JՀ`�RMW^U���/O��4 �n�b�8LѓX��{�_N�0��8pe��(�v�L�b&䅸���_Pºp6F$g)�eW~�	�#�(�0}SM�ϻ!S��=�M.E9�<)P�'m��(���^n�Mފ�������̲�J�@[׷K���Kl�}�N��n���#��'�d��v���T9��Ƀ qM����/O���ΓD�`���AQ9��N����/��9����
�^���Dq#�<�YSS� �(`�#/�
��g��Τt��>�,��S��ra� �z�_ቴ����"�w�
Ga�Q��;U.@eZ��[�{��P|jo*���1��F�V�M7�..����Zwl1I�䂄b�l�y��KcC�A��8ڮ�Ո�j�s1����N�Q���� ���!I�cf���?n��#)���}���,�X k@���hfܶ0�3Evg]o1<\��#[ͮ����T�ɴ��ϻCax�1�P�t���}O��E@ÿj���Vd��RIm���9�kC�0���5��~��,���U�9�~`�)��(��N��n�6Nk�l���F������	�D� m'��^��⯿=��O=l�=����x8�Hh4��ˀl�����T������!9M�;7`@�V�"�}_�	v[���Ps�u4�`�A����d��j��2dN-��7\�w�YղHo���v"l5�^��	g�\���޾�[Ka�{�>���V�̶(Y�G3A��f۱���:F Ⱥ�q��c����I!�d�L��2�<����r��K�]H�4���+Q�������H����� ��^�|�n��EG>��a�̶�����Ci~����z)�s�D�px���f���L[V�z�h��$�u,�}�Y�
��Ar��#�i�Rm�Jzf�u!%��N�"X�s��[akE/�y�Z?����59�M��
�O��PY�)')�X
`��ڡ1��f�3?�{�}�m���Hl�~�	*���*a�1�;XV����PG�HBI�'�k��H��Ǔ,�|�a5�3�K�Ѳ;K|T���Z��A�u�.���V�W���n*�Ɲ���$#g�!,��O͸S�4(�fF2����4~�fQ���x�����]��E�Ms�}���٪LDβW�!k�f��vS�W29b�1�c�*\��
%���1��m.�)�U�g�[s����#{R5R�Z����õ=�kVK[X�̺k��7A��݌�{rB��T�*	�[�`��C
���VR�k! �����j��弃MuFF�d&s���)T��~c��Ĵ���2��j�|H*E'T��5?��"��>��!iʹ�jߎ���W���|X��䲸X,L�Y�VJ��=x���@�)r��돤�o0�E�I|��@˧���Ε��-�Ն�-�gOE>!r�a�<>��O�vL,g�����*ǪǫV4��E��#*�&�Aqk�Q:uнUe�-��N����ȹ�"	�G��ƚ�L��3�J.
)4�����z'(����4 8��a'��oo��G�\+��Ҁ���P�*�sM�>W��Ϻ�*s�%7�5ԉ~5	���Csn�Sc�/�@=�8�W���8]��,{�C����Xs3� �*E;�J�\ e����,�4�kd5�c77���~����$� QY8aġ�d3\���3V��I�S�]�L�qn$���<h��Ta־���l��я�B�F��d{��Ū_@<]�O�g:wg�gj2$�Xr>m��Z���;X$�����mEmV��t�:�)���1�̨�H�0 m�_օ��Mݣr����+��:���+Zfpl\��*��/} l�
���@m�CАd�ih��@3�6Y�*�%���5��/�i�$�6R,`g��G�� 5mQ_9^~ ��z[g*���"N';@�����]���:�}m�<�u����P���q���݂4#U�bW��Ţ4|VX_Qy��@m���d@fx/�So�J���1�|3��6	��Y�]fl:l����VC@-6�tH%.#O���a���8�l�	r�2�b2�4�������0�@�Ii���]*TZ0�mo���z}���J�|���iI�� W�ҟ���#��W�J_w�=Z0,�M�PZ�	�6-��)IŊ��hD�?&"[c7J4!�9�{��3�ظ�+�i�ڔ����WF�q�v[M�=+O�OW������&��y<w�P��e��)�T>?�uD�sh����P2�Ez:kR��z!�+f8E��k���Ǉ������������X��; 1�#}.<��h�L��EQM��O��s�СSK߉5��e�����ѷg�����Ð,J��Ϗ���F��.���I��Ǜ��'�{���[ҿg����E���!N�>)���74��ip������N�,�b���-x���lB�N�Sc��>�3ҾS�B����)Om<q��9���9��U�bWi�^��4E�kQ8�����nu�˓3����.���(C�٪C�j2*m�2�:t�9��XS�sW^���z��U纁�&gF	��xp��R���a�Zcפ��J�o�!�
�S�b��s�RIX����4�.��1����C��"�mS� ���a՚�O����[j����s���9=;�v$��m�
�>rr�Md�P��) s�1a�����I0У,e6uĽ���7�Ey*�W��љ�Q�/�@���WL>C�i'�h0��P B�VW?����r�	y߭�CV��ū�9����(_�ی��j�����,FG%G������d����<�A� ��FI�Y/�0g�&��I0�[�iB�EY�RYL������H��{C�'���{�|�j�E}洖��_��9'��Xy'V���g��rfϝ�9ui���aq+1tz�Box��xK8Yf�j�`��xv�%Dd'�����=�6`=TٌǬ�[�c��CtlΕ}H=� �ľ�p�|y:���-*��F�+#^j9ov����N��|e���[��l^V�q+ԩ1�;��vv��[�N`�V���,Lb�L���=�}�T\k�z�'�YH}�vɞӱ~!���Y�ͺ��UE/d�_<��8�!��D�l[�X��A��Y {�_U8R�۵���/,�����k�PvH;�BӠ+�v9��L���4
j��#�C�Y�[I[B�8Z��ci�D@z*��>+��"���[�a���������z��Rxm���Y�J3�KO+��RCM� ��0%�H��F�ؙZ���N_P(O3��kqX-���dY�����+�VZ��� �An�i��u�/y����^~�����z$�0ڟ�����e ��q�Ȃ2�����>�f({P���!z(fdF蔇�m^�
��ŦY��+�(��w��x�������`��C�=�Ej��[2$��kD�T�^�V(p�u�c}6�D�T�>���;��(L�ŠJZ���Gp۵7�<�$�(����с�������������܃����-��G�Y�W[�\|;_�һ͸"y�6C���hj��bL�n<�HU�)6��"^+�66�1�	��C�H-���Qc>�;Y�n5UZ`-C5�5g~r}�N��-�6�J݃�)͓����v�^� �]Z�Z��G^R6"�	�ky.VJT�ʪ^����*�;���Y�$���Zo�����V�V��=��|�M7�U�I����k8<�{������lbZK�)P�'D�U.<]9e�j���Sw~(;[�\�����E[�8,��?�v�F��oL�숉�PP�,�>�P�	�Xb5:+Х^&)/}1�tf��e&��)j��V(ٯ�Н��e����-�Mz�Ԝ8����MA���>���q~�����,U8[���]���;)�K�n���|�G�5����C�%��j��`q��3+��{��㘚1�8�H�g��Ў��x�ub��8���#*�
ܐ��{���dR��-��
=�x�4�C{��x�y/���B,��mb�Tm��/a��}f��-I�VeB{�����H>��8�S�.��R�b�W���F���iJl���̖���ox>�NiF�h�R��e$�
G�l@�� ���lW&�S��C����ɋ�j�`=ߍ�n�t:)�v%�a��l��\��ѷ�(��Vk���V����_j�x0�d��y��Oۜ˱a�j�ş��6�����Lx�n��o|{m�E���(����ѐyF�e�S����r�0�7JY4Jǅ������1�����'˾��?���m���X^i��7�ftH�3B�"7��Ͷ�^S�� "���P�flq��X���ի#&�>Շ]Pd��J��nfX?�Dn�͞�����ka|As�G-[<���(�D��j $���2���� 3����/�V<���ݷ���a�%���� z	�-��`�gc��O�!DFK��N������?h9��y��G�2t��+�F��з�r��^���+���<���`[��+6���t�1w�ATDȣ�U�v
_�Sξf*���غc�M��k0�ց���C�|^[��˳��}�#�p�k˰�@`���M�;"��Y��8�*SF;�)�
_���\^��In��c-�(B��֪�����»`ܕ�̉8���u��oV��?� i6^!�qk�J��"֐�ہBsr2��׭��߿M���S�O��q�[�&C���?8�RLS��f�X��*�Z7�]�V6���_��W��@��^/�-�������߆�#ŏ��=#p�(�w=���$��qrś�[TJ��bγ1��`@wf���Q�_![Yc�k�f�-�z�^�ҫ��J)��G���R����)*��S�2ٳHbǆ]S ��+�$��z�l0��L%�!E��r�������kV� ���AY��z~���~�����s�'ua15JO,�̜�=b�������ڲS_���'e�j�����x��`R�i#�p2�}�����n�&[C Q\��ָ>Mp����4'��
��ܿ:C��%�-S��j�����z���릴v#�j�]��	T����%=��a�U�����w}S ��Y,UА�ߴi�1t��9�^Z�r<�Qs)_p����{ �J7o����쉙o{�E]v����a��W,� ���"p �=�����ۥ����M0�K�a&O��"n#�O(��u��qЋ���U]R�l2xa!s��@�ٮ�&��|ּB� �ׅF�ƭ5����P�����>J0C;�9�z�:u��Q�O
���a��7���a��a!��^��I���ຍ��%X�V��qL�v"?+&t#,������b�9ɺO(µe�Ǧ!��6��ȯBb���]���� ˮ��uD��S�� �$N��=J�zE4����IH4?m�Nz�o��h ���"lO�����;�x�FSY�9�����Ζʠ ?Y��_�.ogQ����o�O�Q���WL��W[�@�iIʄ���#yl���u-�W��r�	Dz��*(�+�ƶ*!}�{O�-�����	�e������,��b,�M����?�"vr@ڤ5�x�`���L�!�0K�Rdu���%�'��χ3�}h�7���[��$� *�(iU, sc �@�|�j+�����_��z���H4�����V�7�;D`��S���2~h9:�x㾹Z �8J�4�S�o���8i�k�N;A��yc|�b�0v�m.Ji&"��M�<{�':�s�ʹYo���� !u�O*��@+�&;�N:��Ɍw�iD�����V�H�����yvW��_^������q(Jng��l���z�X�-���W��<�(�~/5G��jr�̟ukϓ�����s���<�j��� S�k�F���C5LĴ��F���!�:�.�!��ٝ7������(�B5�$� �N:��9�~�8��u5��ZA��ӗ�d7*�1�6�������6h-˾�w~�Ѳ@��4��K_1��)�HG�����<ݪ��Y��E�(�C��pd�AqO�I*�?�{q��0@�����{��I�~��X���㋄�`������F)���b���L���'�^��1�x�i�]�r�׶�u�<�?��K�� �l/�XB�TY� �	q�̜�z�|q��_���6S���%K0���y�uF��z|�VQ��{�$D ��G\f3��4�HRR�b5���习�j��".�ϴ���+ ���X�O����������{�[iu���#?ʡ}TFmt��T���� ��������G�-T|��\Z&x@e]������0�2�X�kYs+�nؿ{<�YBxˇ�@�휬�X��L�=Ǆ���6��u��Z��/�lq�r(�F�z�Yj؛6��B������)}D.X��҃>k���@뜿����N�N���?uy�������#���Ҏ&��0�f�����"�Ó�O�X�I{�A[ �S潊c|����2��O�|g�ݠ7O��if�b�rL�@˶K�>�3f�>M:3HvyF��j�Lע~��A�����y���!_�v"]��Dq����F_B�\$���y��o�4|��	@&Nh��c�&����Q����k+��D	��c�I�s:�V�5����m��c��{���iB�p!-�[�T=���h�Q|��!�OjNE��3���Ex��N��	o��`� =,�ZUbg�ZT����؇rOP���y(U�@�~UqC���	�ؗ��X}}���2Wt7�X��!�kH�c�4�
�uk��(~ AX�zf%Bݛ�!)�,�������äQu
 6'��p��w���ؙ�້W�<Ӈ��)3ƿ�,�[�lR���!�,H��n�6�
gxi2�s��(�tx0t �$��%�����,y`5�-�)�,�=���϶h���j]H,|v�sɫ6���m�O���v] ME6�`Bl]��g�n)W�τ=��f�A�ӠK*i�:R�纘�B�������&�!���ӆ볁�ƣ���X!Z�gp͏iE��y�~�y��3F�0+�e�l�j H�8�E��L���0�v�r�*E�
~�~���O���P~�����e���"��3�m��a��� !<�;.��;X#%��S���O��J���қ-�A����h
��>x�]���!�=8]ԖP�Ƙ�}��
(5��3��n(��/���|���g=���oj9.+iAa��Jp���Ƣv
��� aBZ � `T��΅�A`�E���dD+�{���.�sm���*��G(^n�|}�4�Ը8rE@
��9�i�n�.�j����2ok�v ���HK�&�Zxh�S�p#��=h$�����yb���R6�=��q'5�4!�L�d��Ԗ��z3�>�݂C|E�i/sE�����w���:7`>":acI젴��QE4t��B2�Op���C�ݤ;��ɸUi>(֘����=��cPґQv��w���=�f�aab�V����9]}�#����㜄��Xc��LӀ&5������3 �l���#��uW�025�`���wX��V��*�%O�讉�=���	�[�>b�}9��d�k�d0�ӓ������	�7_���s�5��,�T��ڕ'�4�'��1�
x���:?�"=GM�Ĭ�jI�˔�Ụ+�uD.�]F��.Dq嘃��g�%�)ٓ'�ުM7x�@�yo䶐w��{1�Y-7�JA�������������-N�o��	��%Y] �&6���