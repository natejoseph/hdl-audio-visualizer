��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�v�-Q�Oͥ뀥d����8Ȭ
|���Ye)��	o��y�}��!C�_r��Q���8h��/����@j���/HV�Q���{Ǌ�6��m׊���!u}d[QN�VĔ�Ӵ{�����(Y��yH�G�Yx^=����C;�&o��Py#�}��%��^����UP�`/��Hj?����!��gĿ̋���Ή$��Y�����r
]i���l�f�E��M3������I1�d�)\��2W2 �^����s^,V��w?����s����W�`�*e/[�`˵rߟ�)U���.&���ےs���8+"�L��`�`����Q[��׆���#����v�Q�@�#?�:|>m �H2F�-n^�m�ń3h�k�8��T~9�k��޼,&�T�)��[#![�fiM�Y*�T�h�V}�k��#:�|�c����p�bT���;�}Uq�jw�Qцq���I1���oi]�E�<�akC��M�6%*���
즗����e�2P�W흇�H-̜���]�=Ԇy��Qw�{�+8�[>�)�5Q.b�� ���.#b9:^*���|��@�Y�$��XO�c�;f�C_nɨk7z*.�	�f�#���{	�N���z=q~C�\��i�}H˵���?Ҍ��r����c����̈́��ux���+�#�٠Zt�Cw����N6�N�5S|�л>ٽ�b��5���1�x0Y�A���d��C`/c芻�7ctt1<E6p��8�R�Pw�.�#��� �Y�������~��+��
~Sl.����j����d��i�~��5b�ČB�REwh~����?��g�3-�(zRGh!��$�|��e��B�ƫP���Z��26�,/W��U��E�����X��%hm��k��#s��(�C��H
��C���HbJ����%�����m���8��֏v�����2I����JkZ>� �ٹ�U�z>���Ь�`>�_��]aZ���7�S|�@�ܖ��G"�?h;��8�k�c[�6 ���i5�Z��_��� �T��N*�]��� )ۦ3�ϥ��hL�	������R~��T�Q�`���� �����)n�qք�e���h�����1�]�״�P$K#�emuY��5;<nh(���V��o��-Cb.k������T�0�ȣt�����Z���)fPo�ƹ������f��`���0�q&P����?~S�����39��<�LVM�K���a��-�iEG]��Ef	�2^�;������}�������/|����w�@�;zͿ�ܱT/�v�>A���rH�}�co��-�@pH^w��1҇%����@*�Cv��Dw8p&���3�t+ՠ��yߒmKh-]FxJ��׬U�B�Ӡ�[������>���׀���?Y���2���t#U�R�|���'S����-�O��c>S��Uk�_�~����|����r'��u(/Ņ^�M]�P��������\P�
�d��ҏs/ڵ�����Ʌ��Hxh�M��cl�]���Hs�:F�l�0q8�1Qàc���n�&΢	�Q�`���'L����CN�o±z)9�f��l�i��m���`̖�&k�j*n��%>���c�ȾUv L�h\�R�#?�`�}��7g`"�M��U/͉��+���s8�\��'�w�%G��[`�'�F�X��ػ�ȂB�g�ↇ�	�I M�)6"��$&Q-�h�S8o;6)xr�M �f��c����}]�>0�
�q��������	9]�e% w��a��3��>־�gr{��bF����)��r�n�N�A����<E.?�:�W�?�'��bi>�u"�1@�Q���W.�~��5��v���ǉd��_�e6���f�VC7��ɻ�O��f�usՒ0F�w��c a�2#ك�#(mچ�*�d�dQ�����[i�6��\�ĳ}��uz�A�r����P8.{c�(���b�.i�/ݫ%�`e���{TL���>�ƪ��ߏ�ޕedMMj�+?�і7��_��)ϼ���>�������P�%S�TE����/��"�+")�D�C�/�|#���,�f J�s<v�󍓻���
�bv	v��Q=;zV�2�v��Jl\?�0S*������Z�bdd���QDB1��b �
��j�t_��/6�5���K��@��i�4�eS�`�x?� 3�5�p�o�}�;�3���̹zH��g��#���uI�����vݥ�ાVG��h	=)sn	s=�_mw��D�6�U?�-�>�Ԝ:m֮me�Ҫ��Y�״�&$�l;_�q�s!?5���U�-;�K�w��=��CmL�$�C��+};�?�;��7+�yw�ֵQא'bv!r�
Ƞ�	��L|6Ύ�d(h��Օ�ɉ��BG���=�%S#���E@�V_�tؕyФتqkP��+�"�6��f`�Ѿɞ�督��O�&����7r䳙}��J
7-�&>ų���]ԟ�����ƈV �E�#��Ղ%̅��S(`���0�K��4mNT�CLp�I�_���Y��Xԉ��H�o�X��4sU,��?Ɓ�\�al��T�MB�p­rD��y�L���f�w��q��*d���{_��]t�Z(�՟�+�����黁��XT��υIQb�Tt�}n�;�@f��r�s[iE�Z6 فIi��Ɂy�݂4����}�DO�UB@s5���~����7�g���Z&��g�CQSVS\;��8WF6�Y5}�ɜ�N�F�c��>�Xr����B��?�1U���|s�~A�%~�x���MQ�������F�� ��=c���Ƒ� ���@��P�0�޿'>,�X��ԅ�&h"�߃���c�n�V)�Q7��(�k�AZ���Y0L����?V(?�)��1�n�s�Q��#�C�I�\|�}��z��z�j�fP���$LlIt�<�h����)���h��Q���u�{O��0`~9l�@eE��һ,/�PY���������#�����3��D[Y�����D �������_r�E=-��4��{��5�脱a;� �%��?�
�a�G!��<"��S�z^�}ܿNge4'-�ҵ������"F'�R����S��r�z�5��*O�;�\�:4��4R�؇�!���Ҽ4bqY�߫�a�uȵ\�&�����|���@�%�pdK�����h��d��ε�z_r��?}\'�n��1��y��=��|<;�o�i��V3)!�-�M#��{T�1�-���.�t`IWs%�p.f<��=���1�>�E���ܬ��p���4�^6(�)�
����i�������d�:��i�6��ϴ��{� zH����]/Xz\79��:���f�+���,��G0Y�["��38/���^��¥�S$��{��T�<��Ցhn����VmW7R�� ��ŽM�xᔁ,�n(A��*R�,U u���2�`]�&R_���"_Si�WR�T-��5����#9����q�����.���P/C��CG����;a_\���"����Z��O<�����,i�?�@�.>�g%�#�_�jǺ"������f?�R�\I3�
B%)��e��_4���Cg$�x��g���hМJ��*��_1͝���&��n�R�>Ñ��|��/.���	�me���Og���S��쑖g:�`���@J���c�3-m��[\�ޗF���5�q��e�?��@����nub8��Tm2�t���xv������xfdW*x��(�����!��5s�5��L�׏�o�j�@���Z~�Q�����ۿ �1��syZ�̊�ґ�u,"�[0����r���/�y-�G�o��#Y�|��FyR��~��)�`�Wes��e�� ��̍o	�3o_t%�[`��*��l�ZM��l�l���'X~u,.=A�C�r?����0n���A��4���t��lT�"�A�3d=�*�� _�� �l��%Ŏ p�Ws��oa�uMièӞ��m���i|����˫-��C��
s%�/3Z3ՏX3k�_L��N��"�ۂÐ2^o�w�lx�\�����5z�r�ڦɓ�nKbPՍՂ1��C+C$��x�e�'�X��]W��~h�a;�i��/Ǘ�?�Y�I]�<V.ZGw���@�o{��f8��脒H]9��eB�ш�=��I�Nq�S���$�(�N�l�q�P��*�⏀�f�(�����i�L������5��;�,c�,��{0s��6�4
��y�=����]eD3��<��� �0�B�Wy��0�b�3)pP�G
�{��\h�!�7��I�w�G�V6����3�\���A!�`�񦪼��Q�3F5�4���z��T"�U������UY
���,}V\b��$Y��d���|���)����ʧr���}���&�%D�_;��5���CH��
�zI��K��JL�kl�BpgP#�����}V�n<6�H��Pِ����0�Y?>�啗�wLqvT}�����o� H�L��.��j��d�"zA��~Q���Æ���	�=�T8��9�n�	Kl�l��B&�p�U��P��fWΛ�<	�m��5�D�W��K����;��c�qKx��^9iH qX M�>󯣊KN\iK�����6dN��{s���H^�,�6��H̒Y^;I����lΦb�ڴ�me�hܺ�ʲ5�h�5����ۺ�$���,��J���A�v��[]�	��$62o;)��J�醠d؅{o���Y:���-���K�����]>�M!��K��]W�d��8+)e)yn~��QT�<�8���W������b��7I\�.���|g��gQ;p���o9���Lyz4����*�K��_��@	$J��pmN9J,��GA�1�C:�Y-���*�7��9��~ݰl��4WB��}�v#��͐�j�DP�=8��e�ucxx������Z](Dh=.0�hp��l���q}�=e�a��=���Z\�¿��dۑ�U� ����j3���a��<��Z*p���Yƪ�;���$\h+����R��$=_ ����Hc$�ԭ��%����w�c?�5=�� 5��Ā��Y���*�==y�Xd�@:VT(w����5fR�K��պؼ�����,�캗HG
�l�����JEԞ]\`�0T�'��]l����R�VOw��"� [i��j���a���EF�ȹ��-˭�(������'�����G/�tkɞ����/:��u���	:�"������_��(�fdN�.&��Re) jb���In�c �Q�����A[Y�s{��N���� �-I����/�m0�M���~�Đom�FUs�Yz��4��U�Xm`��JК�x�:�)��:d���eP���s~S�/�eĠ�~�G$�#�;T�^�!����a�/����<f^����=p�	�ۿOW��U_��$��(������A��I!o�Y`Yx[La�n9ZVLY��~k��l�m4h��ׂl�;,�4��ʮ+{=T�3y�a��,>���<+�������N�C1�w�Ȓ����V��!ޖz'���u���
����>��f��K����ğ��= �f�=&���<Wn+n��j��U���ꩽ.�x�A�G�7�%& ��C�hY���k�-�J�.�>���l��q��w�?+~���D�S(PaC7��V9֖u2�y��z���F�!���J2��ֹd<8Y�� �c'm���L7������Z,(����w��%���H��}���Z3����#�\��Q�`��uo)7 �AǑ;��gE`�)!�X-�F�իGW���z�Q�+�3�	�1�ʉ�b����b0��
�ݥTf;�.�G�9*k)4I3��^|�0��bLh�C|�D[6d΃�p��b�qۅY��h1�z�?ߕe�����)�W�iςW֝C�`k1���r��c�d��r��(�REp[��:����"ϊ`Ȣ�+ �q�<����Iy��;��F5�zi/��)C<�%�xci�hAN�rcMtm��;���52�6�DP��\q5qL����۰'{4ݫ���8ȳ�|1��$��Y�(}O�ֽ�C���㨹���R0��*��d��^��>k���y�*��a:ss��@�_*:!˕>�L�S��:UK��h�2�3`8�T��%����e��Q\�k(g�D��l���Hg���#�w�ST8�^���YtꉰjC���_�4�H�$1���e��*ջ@����(��"���t'����!�Q YVU����u>��[��(t�?�I�3�[˫1�h:O�)�
jے*#��ME4����.E�����l�.��=?������u@~ח���u�λl>+�>4�~u���m�����B��c��>�8��:�+�W�`�d��%jA�e{L��F��R�����떺�28ő_(�>�4,|�8֡c )̌�z�T�f/ymG�Ɵ�������C� ��Yf:��i����!D(ʌ�@�uKv&M磭�l���UZ�ч
p�?p'~�*D���hH�#Qw��Wʺu<�8��`0�|qF�x1^N�8������9~���G{՛��$�Qq؋��;�췧�||t�:̵����1e���P�J��.�I	4-7�>zgXBs4< nVBX�t�I1l�����&���"�Me�J�Ҋ�f�� �\%vC�4��Ɨ&	������e�o4}O��^�(�H���?Ђ~���g�;g�-�2�7S������QV��tmi�4�<l��T��"'OP9(K�X�	wS?CAG�Җ���h��f�~{$Ǒ��JO�c�y\L���B��m�r, ����amY����7�H�Ԅ�xL ���f�-?B_D%t��z�~}q�ݸ䅗�,`��jB���Iy��ntneo��W�.g��4}�IY����ԋq)%A���x�|J��P�g"_�����e�@`�5�o9�D��ە&���0�SO� ��shx���Y� l���Y���w�ٍ<���-19'\VD%a�*�פ��-ަH�*�)����XQ1����%{�d����h.f������U%F�ܓ�~�f6�� 1@/ ���x��w@��͋{O �Y�Vw�P�����gv���՞��L�v�@���[z�~�-Y��d7��E�^�c��<̀u�iI�,���v�$�9�f�1D@��Ǟ3�7�GWMߔ�;��6<���sMx�{[1�:���W:`���8�Z&'n=��L:��B#�X��1�\�.t�������iA~��>a/j2�=C)�
B����r��o�^��D��9����?Ɖ͉��g�
�$G���N<�v��J-G~�t�8���'T�c�c�1m����O��>w��cn�1�l��o7UI���U;k��\E`�r���?�~����
�C!� ��l�!������E�4����2&�y�R)�@5�3OX��e�S+��)z_�b��ٻd�g��Nd.���]�t?ȉ4�/+m��ƣ��Wȫ�_��S�5�B�_�f�z�K8��N�XU������@�&*!l�E(�:�%�B�������s밧��\4�	�/�lu!�a�_Mh5SvP�KGZOm�q�{���TW\l���\T��z�!�2�b"E;%(G�W��vMg���m6�iߣ8��m�fG�0jߑ�c�H�0ŨH�:��}N���g��V��t�>��K邸��f߻ם�H<ohDk����Q6<��	J63�ѳn9|�Db֝ES���Ek�juz��(�oS�a�r����(V� P�1�-�֩ø����,ׂ}��m.m��j
�R�q��O�f,|1	�A�sƼ�����˧�)���UQ3ٚk�3p腛F#.�:}2R��C<�K��_���%����^�~g������ESь���Q�OьWkq��w��hxȲ|:�u"�rCv��}�o�KmS��u���]��K>N�w��>�z�@� ԭn�/�mݔ���ZX�24�532�\��z�����z���.%��W�K&�ˮ���o���!>�À�y,�np��L+��T�`��n=7!�U]�$?'��bh�}��m��?�v{�Ǳ��/�Eˢ�\M�{oh��Vl0hGV0��+��Ϭ
�b�L:_NJ!��
�����.�OK����q:QQ�,U��
X�kp�D��jZ��L?R�l�B�	�`��!��X��l����1ߠ �0G�4�̔�V�>'؁�.3!�)8�Q�U~��I��.����a�fa��`b$C�B��죺>
�0���A�����J�q��ʹla�7����f_��>�n���;̥�+E�a5
��_(85M�J;P���5|j�V��xӈ�(�?��[��E��,�lك��]_����O -y���}u�j�8��1.Ɉh\���1��o�%bp8׭���2�5ɿi;���)�)�Y8kW*�WTH95��x�+����zO��u�f��iŝ,F6�~c���^B�$��l_�zi�z��/I��J��a`�b�E���9hVv���������V�ԞEc�����S|�R���- ���kL+�M��U��ە�M*�e�?�r�H����K2T��l���П��u�k�j�,�nxm��ޅ.�����'��﫴���L#�.��r)kxR��$8+���~�A�EY�2�Z�[���l�O{'��/(����9CQGPbT������:W�{������o�f�X�� �]���ӣ�>#VX�cp�X�4n�l�/���֞�ͽ�gV~�4�~�Ɉ�f'%}++�_/��/?u��YAk�z�c �R����ܱZ��7?Q�ڻ���1̫�"�)�k/e0<��i��c�0�oUQ*���!j'"�]e9#�j����Q�f���ʓں3)�ß|�d/������f�t��̆�Y�:<��s����wg��i�G�����9�Q����Li���	^O	����&h0�9|8�w�Q�a�r1�z5�� ����n^��(G��]��?��%4�XX�`��`���������+*̰�1��r���{�N�3�H����eY�w��|�+z~�3��2��2?��=+I�^�K���؛,Ysp�4:��^g!��Ȍ�Y.���t=�U���⪋^��Y��UM���a�a��ݽ�K#�+�����v�+ǆq36B�[����lfp��0���,��m�0WD�� v50��{QL��0Z
h����gAW��hly��E!��-����}m�1�1Ѹ��'����iϫ�Z�X�OTK��}V�q���}�� s�zV��:ʼv�nk���?�y�{�nth��N�zqU��s�Uh���h2�x~�l$�"Z��I�vJ�~��Ƈ �����Q�n�r+��"�v/"o0��uw0<����B�π�}�}�� �Vu��r�����x�܏HK�h����,�=U�#��Ӏ"1P��7L0EO7c�!D�8g|���>^޲��0�x�r�ߣ�����H�ӀN�|͹b�+�oB��2�̜X���dv(�p��M�7�B@�b�����V.�u����
.���B�mC?��1�Om(1������y� �����A���[�Oy�Q�J�uc�^��*�Di���Tk���ҧ��#��K���M(^@S���!��@�A��v%9� �?%��j_ V�$�x�k��U8Fvx���a&����U�m p�A%q�чa�b�~"y�X������}��d��F�Lf��h��;`
.��%���'�_�f۞�tw	�l����z���d����N��#�X~R	�V��I"���G�Eb��=���O!h `�Ń{6&dm�`���S�7������vA1�PQ��`������$�
�4T!���q⌽^z�"K.O�k_ج4W�]�O(��-��V�g�u%A��x�"�?$�n۟D����#DxB�T��v,BH4y~��.n����
��Vwh�]]G�PM�E���I�1���F�F�e':1�s\����ko��ꜝ��W�H\Ej�2��q,?��`P�o�P��O]