��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��ݷ����M7P����˱1W�����@e<���vL2C\�]'Xwz��6)�	;�j���:ݥ?ܲb0�*��qd��=�m8�edSpE�;�;!��I��R�e6��ܯ����oP��m��Sj�I��µ�_h�5+�`�9��y�w#�J-���S �-�B�2�7��#�{��}�.��b���WJ����I��E.�x�j�ei6l_���9^b_�TNF[�kw��D���)z�̉�k���Nz�Vc*Q�i'��e>2�v�KJ�wx��Ӕ7�I}��� ZePw�D�R�߃3���Q6K�e��rq� ��fl֜��rw8�$щ�R�E����z�S���Ѳ�\�f�J�y#	�P�Ps�V4�X]7�w�d�n�U��ڒ�Eb�a;������#h����8v��F��+D�(���ǲ�(��0�"1��iR%�ͥ9��B���^ZH[Y:�7W�H�+�=�n����Pr��=����(3)U+Ah�[��,`�0У��$�4�!C��;�?d��=��d�Lk8r�R��:�P��O̹1<�����<cYF2o�ߒ��!��3cφ�T�
���
B_����e�.w�'0��I�(J��wؼ�H���`h�aA`Y�� xG&G�Nb+�ָ�^���Ov�����L��T;Y��}9�$[0��
�n�U͌h/��=7�����fŤ�1PG�I��C�%cX���<=c|#n���	����OT�xe�H\�TX�
��Q��[�y�eI���.�*�!���퍨o�.p^� ��^M�/:y���W�������D7�cP{%:Eb�i��ʕiZ @��p���!n$���U�)4e�4���.2w�J�v��O��i]��f6��3!^c#���v�
�$�U�m5��X���NO������>E�v W�,����$�Jl�pZ�����P��7J���İ���ۀ���Z�MnFǒF���$Go�-�����L�9Ώ���v
��qkr~y�eunS�2���f�9{S=�M|��8�0K>)oNC��yuK���^`�L��@J�ޔ���X
���.�K<�Nv���/l ��<Ӕ�;+�:��sZx�[�h�vq�#z �3���b#:i��<�Ӓ��5�C�xs�uը�	؊$K@U�UDMOߓ�����}V�S8��F��2 ��D?�y"�K�.)L*2��XL��r����H�cъ��y֫_�]yz�� �jgs̼� ��aD�'���T�|=�.���S���u!�RVd��&%{u]Q[��	��u���K; ���ȓ[`g=�_R'�E!�������^X�B���x��2�&Mǐ_�����IF��M���X�2�^칎l��+&C��~mJ��ƪ�����������el4#�f�&����q��,���,j�}�l�cQ4o�ٔ���T禮O�8 ��ø��[U�^]ҨY����I����XR�:zl'�~-�,�x�=G̐��AO��aΣ��h�/K~d�4�@�+"-��V�3�ܙ���x����O��(EZ�=/��	��u�9�@t�κ�j�#Q�{��M7?��E"�>���0�Y����t�";��
���;��C-����OfAw��6@����&\��ɗ���[��~��!D�t��"�+|��Z[<����eK�X�
;eUFT@]�!�D ��װ��w���4��%�y+�n(Fa�N��Ր�_�d�Y��u=3��=%����I�Mb'_��x�k���ĥu�/C�B���kv:���K���t՛ ʈ����Ov��vz�!�_X��d� A���ؔaBg�ѩc[N\�m��, ĥ�)�|��\%��J�>�{��n���h����h���r����c�#v%���)�2֖~�#���t���OS)0�ߊ�\a�o P��P��R$��0�Ö�ԃ�8R����ϑ������A�;v���0" ��>^*�mi&Ym��WX����['(pJ�lBC]��S'�6���m'����w�w2� sM �+ܛ�,�MG��O���, 
�q{�g��}ުa���D9�����'�h���Ohc��ň5�����"2u����ι�P�Jv�-�EB;�%x=9`�����o�%�|����5J�О���B�_�obR�$�N�&������4�[��D��*��W#
�_`M���]o��[}�r3:g��ݥ��a�1g���v�5��Xѐ�
Q���ޚ�'ϥ�Nb�X��s����AI�|Veo�Ӵ�C��!B!k�̷��
���;���I���I��u�V�����&H1
��x�RN�dF����(��lg��΄��?v�+�#lk4�j�� V'%�D�������k���}l�S	+��;-Y�
��f�-"�]� �� ��L n:��ŕ�}	�e7���Y�]�jno���C'�;[�*F�$K,�����j��ޗ��;�����"���K$�Y[�LD'5�DF��_*��]SL�-�m�I�[�P��҇j� z-+"a��1=������d%=Ĥ?{f���xq7�U�v�O2�\��ޫǳ��Vؾ�;��L���P�Q��F%gR+L��:�^���/X34�O��𵗷�Pǅ"�e�a=��H��嚿���_T����by�7��P�#\���
i&)�k�n�2Ajh�X�mc=���%5�A%;�1�$GKLH��6����e��1Z�h�4���s��D��Ò���S�����禪Ư'lN1��N���R�k�_�D[�ne���;�E��'w��2���uJX����PCҼ.Mk�0?��>��'���3��"�=����L��(�W�0�l}�v LS�.S
�@(�w��a�9�a�i��X��Hl��b�+
Ip�]�G����܆�y�K�ǁ,��toP������>��~�h��u�6�>oe�P�R(3C�X�c%��T4��/{���^�z��`>��F������+�U�-
T�ǏV��ɮ�up��\g��];+X���&i�x�h��涗R3(,7���G>�!��x�PB��W"O�D}T�:?�V���qT��0��ݮ���%�}!��r���QChV]M��w�sH"/cϻ�3�OGb����?h���N-7Joݝ6�͋vvL����ΡBW��z�m�:!
�'��9kǋR��-�[���� i�.�12�����: ᶄ�
p����rY��Z�x�	�i@�?�W>ΧV��8It"��Ha7K:�6��$@8�Y���AyD��b`1�^��ɪ�n��5�F��2�N[6[�}����b���Wi��"\���7��G)DMı����$TE�I���̮z���4��/\�3�O	�W�����ͼx�`�vp��ns�����xUL?H5�h�*��dD�����,[��ݾ�v�;Ϟ��,+Ǎ`�-�	`ť}�Mi�Ӛ�]��Qj}-��چ0v	����|�)�n��b%�d�4�D����y9+��1�zv,E�5�un�@O�,_;B��EL��d�Op�u�+�nq3bq�������<���k9,Y��y�r���#Q#n+y��� S����n<j\�|(7L*fmbSO4�t̡�>o���J����t�ִZϷ���F�O������Y�w; $�|�ʖ��>�VQ?�1�ն[)6���$�@SҜ�?���2DōO9��"�GN'8�"�x,l��q�k�7|��F�I;B�%'���X�,�L`G_��R-�h���2��4C�,�E?���I���D0�~�V�Xa��1�B�m}��Ns�L�3�!����E�1Oeƭ�������rc� \Ww��>&�'*����p9�f�		k �f�� K�I�񋬞A����F�$�jD�%o��
a�_gO"�yӆ�7-I�U|�R���ݠk	�I��+(Ĳ �n�Q���-���֫��Py�?�iF�x5��\�,���0+�sny��BA��+�&�@8��8���*!G{�A����J�ǃ�C�^��9�EC1O�o���O^�z�"�1�]Bˁ�8�Xs���<�X:��QF55"�􅲨zY�l�k3�}�����������N���8!(��aI'/'���{���՞
�@O�	r��F�ϟ�l�<�}qW�s;5��*nz�W�{�y�/�ϸ��/�UO��љ�)��n���늻��\>7y6S��VrBζupG�B�XF��d��ן�����	�ܚTh���������}3x苜�ԕe|blK��T�.,a��?c6�܅�<���i�Kx��ڍ�j�g��pf�����?
�jM�\��\�Ntĉ磂���w��\Ş��7T�^Ǫ�`��������?ȳ�à�Ԋ�{4��%�	�5l��)��C^�<��/<�jO5і�%d헤�Ü�i��J��':(4%��<ܳ>7�A�iU4 cRz�S��N�t��_�)�E�: �Ԍ*�e�\�_���:?�[����29ή���#�2��Um�=Y�:�?��8^I� ��-$A��:�%�W�C�-��ܡ)=ۙ�	1�m7������԰� $��hk�+	�ޑIr��D��2��B`��T�z����w�w�	6��U�,6�F�h�K�e������������D���:����m�W"��]5�T���o��>N���V� ,O�q�:��nG1�P�������n5����9�n����]'H��m������|���R�'/� ���}5�n9����0<M�'#�'���Ja�I���R��L^#�#&	m �{����,Ҹ��<�H/++_p@H=RS�RcN%�z~q�5>����Ҋ@&L8�@�#�\�7ɰ�\D�1�vV�&��لAw�j���`�<�C���	��Gj�..�%�{F]JK� ��h\̍��:B�Mpw��ʬR�6����H���M;���u��wُ��OW}�LwC�K�t�I9z�B������n=��1��%}J���Dl�����c�Q��}�������iQ�X��{# ��[��
���q1}���MB��ܓ۸�ql@"�d�`�]���_U���������[T����y0j ?�*AN��c���*�;Z��?#���!���D7m:��Z��6]T�>b�a~H�D�XX���Z �W������̽~p5C1U���(5��$���-��[�8t�8���%�Ӥܭ��������b� �6��
%�~
�
@��A@z	y/b�cL��w�T��I��Rf�P����C9��Z�pDj��p��"��o�j���͆�>\��T��Ӥf	��>���b�z6��0OxJo,ZUze@t���x�\�T����j�s[�7r�{��'�K�v�G���g��/ݏZ�q��%��M��|����Ш����p�M�Y1��ܚ�к���0.�I��?��������'D~��J����{�E��l6�$ſ����&}���63����(�c&U����37�U�DT���4�$IM8��^�ꡖY��+���~钲&�N��<�*f�uW�Y-k�1������s&�sf@�+<�+;����Zs�d�:�#���f��Mh��[��3J�
U#�Up[|���I^4�Q	r��;Ӡ�k��=(Z��d�G��./��ܘ�pA��x3D��[p������yY,�+��v�7<KnR��3L[�]��{Kw�=��$�h��I۞}��e<~I^���9�J|��N�܄��;�tV6r�v~5`a(�.�X`�1rF=ݛ������oZ"���lY�d$��N���[Hpf��RW���%�������D�=�2l�d�i��H����eXIQ�D	�!ήK�,l�h����Mc�6x�̞����q��.<�)���ԫ�A�#�!�՘Y*?���XnF�0g�N�y�d�u�uBƿ߄n}��	�L�%.x�D���ڀ,��<����Ѫ�K�dYZ%�R���*.`�-�9�8$��	�55��I���\�� ��O����O[���@|�j7@��t��&�99�שjf��(�L"��l����2���
Ш؈�:����S�mY!�Fo��+ j���!����nI�M�	d�����`��s5��Yp^��ӥ@��[�1e��J�6�bKR���a�A�D�6n�X� �����%�u��ڡ�At�����(�}V\�߁B�捋�'�j.9����U��[��u�뀪λ�,�۴F�26(S˷�H����lͬ��κ���D���6���N���/����U3��x�aK�cm����C\I+����=�G����� [�v�^�2����ř�q�	��r5���*�����f���9� �۝4�_�{�uL%ߵr�l�`%~ ��AY��_֥Ǧ�k���k/�T�/���'`+{�'W	�ioBV>�{m���td�&g�/}p �J�2�Eou����=ց�&��WYU�r @���;X�a�H���Kl�c_�DUEq�҇�(����昽K:濳�=�PًL��ړ0��v��å��\����I��i���p�X�y����*�:��?�3a4��GAQ/V{ij�f�%o,�(����h�7�>#m� %�.����hu�n.�<�<s@,4�����R�y���ѳ @�@E�Ĥ-F�r�����{m�3�5���:�;G#� <q΁i��q��ud�!4�x�>���`<�`n�V������#��ˊ0] ���]�H�䰇&��\=?�zA	,A`���40��1Q�{f���Qx^p��"��)���gy0䋌��&�f4b;V��N��4~@��3��]L�V��+T�a�)v�~`)9i/xe��U���y%ԏ7�s�CS�ѻr��q���.�n�
j���Ms\=1|H��L/w���9LhL��Q�(V�l��?�z�ճ��L%�t,$U����M�y8�<l�I�r@ �@�-�Џ!y\vY��=)�E���/#u�Y��0�j��/@���H��2tF� 7�I�����v4&�'�W���N�4���n$��8�#�����e�t*���Q<�Ҙ��:�n�B�<�)����2�����b�����Ҝ�</k�#�.8����e*���:�v8�;�܀���]�Iٽ���٦]e�n���]HУsE���]���F(չ@Y�"���Ч�>tK*��Vz��L�ސ?_w ~���D���l�p�01�W!���隡��+��6,'@�HL�`�E�6&�������LH(�~}0lo����r�����̇��$YY5B�/�����JI̾���E�;��J:|�8�ɾ�:�ke���{*�rp=m��&��2y�D�������rb�БG�����b�7��;?MB'�T��R �{�{	�t��%�����PG��� mi:��R�Z|�>W�f^FR,<��8^�W�Tx�>;�9#5!�ݹ��`7�ݡM�*ͤU�K���5�HV<q`���R+�PC|(�}��f^�����k�Ï�kӂ͏�9&����%Z�K�����xuk����>Ed��f�1�4�@���%6�l6��o/s�TϽ��r���Cm����aWOu�w�z���^������=��R&XYm��ꡄ.������NɢCY�ϣ�'��s.�2b����F���d��nqt�%f6��$���荮 �t�U�?21��D�S�\�T�=y��b8�
�����Sd�hکV�M��Da�<�S�PG��]��cW�o��A���U��O�L4�����_�k�M���fi�5��H�ȅ�(��������lغEK�������r�t0�	�t�Rˉ�h�ge�ǭ�MJ��������/D�ű8C.eԋvc�h���<�-ϟ`2%p|�/<q�+n�`*O�i��g����Q{��K�R�#(�^�lO�\͜�u�0��݉�z�܆�1��q��#�ނD8�3��)�0�����z���܃g7^�N��>8jW���e������,�%����h��HN��I��I	[�T�%���Dd=����� �cۡ��9��D���礘��D�3�zx���Ev��"��P�� @�,}�(m�=�Q���a�j��6[P��Q`�O�����b�r��|����t-Z!D����]���uy�3�f��3��C����#���DiH���/t�:[�V��`4;1'[�b,���V��Ee����Q,~��<^y��LA'r��=�
��C:��k��na�o4ܸ>S��90F���\������8u&�|%����zcXN�yd�+�е�9S�HK�\Rt�PP׋Qɐ)Up򕸦��dv�rE�ɏ�P�J���(�D�֖]p�Q�P��g� {B���5���3�C�q��8��rY�&$�r$���(���d+�_$
Α^^����O���P۲��w���\�� ����4��͜8խ��d���C�̶|���:w��^��df썝&�˛�k\��,6|N��_��Hv׀	�dAU�}i��.,���*C$|��Z�kC�I�L2E'8rq?x�vA�v�"Q�#�Yp��b�K�ۅ�y{m�˛wS(�gpa�l���m,���aq׾�w���[	.��#��� ��z<kN욯����!��w���NA�d����p���ۡ����U;�d)����3�l�J��=hbl��T���U���ї��ھD���ӷ�>�T]Q��aj��^�Q	W�ƒ�n�@�A����+e|:����#�f�VN8�ne5,?�q���c��⯺�}jD����!]g8R�����\�%�$ק�Q�~�2�u[J�����Zѝ��R� o���/&�z��X�of}"o��S˖
J��x�L�� ��J��aF�������@�n\fb�ɗ����U�:2���O���c`�ֵ���U�aʇ�y�J��1���8`h���o�w��T/��y� �C���tF!h� ��'M��}�U6�%��1U�H-�#
�(檹�[H�D)�	bsc�U"�7�fO��ھ��iHΑڨ��H&��z�J��e��z*�Z��ɮx@Sڬ��D+0���%�K6>�ˬv@u&��<8{y��w~�[-<� �	|�nH��l�&T�Ҡ���}��x�i�޼'��a�0sf�w��\$mr/�W��J��/�ϙ���)[a��S�p�<zd�������z.(�r�3=�&�lDOC�P��om������7�r�p��b ��lơ���	�U	IidI� ��ƪ���-�|�?����a[��&9�x�<�5M�F	B����I��M��{M��g�a@9�3�e\`�d+(�oUp?倶i����=#�Y�~+rmsZ�xm��_�$��{=O( yH�H��3E��!�<��Ĳ4X)� \e)Й#���kH{v�;Y���Z�5:ү���|����s�a)O"���j�t�\�Ŵ��vVr���hޒ>��l��K���q]�^3�����$l�R�%�hY�G3�:���=����
�!<�y��˒Tn:	0�� ������ �۞���Br�po4�����:�	���?S�&��������j$��!�˒��j���v̔2��˴��lV�`��+A�m���yHw��N������!�R�Za��.ztG�xg�\����gȩ�r���$+��fI˯P�k.��D��K2 �A$�v�7�4T���ذ��mz�fn 5�O������Ɖ��_3�Jɖ�q�B *+m�7J�4�԰?�o[��k&Q>����}.%s��L��Al`�N�8;�Jמ*�}����`y��jy�J�7a���>3��P�r_���|��XnkF��o����WY;�* �rמՓНj�iG��%�S:�@�V<qЊ�I�����evlgxˣ,�R�"��q�Zk	��_���?�/K��Z��U��!R4@Bx_�u����cn��/�%\�,ؕ1P�J��w��e�����}��6�/��e����0<�'�/#���pM3��Q�� � �m�݊N5d�В1���M�.%J6A1��o�7)=	X����:ݤ���j���	Q=
-!��%��Ǳ�+^�D�� ��b�tq��0�g5/#�����J|(!pa����T!�Qw�� *����_8;���3`%^�����LhYl{!��uE�@i�~2�c�q�Pd��j�w���¡RB�V�A�˼���G /�MW��/���03f@]�~}���@P'
�O�R�bFJ��b���3����f����}��9��7q#>C�x��1E��X�x�ef
��ΈQi��K�qe�դ�?=��̽#��ź��'v]giT�.���t�|�zZ^1KE_�"��P06�"�^��M I�3�����+zZ+���*��1nx��K�U���=��@S+��;��9��0��{ɣo/�r|�4��Q�KX/^Nfw��8�Ѫ������{e��\��!�����ˣ�����$��oC{���=3S a�*O��k�dB^qi��-�}r���+��u1Hrױ.�*�pZ��{.���Ly��r�����ȶ�4�j�TV�1����P�2�M�	g^�0�Z�������_���0� �5���O��C*��t�i�׵oTUR�#T�:�a4�����woh[�,K�Rys+�@+�N���PM�O-�)��EU�H�}�Xc&u$J.�� ��C�9se|�=�n���J�7a� Y�u*7�w_T<�7�۽��_����z)Ӥ�"���@=|e^q�s\
j�؄�ĺ�������?��˸�s�^e�,&rS��8�٠'�hr�f\��J��rl��>��_˙�
�~z����F��4P�.�l��f����U�z{3��oA�t�5Wl����Y�[8�4��!X=�_�}�ہ���}����W����5�l؁�#{����[5��x'"���Z�ܒڡ�r�
�-J��ؕZ�k9����-�P�8����Z�a� ���0rƹ�Tq5"2�/ո�N�W�:�O�_ɜt4�����l��xԪ����F�@�����-���Mr�*
�F����1Bm8��7|�ǂ{�ۦ�u�PU���L�E|��$��J,�'��H�S&l�)�!��b��l@�D�9~��� Z%I�"����Bǰ�[��{N�����;
d%��Bb �$���fp=F�OW1t8U�JƊ���4	'%GE�և���/��7���40N6����!��Îa
-����pJ�����QIs�:C��w�7r܌�%�]�o(rk�!h��0zUw��]�⫢�)�tQ9��.�����џk�
�����ĤB�xX�b�~E� Cʓ�o���ny��hՙ&pa�V���3�LL�9^j�дLI��A2��=[ӳ��B�9H��)8�4J�׹�ώ��͒f�Pv�z<��)�� j�z�sr���Rƽ8�a�C��-a
��O�Ģ�<�G��VݼM��N9��	�1>n�{l�֙,����v.�*�tj��̶��#Ia�W��n;0�_fS�_�L(�XGn_f�k���|�~[iӴ���p؋O ��>EZW%[	b;�S[�!O�'M6��L�"ٹE�	5c	b10~W�ͽ9%@I��Ց��>�,��p�s����#�i��*��l�|����K�r6I�
���an&�518��;��+��V�1�Y���H�� �/�/4}�z��J���m[*v��:cY!�-�)4�\�#��
O�J�)7���EaN+V�k"�i�.�_0;_�8w����o0 ,���[��	o�HŹ�H���;2�2
��P��,���Xt��vX3��«:t�D��G���+>���]�ًL$��h�����ٔ�z�$�$̻�%[���Cϯ>��\u���&a+�%��^2����1�`
��x"�ٝ��<�w)�0���^����4�4k��ȃ�ogӢװ����y�����d�Ҥ�_�IH(�h,�����U�lc�+���h�u7����3_#���;$BJQ-����,e�y�䊑�Ó}��%���=����4�<�\�b=9v����\��+���`%�gS �@�F�'�I�7�q{1�.�����������0'�����I�������_�G}%�a`!��ϊ�zz]��g���w���G�P$�$(vLH�ʨ�O-����t�����7am�2���'��ó�ϛ�Y������Jy���oP�.��d��eO��U n/�[���!��s!��^�n)	��M������	�P�E(���l�H'� �%b����hv�bs)]T�sl�Z�]&��b�q(�w.�7.u�`d{(բ9�-�m�&ܯ=i��Y��d�)3)|�� z�`>��H�j��'�W("sL����yo g <6YdջU��=���ߖ�r�uT�%�UF�>�{𽨏����k�i���F�Τ߻]�ӱ�����:V�<fqq��(�w����̊�߿p�g��(�ּgg��-�L U��H�G��qI!0��0��b0�F�9��s��� �C*8�
����ß�|8=���F�6�<٥}�D����$��4bs�����i,gjn�KX���RjMf�$��l�m#�tz���N~y��
ϧw�a���ŁL":��yG�*���������g-�x҃����<�Rk�2+
�;�̒�섐��pr��A�ƥ,@�r��f\�O:��Î+Ow6�O��^�kgd��	 1�)_sH�Xn�嫋4��OD��JhݳK럱�Dm��KZj)���^����_
���k(S�;��c�ض�
4Vge�W��un��ì. )�v�g��|n��	{qΝ��N����DHgR:��TҶs�����Ȃ��#��؎s���fO{�2�����m��LR]ҏv;�b���� ���j����������S[th�2AJW�Ҕb�#�����ȃ������|v�7�}���G�0c��H2�mdsT�`F�=@*=�&����T��_�l�ur��קڬG̃s���g�J�����A�Z�j��������O�꿾��-�W}��C� ���z�!�����I��U,F^6�s�C,��?�W���g3F'*��Z+����G{6��>yv*T8�8E��9�Cz��P���H������X�l<�8��+b1�%��IA�A�3�F	^x�݀A��J/Ծ�tux�$;�zҳ�"�B�������#zm��љ��Ҕ(���m�+٦����_! {�B8&����q�s��]ɿў
*�k�< Q��uG�gŇ��j�$�HF�(=��>��z!�d�`Y���t�$��RX_�(2*Z��{((�B<���mn��ϼ%�2��D(�ʆ�e׃�Sϙtǋ�z<)�Nt�z�Z��2m����k�ah��V�N�-��4�W/{n�t)��Wi�����J(K���ï���s�j�iVMp!!�n�w�-rgż#�uW^𗽥qn�T)hu�kꤲ�L��v�!j. :�Iex��c����ż ��S�"I�g�W:����?��2�?k8F!3�{�S�R���m0]4�E���pC�ơ@�THD]�ڋ�1�߁���2�dT�!T$�l��p�Y���
�l����yd_��z�}�V;g��ǘC'z} � ���H��\�*id����J5Q�Y�P����7g���Yԛ@���}d�sٹYn.4S��o,- �k��w�zb�v&���l#2�S�����VE�����
H��W��T5��Y�I���lTb_9E�&R�a=��O�:CF�EO���f�y\�OQ�r��+�Od3;���T1�,�?O���QZ�q-���#����a`�Z9׊����U���Aч}��ۈ��IΏ�4o�>x��ɥbg��+[> ��ž�X®[d�0D�sA1�<~� P�)g�/�4[v�=����6q,����ȉ-/HkPm�&5��>ӏd����l�rə��}���m�S���mc���_4��/���W�I�G���p�;����F/�#�NU��95�<�O���5~y��y�l0�㵗=fn�VU�f�tBi�l��u@&i[�W"e�|�ڧ1�
��W� Kz��f�[g�I���s�o_[>T��w�|�#=�`럊��Ș����
���x���Em���.�-����m���\-��fA��4h	J�6�i�5ɘ������Q,_�?@t
��J���d�y�fy1�X�������S|p��&es���
���_Sm��� 2i^N����k�Z`3�/D���if���H���dG�ٯ*�}R���������C?9��G)�A��"�د��͊(MmM/����q�s�A��D-�
�&���PF�l����|O��c?�o#�b�>�6�����P����vF�P�,�NU������8��ki�)^/Ά�#��;ƴ[77�0��^�{�����]�5�������Ij�r��i��+���9��;M��xl�l:}�6��R���Ǡp��U��-��`}|	�T�� (}fv�{s��ILA`N��_,�0 ��&��j�8]ɿ�׃;�c|��p��~*�E���!2�dZ��zK�	H�������^�����T��)�����+^�z)Ќ3�$q�Sr�P��tv�^>~��x���$hݜ�1�(�4S�MW�-	��l�IFk�0a���m�M,������{͎a
s��:v��_���A��H�N$5,�%��t)�G�i��s ��wx0`���D�9��o��^莑��ko��L~o��'r��+�I�!�s�Ջ�1.�^|��P3�{�l!���P����4�8ѣx���������q�&5�Ʌ�\m��jp=Yb�$�)Pх)���*dD��K�5���y�x�iƳ�`�83�.��s�x����2�l�X�*(�󭳛��@f+^��Ak/~��mL��3�cO"<�F��2�jL>ṞY��w�7sG3�E#�%}�'Jr��C����V��x:"X͚p�>����C�q^ևh�8s�\5^nPV�3������'4{X���ܛ2�p+n���T-��$�N��E5�k�k�
el����K��h/��O��6K*�wϝ�B���(	|���Ňm�Vs��hX5��<P�����U�N\�����}1�k�W��>�+{YX{�\P@�Vsî?��=�K�,y�/�')od������G�`T���
���� ����]�y�2T��lA >�O����r~ޖp��!�@e�_m�/aK-�I�X�� �Q���ad"v��Zd[��T���/�с�9���h�M̝%<6|�r�9D��� =C[P(�X�"wqg�;�q��DD�S�#��Tq?"�ai�	�j���GV��i��c���^�&���4��/��ÀQ�j�����0�H2�6r����}":��;���;?d���|��,���^�N�M��ޥ#๠�'oq��ڵ�HvR�Q��
ƚ�B����p���"kӧ��Lŋ��w����<���O�_�GC��?�L{���M���ʫ&�Ϗ}G,�F�vd9#
����OV�YWOB����� l&��S?�nێ�&tu_�tӮ���}����.:&w�Ḛ̇5^��rJ��F����>�1s�/�Fp)�Le$\�D�����e�$%��@��~Y(_��la�./�k��Sa��U�o��<zD��B���Z}H�?6&úMV)l���[pݛ?���BA/�|�eQQ'�����;� ��� ��\P�����x�C�R�sr���?)42C�S���`6���uA�`�ɵ�B��}	U�r�3MJҞc�y���u!9,��2RV3�E]�?Ūb�L�1��O7r=�����^�'�<7rf����#��.cv�����rᵩ��?N43��7�YߟWJ!��.]Z}���-\���L�%��@�Y�� >�S����H����aZ����.���Y9
-�neL��d�qQ�!�8�E�����*ޑ�̐CFG��[P���X���%vA臭L�T����b��q��Fd��'_	avO��؈ϓ^K��=D����Ѝ:��(�=(1�����4����O��Oś6�`����a VϵV�k9?�0�iY�Jo�hw��_���b���j��j\�(c�`�3���7�;��G�"B1�.�J�.z�(���7!Oګ�m���!�ܶ�@`ˊ,\Xwt¡��ʸ=vF��wsha�T�9v)`ЊS��\&;���>����ߣV#23��)�qB����}Θ�2�_<uL���?�'�R��ץZn0��iW�_r	�:���L�Մ��~�ǅ,z��h!��G��#dhg���(l�t^����<9� v[��jؗ
�J��y�԰��Y24�%�t����Oӯ�ˎ��N��%$۰��k[��}N5�T��~�G���"u��M|�>�.Ÿ��s��"zѢ�M� ����n�Z��d����G�޾wc���u8�+�`Z4*���5�����ZcH4��A�^k�(�vj$	�P�]8�����	CrT�k�
���M�Rh$��-��I��C�0`�Lc��HS|P԰sp�W�w:_Ui��E�0�N�`ú�����mlT�bsw&��'A�1iA�#�$���H�lP�����U�`7$�y�0@!tM� ���G��A���5Y�1b�xXN��_5�<xT��t�E��b,���Aa�f�,ʎ0B�y�.��/h�*��KD�(���֧�A���AŅ��2�B�6�#b��< }��J��m����Ji� ���|T���,t�3����O����s($Y�Z1�(��L��mW��̰�Ͻv]x�n�Bn�o��C�1y�9T>�5;W8mr�Y����h�(l~�r��mk#ޏ�uG��p��������2��/܅Q�/v?a`�n1����b�i�:���J�;1ń!�oDͲ#���e�cxdP����^��P�=d�Z�c*ʩ�u��}�D��o�aD���v���X�R�e,��"����L�~��'NPwT�0��.�%�Z���y�=�0m���o����;����i�?S��J���&��[�I��M!�)
�uܜ�q� �g�u�K�	7�:}d�'���N��"-z����In�,��d}��+�X�,��[���G�WK�Y��存p���>,��x�#���BD�8��!b{g���(�/��`��DV"��(�%Y^F�:P�AC���5��I�|�W'm�������!���s�k�ίI�%@")�I��AC���`���"���?���[������5ld�ު_�[�3�r	���9┊_�i�(��)a�>�O�?������-���-}}��7��(����������(s�a4���o$����m���JV-1�#��u�^���o�e�U#�v8s�������;/�p�z�`	�s�VJsXo����=Z��SZ���Pv�G���J0���ިrw�N����.�%����m˱�/�H
>�pv�yt�K��:��يr��%-4������ٴ��-_���!�)�)��0$����~.�P]
p�p��Ö��`[�1Ÿ"$��]P,x*�j��,���on
#���$3D½����囔!��ь�*3��y���Rq��,���)���t7�8_�⚾�����]&����~���Ⰳ��o5���/�3aq/���ȸ��Go�3��i���Q��!�(6�����s��M�+K a�垭m��Ͷ2ӊ��k.�>=���=���[�^�7���5�@@��@[��e����©K�Bbܧ}��&a���VF#B�پ_������:�{�قY����Jsz(���df��Z�,;�̫��iܯ�3�R��̱]���������^yMXI�1�pq�>rҎSQ�9)FK���-�1����r������}p:cj�W�o6;㢄��U��}�k�5: ��L-��~ۄ�!o��|��˕�ނE�&����6��\���8��������RW��f3ݾJem\�P-�~��Dڋ���C�f����%���k�u����>e��Dˬ��=��T��j�+16�
o1_J��U�V�D\W�����R}��i��4����qrD�9�8+��j��r��wSuv����:�6��b��4v�_���kZ��*D �Odt���E	Y���q1u5�f!�w��`����ZS|d�1K��LP�sr��	�C=�U�q�F���E���LhT�*z�\d���oLX:;��������I<_Y36��8�������o�v�~��Y�j5.��L9���ݳ83��>�r�0S�霄_�n���FpA<͍:�I�U+��ӎ��F��̛	ώ�{��j�Ԫx���*[�g�j���㮥F0K�T�m�����������z����u�N%��'1$IFK"���!��ګ�E�3��N��^�v$��P���v�o�O`�'�Vo���(EQ>ў���^d:��X��m���r<�+K��Ԋv�&���@!D���halk#��U�;E�i/=N����\�B������+�9�R :O$aj{�����Ȭ���� GB���һ��k�����3�ށU���3Q��2𜽤1r��5�������1J�|7�Fd��ý�m�LҠ�g�wҺdW��Ĕ���g�H�q-)b�k[H/���k:++��I���5't�G��O��H���5A�1>���H�7)���e
,XԶ�����F���SC�f�UA�߳�1l���:,8�1͉I!�mO�0D�u��Y�l�tT�ò���J|PՔ@t|%��»H�آ��	^"�U�A�߻k�a��]��1�_����ח�-%J�ӊ5e���n@8�Y�iRz�G�<��7�Ҥ��)Cc����!�~B7[�%�?S��^/�䶥��w��ςM6*����9�������'�6y���8��߭	����o�x	�F�۫���g����	����H�h��5])w]<F�& �k�G'�K|(��nQBN����U{�n�EyQz.�B�� hH���.Ϋ��=�|���W���ZAR�2�˕�6&tO�)��O��jw������ �BbusД^��0x�[�P���%�&)<�z5��������p�_������J�r�|�!� ^��%�E=qqnWN�bJ���e
bφ��+���:(
��,�%<á�)KA\~i"wt��^]�&�r9I�Ȉ��"��o��J
$fё��g\�$�g�7���|l*������*����ܸ4�~��*�Nn��/IN���ў�ϭ����۞S��L���BL����o]�����	�у���+8<噍/��u|}fc0ƾݑb<d21Q<<���D�`��2�s�����D��|��I瞴�gȫ|4O����6s:����Ǔx�N��`E�������>4^j6�޺�f� �I�oؿ�7���N��@��7��<�
Y�GT<�y�o�c�U�wՖ8f���#���ܮ#�4�}���{�ἇI+��aHT~���+��ľ��"7l�_T�	�H�;��6ZP�2�o���;�kKAOE���>lV�x����XX��unK�*M���5��P�:Oϧ�m�΋�s���4��c�W���)�&VA�2ɓ�V���WB��֜��`{�O�O�]��=�d��G�C14a=�P�0Ն��M����7�lќX�\ ��ٯid�������1��P��޼W��@'6j���� ��i��+�<dE�)��߀,�Q��h�>�����Ā�UAP%iau���q���.�M#������}6�Y�Ú�v��OF}'���N0������2�ky�8-�~��+���ur%�#+5�Wc�_b��6�=>7޾CV̹Q?�V�R��t���~X�*�N��fv�/��
l�+V�].g��r�7P|7���>�v�a�D��d�����mgO�	�IiM����'$�I�bހFܓZ0)c��$�1 �R��bG�Ƹ	?����,p�L4�xec��\��T�<[�W��g��m4���NG�A�D�d:�jȐ�Yӣ�o]~6���P@O��� {W�U��
`~�0���I�if�X?|a��P�gU�D�M�)���`j�\�,;r��uI���~��Dv�9x��L�YN0q�!œ�O2x��A��4�ov< �_ȁ��jNz����`@X�2Qs5ˤ	N5) ����9�YߠV�+g�8��M��
��yJ�B����iи�D�4����D̨�~�zոJ`���Z$�����L����c?!%�eD$��띖����9��D��l���j��Ō�Ѫs�O��uM��}�r�<�
�Ksh���2yд�.bp��C�C$u���y�^�O@�DRh�g���ǲ[~��r�I��#�#u�9���g�6?�^�͕�m��"�L��]�%3�jUc{���� Ȁ��;U���9��?����;-Й<�h�`�ی������At>�X�8ހ�K�2��z�����K�SfG8G�:2GK B3���aN�B�J����au��:AK(,����ei�3x�g���w)�j�X����4�mEVt$�pu�iE�������;���I1�W�uf�+����x�ϕs ��ۘ�SRPG�Z,b�,��|�z��v�I���C<6α�j�_�G�{�B��v���t�- �`�i��w;�8*���?����޳�V�n&��"����p�i�zX�0�!��ɼ�������{�M̖Ifz���c�� ���{篑A�Ӧ�S��D�DJ�MS�����=�FG�	�3�5$��}27KY�z��Y�X\.��g��m�c�1/@�k13<�-���� �	���]���7P^NVYf���r��	_hN��TŴ��q�:�������궳ͪ#C]NG�B|�g��>W�4{�y��r���5幤W��ёÀ4���'�෨o�@�/xK\���p956/@Oj!���jא�I��-g9�閱)�+ֻI�X�[@�^��O/DҲ,��Ff��ks��[َSu0vg�׋��"l��+�K)S���bF��VB0��	I�k!�5�oѯ����d�4r��8��7��y<!��wy�gQ��=��<ճ�P����\��.��*��=���I
|=X�֦Y"N=Xe�ӣ���� ke��-�]u�Q��E:;��I�f-j��9�5�PlB�85Q����g����l���6E������
�A�V�F�x�]��oè�_��-���"�0V��ȳ�m/�tx.,��n�vhU1$�5�?
�)H���ˁP���M��i���#g<��:�+���L�*[�7~��:q�P�����n=��x̟�/��S�����tj���"{����1ja�����DË���ֽ����[Q����f`�Y'4���\��].e�-Ev�Sk�y*�Kk"��)��@�p���4;ӟD.4�"���������<�'�_w(��N��n�x�t@��iA�°�`��}�P\"ڈrk�Q7���oW�L���q�9���@�Bo$�/k���m�.֥�����眳���/�0��&�Z��4���8k5��^m2���Z�[�[2%G��&�5�q�}\
����ŝ�&y0ؚS�����^dV�V��2��`W�����N��l��g������R�>�D^�q�jL�)틦�i�3��mfiXu�*��p�[�W�}:{[v����g�J������s*�U>�f��u���\�V�����^Z����(\/�l�z�� �Z�Ɠh�󴥭Ya��w����S�O�[i'�T5��'�^�4}������]�%�&"��с<w�;��j\�(J� �W��뱜
�iH܈�4*�f��4����%�u��Ž���Ӎ��Q�}S�?�\(���ڪ�a�}Z����<�7�MF�ƿصnv������rw��ધn���Ԛ��6�uΨ�PR{l�'�\Wfo�Q�}�a�_�^t�ò��z���f~2 [��n���ӛ��fb�y�`~�:#�ӧkN�FT~H�z��g*����AD��F�w6M��2�J7v����^V�Mg�ϫ�gm����s�}LJ��?|�xQ��[��×�j��׊�*��@l����iN|U,�vv�P8i�v���o\����Ll�["�`{Z�ހaf���B7��,Z���@pȳ6��"�-�� Q���=|�ղ"<���4�o�Ku�:��d��凊�݌�¾�:�>3Y�E���?a��mB��Z�F���~�F$*��Q��H�A>�i�k:>���;�Q;�آņ�=�Lژ���f@���Y�v��!������CY�j�!ǟ�w9J����=��]��'@ӽ_�3��BHg)�%��Й��v�돭�@>)�H;�%� [}�M���R��GX�t�E�I��丬�#|��o�g"X�'L�mڠ�����/�Ɯ�<�Y��@��6�Q<�S�l_E��`�G�GbaZO
Bq��(�|�h����.��]M�I��~��3���79R��En��zã��G�jW���{E4������� �T�/$tD^�$�����|�sWJz�����5���z^nY��_�:�'h�Ŏ��Ah	JQQ.����f+��+8ȴ!@�kU�y\�+/ݝx�]l �.=�?���IOaV���?�N(�zZ.��<)5����ǡ>9��P戧㕡n�Лbny% �u�������
j�\,�7����Pi�ۗu'� ��a)�|>@~�}d�w��O���2���_h!�Θ�M#p�s��	z�`-}�KH��H�����s��dbe4!��gK<j��j=}r����љ��D��-�j$�����6�j�4��,�$�RE�s�*�qۅoFi	����z��	��0��t z1�dܑ:س��i�L����ja������Gr��g�(�kK���LT��������u�Q:��6�y{w�.�:�"Y.%o$l-���q`ЍV4r.�±g�+ء��	G`8�,bp':V���kK/ї0�m`�
�p�;�R<�I�k*#��7���;s���8�p�V����`6S�����\"���������kTJ �>�, ��U&�U1$~��F��(�Ϋ���E6��U�t���-�b���40[>3
Y�R^���Z����Z'��{9�zL�8@_�Q����g��J����6�RT���ub�B�f��ٿ����4�y#�r왚���$�ԙ�h'�tȕd�������',q��a3��Raۄ�k�n�x�j8��}�քN�w�H��%J���W� "@��t�j�;\c��ض�ON`��|H�m�U�f�O7&aB_���4Z��?�%��\�����^X�ε!�~��>���XkjV��Ur܉WC7��F!\�j�����⧸�0���~����
�K��+��Z�A$@�q� ����Q	 �7�t��C!�v�ƳT��],f$ց����]�q/�S4:�	U�k��*^�`'��s���W�H�8�Ri���E�״b�+��6b�!���?���-K1���_a���iIig�! rJ��|&�]�f�U�p6K�Ҭ�{��-���U�GW%К��A�='��_ �۸��<q�]Iط6�����=}��<��1���gс[�¬�J��7�&w8Y���[oy�៞̎�c�A@��_j��xN���f�)��ᔃROf<�Pٞ#�vٮW+	#�v$��X$\ !��Pq�%-^�G����Z=;���B,������R����ȵgZ���"����K 6b�R;3Z��ˡ.N�Ҹ�;�A�Mr}�_��I	Ͷ��Xm�Ҋh�kD'C��gpSBZ�#uWA�)�YU߯c����x8@�JLˤ8;M�=�P?�A����"BaD�M�wcH���1+o'�E������ЁN�Kjq!3я8Fg�U2�|��Dff"(�ͨ�gy��s�R�kݕ���$�~��U~ .a)���ᰊr�T&/�0қ��sE�&��A��r�U��to?~� �"�E9�6�^��"��Y���]�p,b]Q/���5�B9�z\�^$p�7%7k�m���O�՟��)��8fkoa��4���"�Փ�d�Erq�y?[�յa����Ǘ_�L&�ĭ�
�T�FE��W��f�&ʓV��7�S�~)PI��|ߕR�<�;
�gLZB�mǙ���m[!�VE\�!���my��ĉ����,��p����B������@�j2�K��#x�_�i*����iCB����OL�g�	��O&s;Y}	�6Y�r���	�|�ZH�Nǀ�.]n)��:^+�p���.�:{Wu�}B�$� ~�����ٶQ'q��邐|�zT�kK')�#�7���!x�@�k�zU{#.}�a�J4�ֵ��Ï:t{�Y�NQh�]<�l&3�{xNND��9|{
� ���r�п��sÖ�u�d��b����4�iֳ����l�3��E�R���^��[���İ�C�]�kP+~&��0܀�t{��.���`�H=}��)�w�Jљ�Y�Ҟ�g�=�ma��/�6�~��Y�FJP�
�Jڹ^ffQ h�'�=�d�Z	?Y��5ҹ6��c娲�" �f�J���y��L���z��w��G]js��Q}�ݻ��R}J1g��������V1�"�;k�R(�b�"'Ɲ�MHl����]N�
�z4U�k(��Zrn9a��F!�R!�^�'e��n�W�!�bZҧj��]��~���SI�,\�2���T�[�`�=�B�\��7
K=�S�l��Ⅎ�$|�:9��k1��Pz�So���ZkH99����o��ק�O��|�*R]a�C�4���y�f>���u����S�X�Gʇ�N�Qp�5���|��6D����6oO�����hn�z`�e���vGu*��sI�4���)��wM�~ǁF26ʩ��|~�F�Yڽ�3X/��|��,�I���j,���`����v�V9
��+W+`T]��t3��["'թz�2�a�ܶ�9&-W�f}�؃(��se O�}|_��u�A�v?�w�j�5�ͲG��c���K=xm=�j]EWÁ�}$�_{>A��0�/�Q�v��i�g���M���6�dp�W`�@���~�]��M�� �Y�r�ơ���F�t��>�".x�0���断���s$}��)�+V��.�J~�Y�����2Ϣ5#�;��w-sE��R��tD_}~�_/���E�V�IA��EWQJ�%���9�~쭗3
�v���|^�\R���Ea(�Q���4�	�Y�T��:�wJ�>G ��͋�nq�?ӭ�àұZ� e��hA���)V�=���;�3�ͨh��'`p샅��a�0oᇆ=A���"QZ�ۺ�z��yy6��ݙ��|$A���H������.�3�{M�?��g�_���y)lg�Ys��?{xx��_{��oa�o�O�c
S���v��>�h�½��S�Ke��\o�`��"���`c�b��T�����b){
Z�,e�{��ou����bB3��{�������#V��Y�O��]�&Eb��zz���Wh.}���� p ��2?�%���U	��UG����T�q���uV^)$[�з�������-�����*;P*ol5����H緦0ᗂaWAe���$���Ze��M*�Va\�)�Rp=%5JsP��Ơ2����5��=P�Px�_z��y�_�=�����F�H�:_}�'نR�r[X�����������Cl��KV��Wʬ&���y��)'9�0C�;��z�Q�֟k�n��U���!��P�2��p�B�"5�,���LFd��+g{]}A���Y�M�n��k�?i4TLo�J��9�a}f��'�Ǿ�~��H]����FSZӆ�%f������ ��-�VL�V=��z��e����L殛��5��- ��ʩ�D��-1j��]$�h�&�},w�"�jL��-�9��^��[l�[�&�@q�aW2�
����gi<^�jM-);kC
�x�O���&����]���<	��ަ(Ak?!UiVu���m�_hc�mP�	��8I΄��	��nڎ���R;ּ�0m�[���fw��)���W.��F�'�I������}���b"�nyَ,A�vUC��	�x��j��+��x�0�+�Y��C��?ZzR��\��i>�o6��*���(]�����,	 �W����c&`'�C�i��ʹ��U��m�� ��%)�TU�d+bs�o�4B���0m�aA�L�a~fN�9���,k�XM��NE>��z|��J`�Ʊ�{le��.=Z�8�i�+OW�VPݯ\}v����*� �h/�q����50��x1_g[�3�P+���n�fX^�$�& �wt���5�=)�q�J�U'8�=j��qHeS�+g��$�o�4��9���l�1�t��VFqp� '0��8�t\������rJdS��:�l��-�)��Lۯ`���g8�sa�n�s3�z�uFi$�~i�3 k��z�׊�u� %o��w� EeZ|̏��.� пҒ2ԍ�����@�\ǀv�>�4[#e���� ��_��R�A@�r�p�2�\�$Dt�*�Q�S��è.&#Wpw:j��u���n��0�#������?��s׺�͓2�G]<���j�- �����ۏp~��R�X�V��tW6�2/�W��W��f�d0}�G}ke���T%�7ab*�R�~Г=�פڜZj�-Hd��թ~䦉�
�;�ʚ��,��E�DUK_��/�f+���Cpzt+ΗI)��&CpY�
q��a9���o$�dh`[�_T��d��7����}�}::����?�) ,�R�7A lg�܌*�m����+����.�x3w�LC�U�ʕ"�נeW��B�A@H�m��d�����;8�p��$�ڷ�x{�#�&��J�1�`�#����0EW��C��o�V~�JwG���u�S�����- 6�u�R�׎��p���^.�>�� 
kJ���׋3�b�C�7��� /���ӡDs���t��2�����3��Hۈ��T�*���PoN��"��2�P�d�E<�C��M�bK/��/a�K3����#i�߭��ɑ��c��10a:�n��@̼;x�jJ�98������c���q/�:/�I�B�&�3W�'DZ�	�@p~���>*�<�V()w���bKp�\���Nb��U�Q�N|��L�g��$�fe�Xs����<x���x�z���9���eΚ��q��D�!D?�ge����zU��r��"��!qO_[���T�ͫ	GW8,`mn���Y2���}	�u�ks���DN~�e]�AԐ*bNY�x�?�j�+�!r2�u(�5F�kB.�DJ6� �<)+�]�b���jNX7��UӘ(3�A�m�z�.qGx��5��w{ek��X;���U�|&7�J�A���a��� ���ˠ�i��A	۝���a${�\��v��yd9^{Ůz9[�ً�n[�T�]>5�ܳc�t�Crs�0+0�g�7����ӫ@��?'*��˱Ť�@�
Yq`v���*����L?:��u�A�,�1�8+t��a�$?�Io��}+mV<�e��nnR��t�T�C� a!;��ݏ����Ϲ�`I���*�F��C rշ���\��`��#�2v���;��ORu����8��]���3"<�VPͭ�Z�	��AzM��ӪY���6��$������jH�a�D����DT�nT���~[����8����q.��顛 �P!p%@�r��s��:���|��BA�,x��Z�WeK9&��~=O�[�p�������a�d�a��ݳ'�(5��8��uԧ��?�������G1ҞO�U��5��;���A���y*	�4�\~�bC����:2��"&���j��b��>�T��T�aOAvx-����b�z���-jD�!0�TU9%�< �?E��È( �%ű��&G�̯	�Ϡ��暥���h�ϼ�g$���^���9e�;�1ICq��jIRz�;7�fɖ�.��O7���C.�C�g���qB�Su�+�O�hM�7����4-��G ݝ��i]x�R�˸#?*	ڪ�J;
��܇լ��Q��X8Ğ�F��Ӭ4θ�� �ش�Sq��v��µ)KO[N�&�����z# �_��ݳ�g��*�?�he@��&N���_%�E��\
�4������:�z$�r����\���{M�t�f�������C��]�����8���}�ּ;�M��m��E�2��Eq�[�q��C�B\.ۣK�MF������ɚ��A-(n���Ș�B�235��l�C�����IwsY�h=F9ސ7X-�r~���`s׳�+�Sv���)h�䪇O���
�&![ÑcE�~�h������P�C�� OFJ_!���хM��w��:6z��`L��%��+����,\��n�P*�8�_�zdz	�$�O<j�x}UE�H���eXC�-�͘�Ɇ�������"�����VO�v����|W���£�2:���x�uv�wP\��ɦ�����z���T���L/��%�Qk�j
���|�5dw;:8���	rY��ۗ����·�a�z��z$йX����B.��)��8��S��A���(���h� ��oX�NȰzp�ķT���!�N���(�Y&��o����~��ƙ5i���R��4h���Ϫ�܄ޡ�N#��e ���������h�C�K�D�U������*ZR�5p6���:װF��	�̣�p�YV="��p�0�4A�<�Cˋj	�t��Pԯ��]�΃��(�/��k*~�P��Xsݴsq+=�N�s�ѐ�mu�h��2��ʁ ϭ"�;Z!��Sg�w^w�:|o)��H���ȸ��;D�h���H���ǯ�R#�\�~<ɔPM�k�+��G\<��o�ͲY� kGɥ�y��*Nl粁�sĹ����0�<����5qx�qU1��B4܅��{C!g�8���,�F�w����WW��>��o!%ᯰ��M4c����emek큛����j�g"e��f��Y��
�98�a��Q�<c�+�X79�$ Sj������Z cx6�N�z'+�E�-o�J ���#���Ʃ1�L��~�;�]s��\{��������B�՞P�?�Щ���>������if]em�&��V�:n�B(��ܤ���D&0�K5��a�R�'cʜw�#~��g1�ᴭ�`�9d[�ѩ2�Iz�7�gF�W���s�9�.�'�:�0U�3�����>aU�s�b���mlp�=��ǀ��qh؃Q'2F֊y��k�WaE��C�Q��A�����;$�j0�v7��m��NZ߂\[���I�5/%��4��jҭ�ϯ퇞����2��6Q�ų�0�?��u�?�<��2���H���f���F�� #��¹),,�e�`e��%&��jx�o�Mz 1ǆs���[��z*������#�O�+���s��!BH����أrl���J#��WY3��#f��QP��H����2qSҁy�:_���!�ɢ�u��&�H��_E䶭ߍ ��W�-��+u \n	%%Y�+[�Ύ��猠Ǧ Yٹ�g��R�+v���ۃ"#ȑ�A���d-�?&]����1�nD�E�ŭK�=��~[0hg�g��P�y�b5e�����i�'��ՠVh}b~�
�A�f����Ǡ�Lxb��+��UN�=8'G��!�y�ukBǂ�p4`%�G��W�Ј��DO��PL	%�c"A�I�j�ue�W_����c8)ʡ��v��%u�V�v�ł57�Ir̵\?����8�2�
zk�Q��ѿ�F7Fs1�F��.ad�N���Og���q����������h�H.�٬b��?sm��Y��4)��C��&N� hd�9 ��Ϳ�^�+�~uBP$���NT=d@F�Ÿ�f���vty�;���*�-�hw�H��~� �!iA���U��F<;�1o,y�:}z���Y${�xߜ��QO�@�&�cs/Xi�Q�~�V�^�!H��E*�{�O�@��d�8�����2M�j0G�Ϭ�m���`Pm��>��a����[�h^���ˋ@��O(��5-n��\'=�(ʭ��f�� �X����z��z��PDa�й�ܘ=�Ib,gR���A�q������x;��%����o*Y1KDQ���K�$�-\RWW*/���4:�Q�c�M;l�-e��=�z:��u�W`���,o��(���4���I�_�MM[��}��MQ
�k���<���G�.wd�d<����2+!�������\  �;���f�U,���zd;G]�9�u�|�O+��Ꚕ�>�����6X��(���0ݹ�Sn��G�[4��ݩ(|�� �W�*�L�K�K1��Xy�I��p���j�P��B��be{�9)�~�H�/H�Z�c7+]�@&?�����������DJ�VӘ>Hd�y}�a`�̽��*"���ަ7���,s��WЛ�vf�Z�f�߇l��ZPv��Q�;1uN�y�u�+d��uI�L>+&�3�VDQ!97��������S���+���^�� �3D��"Nݎ.�gJ����
s���y�����jZa�&������d��3�e��x�0�T��g�����[-
v�|�?�k�7��Q!?���K�~���$e��c���b��+x�z� �v*��̳»q2�F_�!�@;1���3�E�I�ފى��~a
�������d�bݿPU�]=��)�n��[���][ Xl�6(Cd��\Fʤ�P/��Xk�hF-�1�^��0m���W�ogp��s�[��F�Y�ؕz�x�2m�ed�����������VZ�=/B�v��g��/cA��T�Ԟ�G��*����z0mCu*��>�s�xvD &#Q/�<[gʄa7�����{�X�ڀ�5�KZ�̖��5�/�~K����0<��ZŹ%������<�-h5f��C�.&��U�bg�?�D^4\���m26�.�E&�u�Rd�lGo�+�̍�NN5��f^`����+�*f?��*Uډg!��?{1����� \�3�s����H��"E�Ȝ��*.h�Q'\J޲%��GMgC_4�#P�S>tE	��8�[�+,��?`� 4��]���_&ƣ��R��B<J���ha�Ò:��A���ß�O�����T�m�i)35�z�1���Y2 ���Ia�d�����}(o�OG��Ep�)v��H +��a���nCf)`oG ��|���H��6go!��]i�Gr��oi�|ت��7Ө�i��9��-j�?�1hI�����*����xz]n4Q0&i��!+��Z�w�1^�[�k��������_�O���w��&��ft�bV�cG�ʕB�h���tud�-~'�mG�8�?o�Ê|���P8��q��^��������@�b�jL�$����F���{ECsI�Y�=ߤkk>�|��.��ְ�F�:�|�/T�Sd�@�
��<�5Ύ�$��)��zk��"d
f�:�bm%g��'��6�/�7tP��?�Z�)�+v�|�-;O%8hV���ƪv��{-u�|\�6�ߡ�����Dlh���9��a*��[�)��z�3(��h����x���1[j4�^^���`ۄ��:��խ�;Pc��/�^��w���¿t�A�(	lO����#���
􄼲uvӮd�'�Ψ��������m((e�~�Mw\��;7��̦�ρ2'���g'���������b�ͬY%�*[�=9x%x�I\R���2�l�D��紁�s�]F�����W�ǔg��㍘���ڃ�>"��\����	�e'�5�<�[�(AJ�N��-1l�7����W�Xv�	)E(�&?�ן�6�[C�,R%�D�:�'�>I@�%�/@gW�x�nR:A"��e�c�;�v�����M�6%��T�w�����\���(�|�ݫ^���˛q���d�
��e^��!L���!t!�z
_�4��e�<�!d=���@"�HI��{[�x��NB����#���:�G)��tp~��D`U%����&�/,��˳�2Fi%�x�@�Ǎ�q�>�9rG��S�������v�R���*�mQ|e�6-�JH�G�jv@���n�.�5!x�];d
������
C�0���um޽4���G���=�����p]�1�Vb%����g>�	�5Ig�f�=Z�>J*�
��&��9��Ң�k[v�߯WQ��YS��嚞�Ȳb�O�G�	��#6����X��є�d�M��1E�`t�'O�<x �K�E�� ݓ �̫&��qZv��_)l����ب�bn�}��M���ْ�� '偢S�!�&A�P��땤
r(��J'���d�K�~͝��1�����o#	��չ������B���t�y�,�?��]5���Ɔ!���82��ȌZ�\���&�^hG��Yz�|�K[j�u1wG��T��l���#�O�Z:O�A�@�@�+�N�;��h���l�J�D�}�	%0a�[e&a-�h8��+���5����d�����7���r����/۞v���b&��+�%�b�˄�L�!�92&����5�����z4֭�!���߷z"v���\�
��9-6��ȸ͑��ˆ1�<��E��J�w:�z�BѺO��~��W��+է|��( ��Y%�$����M[�sD?���a)Kr)���\]3����|؎E��������p���&��ٳ�8IXo��!����`�ƙ��E��Sh1�9�D�&� LeفP�Y�F��@�� ��z�\���!9ȭ�)���h@�?d�r���x����"�*^���OX���/^�4�q�
!�y�#�u4?j��TaN����k�xe��Ѩ����b� M��(��K[�zW	nM쿚^ERq�x:���<l�aq��G��XI~/���/X\dQ�I�N�������熌'=z�C���6��Fӻ�'�D���[���V!�aGS�����s
�裲9�R|��6x�{l�%�~�<f^��'\{[V�� ���ZK<1w���<�%����Z��ȃ!d�Gw�<�ðh�Wq���3�?�-��4(G?���#: ���as\_��e`r�9�Y�' a68�:�#�ԝe@�k�W�Ꙩ̠ ��H1��y���鿝�`2u�������z���Y>�yN�)o�9�$�Zr���1>N'n7�*[��;"�'j�av�,��i}����W�#!�����a���RN��|�F���#0���K�W=��=0��%�GU�q�#�>Mcﱡ���";�pxġ�1�/<�2S`��9��/#�	E$c3�Ob곃��5ڝ��SNj�����%l�_/��$����C��<��x���h!��о���_X�?"^@�6�\���k�;�Y%�
U/Y�k�����hyӤ׏�$��kOΑY������O���p�D���WS�*���PgUvdZ���"=��| �Fls�K��ʵ_ψ���=��8�XBQΞS9�&���8^�4��+��*�>�Y�p�HpZ��mX^zO� 8��w���:�_S�2��)H23#,+I�,4"����@,�,cVc��L�;h�U�҆VV�\7:�yjG�[�E"�Y��x��e9������	��KܪV4��Z8C�)Y��~#
a	���s�A-�OH���?X���Q���~糣sKQ��Ȣi@Z[�`:)亖w�Ċ0fu���jJ_K7��SF1�Dm���.�~*A�̆������6B�N��A��*��ޮ���q�+$�n4���9��dtgNOô�F����v{����s㱏>�h��6���
K
��ԉ+"��c���T��>���8����s=�CiQ�s�m�R[�(��+�(8�@��U$�
0�����,���D�4D�/�OFkV����0���������:��$9Aռ�@�͑c���i:�"�t���T�2�odcs����<y�J�jLi�?�7�**4+;ʂhN��BX��e����wJtyw�1��k��ybvIxd���B�T�e��lڀV�	�K8��<E���<m����;����h�U�cW�-^��/B
#�D��ئ�f�7�U���Y�b52�l=Ĉ-�����Uf��VF��q�B7�q}�$����Z�� V�BHH��_}��cK��g1��6�e� �W�#M|��Q+2-�'7/�
�
XZ(2��*rI�D������_���ż���2��/��a�r@?�'�H��1��9�g�#��
���R����FW�T�T�}���	�'���|��u>%�knT����,��w?^��_��j��{�R%<.d3�7�s�}�����n|�����2���,<
�H���X�b����vh����w����o�!:f����ľ(���rr���BCO59d���������e��v	&h}���K��iW9*Y�xqDB��AЦ�>`�&��xA��t�����k&��S�F��s2�>Q�Oo*%\���c���^d-Q� ��,���
�/�8��r�<*c����]��E�<����{�\��R��6�5 ��s�z$�D�ras�������~{
dѴ���r���ۖ��tw9,ʶ��Uʻ���r�CE2n�Fŉ�$�L��J��Y(5OsJ�s��|}q���gQ��Xꀢ��.<DM�Qy����U�?��]�4���w�r8Q 1�%��䴱D�uF2�Qc$Qp�R��L�Hs��+�y�pߪE�hHnl;��)�����&�pKˮ\n~0r?lR��0�~�,����7u�K�$����Q6eiN���f�żR~��&y	���F���4���C�����=sy�1�P<�t�g~��51�!<W�
1L~n��q3ȴ6�Ge�^V�Y>M�֩�ϲ7B�i�"j����N��-��8$�:���Lv�T�����u���.X�KT���?�?�=[.s���8@]�}�z���o�ʌ����^Gp�#���X>���B���?�n��ؼ���e��a� �l0U��mbJKE��j*��J��;����l����D��ԩ��"ַ,<:5�>��~Uj^p}���,�PT�$�^�X�U���4U�����9��������p�^6�Ⳓ�6*�jC�X�=�n�0b�u��9����H��œ�5ȝ�[nHd)5`�c���xr�ް���;8Id[��f���0v�e�JШ�)�fD��(ϭ���i��6��0�j݂%��<��/��֟D�KE<(�nN�̔��l.A��-<���+`q�^a̤q#�bT�4[�P�q�>~Eb
T͖���w�����;�
.���0>Q��I\p�]%�3����
��� U'�Ú�oy5�x�/E��IYt=>@���1q`�R}�7dG�#^bpwݵ�!w� d-QL
9*����"*/����Am]���֩�`u��mG���nŔ�S�D�/����P���Z4�k�LۄO6$���^���oMd9?�i�-��ݝ������������U�c��츮�K#  �<bG#�K�����(�� �4\���ncّf�zscܓб��?q&�H0j��ݏ�K}�Ķ�&�� A��7����B��@Φ� ����3������eG��+|�?��4Xrh�Ɣmy8';���.P�My�)�������݅%�L4�}�Xo[\����l�:��A���������}c�5[���
41��	����"��׳�ɌH�㠐�^�):ph���d��	�;[\C��W>t��L*@Ϳ%��Z�}Ђ��1Ӣ|��VD'�a8#aO���q�J�$X�GY�{��	������d�zV���N^A��Qq^\<�{���e���
�KE�%����� �1��q�`$j�P�m4�V/ ��<4ɑъ|�Q|��#1A�3���R�+����^�.���գ�b�=��xmϖ�9�P����q���E���N���*��4N����k(t�wS���hM�CXO����*�p$��$��'�:���<Bv���dޤ^&ǖ%F1>��JǗ��f�?NO�f�����k�P+��<�d<�k���Q�θ���2�j�sRX`��G]/�z5�)�lP���B8=�Q�$qLT������s��yF��dTH����9����f㞎�j����e�w��}/̰1�(:���C6Ô����I4�AW��U�D�d�U��6z8K���*�wU>L���	ʨx��*��KSD��t�JJ��ڻm1
�"C���V��s�ʎV�s����d�O�_��d��?�HF%ޠ
�LN�������.#it�席;�ݱ!l:,��w/n�j��>� ��Ydn`�x����.���{��3x�sl�Y������(2H^��}�/D�9&�1� ����q��X�����r�H��7�?Ӧ��&-�4-ٛ�m�[�2��j�Hflnؙ������p�9n`�OG*�X�:D�N)���2�o���a��-Z.��/V�F갍��a���iV*��M�5�����R��9�?��כI�����oڌ�F��o��[�k~:=OI祓���o��G�$�H���0'�� �g����Zܬ�u�*U�m�(E;�k"�[!�3��r�c}������ޮ\��M*ZU�)�X`oY1Ƚ��Ux�?�&��?�F�u$0����C����`Y��F��6�i/��b�q��,�O�Z"c��`��Iθ�ߜ8~V+��[��=�E��Ğ����	,	��R����w�3�\���H���ū~���(��oz?�/�.����|�|S�(G��a%�s:�X,���O��2P���v!Jl�!绁z�H���-�u��H�5ʅc[������S%����O�,se�����e�v^��{�� ޲z��I}vZ!q+U��ޞ�:+�'#,O?�R�����
/�Rܱ�{@���ՠ3vz+TR���b92E�5P���͉
��+O�2Z(��#�6��$"��J�Sߐ\�-�Ǥؗ�|����_��w/���h��);�.�!,Ɇ�\�R�"�ɘ�M�����ںR2ڞ��A��H�µ�#C?8����7;�,%�_!���