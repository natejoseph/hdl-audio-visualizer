��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����:�unkw;n��n��x�'�J�1����,��p鈴���T>�/{7o�TŻ��Ӭ2-I�7��vܾ`hB>�1\$�$XG˥p���N<i�>-,�p����=�H(�6U'|	
^4�/\?���'�ر��|�@X uR��Gh^\�E��[Lg5��j�"?�=/j*�S:W{�tc{B�-�P'��!!�c���s �G�%��(}��Al?5H�Aa}ə#��JpH�;�,�ZÖ-"���4@�J�N?VG+,�1r.,`���������a�W/^���N˽��&D]x�Q��1+���#c��é}�HMM��n����}-/;�_�q����f�j�
/���$
�>��$/���-���=�{�lt��,���W�!���r.�gY�u�Ձ��� ��è�/�"u�ߑ��
r ���د�_�@3��)7��O��D��kZ$GZ=|7�����X����w��T3r��Y�O%�P#���`g�	�eT`���G��A����~�v�/�@����{�p¢j+��UNω~�"�����Hݜ���73�8�®9�94�Ұ�j瓦����^�a9��I{#� V0j
G�}�WNO*��t�d��޾�(�y��o��kw���z������u��?�0m���B]f
"g��n����B���7����Vٳ����z)�Σ���$|^M����pγgb���{��/6��# �����p���Y�NUz�6�
iΧ�%$aM-@����������j��3I���su_(_�\, 2�ߘ�K�m�H?���߀�n�\)�����P*����B���?�J��k�����U�U��ْ�<@ӡ�	��H�"����X��Zw�6R����H�X�ī�w�P^d�L��`.f- �3��H�3:p�G��䆵����%L:6�����>
��Q�	XG<u���8��"E|������F]d9.ĕ�$Ð�*�m�����{\��mH�X"�Kg�.�]���%�W���{4f�Q���U��_5
��
���%~u�xG�k͒NHn�ߵÒ���aXN?�SI�W$f	r$ytz�O���篓�q�ޚ����9^��R��7/���T�[
G�tĪ'n�N1�z*YS��TǪ~�M'B�\�CZJ�go�?����1�G������rF��������u'Z�<��6���-�s����ȹ��-���ȶ ��$Ժ�~�"Ê[�i2�@���M��0!�^�K�&@n:�����V��,��ﮡ������fPk�&��@B��!�m���l����/=�[�ն�dK��ſ &��^=��g9�-HУ��5��ҍ�|z��kd(��y�C;�����=H���ZD�<���D�#C4����c��!!nN`O6pq����� �E��(���[19�"�8��,َ��3Kx�k�g�k���������A����a�歄EHW�}#4��ݜ�5,���&��Z������Z��\�e=jϕ���y�i�Jv=*	Z(���w�>0R�\��gn`|ޱ�|�K�5��;�\m��٢�h���uW���z�������r����U^������̿(?���֮�K��D7Ů���XT���E��E�R [{����s��	����V"��Ŏ��a�7��P#'�Î�NZ�2�J���Vd�U���e��Kq�tf9��lQ� (�_�@v;/�2���I�3� EF}n�⅀�.F�9�%U8`*��J-�E·�{g���JY�G��Y搉 e&W�6�,��k)�~M�^ci���|[_~66̗��:����є�V��z���P��Sg����)����ǁ�@�q�D��Om9Gs�1��R9r޴�2��w6o%��Id��f����8����g�4�����@z�ݽY5�*�J�x[���v?����)y���نjfm$�/�3^{W{L2GPuT��P�a-!◾�d����;�P���k�Qrj�0Ĩ�{K�p5�`��G�C"�]y�Z��\��OY�x�Tϩu��w��W@���"�a�w�"����Z���m��+T�sC$PS���أ��n����#�wȜ��+`��,\8��J��o�b}��;�n�"��~��?��#鉮|8�磬eS��Q���4��������&Þ�EHs�f�pb��	gRv_�6������a��������.�H��Vpn�˅���EY��C��!8������O���N#�9t�in�h0�#�#�3
D��b�0����  ��F"���"ªM�����`���-�U�!BC���r:��\��Đ�Wv��e��z+�nUR�vH�k.�:�ٳ�]��&z���ъ<�֒+n8s�(��S�|��r�9ƶ�ɅRq:��q��G��S�S��CI�EA#�:�7�Ĕ���QM)�]���JG�ݿ�Ҁ��w�����1O�4���0��@�Df����� �ʵ�����2�XCm�}PK����q=Z&�$<��i$��P?�7�*����tUm��;V=k[&[��Yn��	y�! �=K�4��2]�(\���:7��`���($!�+���O�lP�s�gcTF6Za�~PN?啬�^��R�s�� #�ڵ^X�5�S�Z�J�3������I�[��0G&�GCU�^��<~�%A���M�x�5�k�*]8^9"h�pv*��W	�9��SuK$&���u'��c�ɫ��z�Cc�R�(u)�����\�Ŷ$��pC��<s�ud��eֆ׵C��>�t�ȟ��zj�G������+J �x�<F��A)n���&��
fqCY���)ry�a��zS��I��� _�K4����z�r�D�b���p�_���dCG�+l�'8���ؤ��}"�.ϊ6ۚ���||���)ai\������>��T�I�H~:K։+��ۄ9���u)[ ;�Ce����ekR��'4� �m�>p�T�fԸ�h�8I���2�@�XOD35�kyj=���9p�ߑ�{	����Y,C=P�~[w��<�~�&�Q]D�hW���ĥ�L���Sy�C�,���@w-V������LI���aI�/�TD�TGNa'��5� M%��k��r�Lc+!�\�[�]�Q�W��$d����}=�J��GTȱ�2��w���0�9�`9�8�-�[?�Xj3v٥e����T�	.������� �a�Y��ke��o��u@gDz?��ޭ����^F��M���|t�����9�_���"8+(w����-9:�]Nd���H�T=�ז�6O�
�6޻	/��~�,���Y����o9I�22��ϑ��Ώ��Hېr��S���~�"�ẍ�]��X�/�59MP��S����k X����zM�(1y�>����죷�e��>�	

�&<�b4��N�ͦ�4��,+E��|��T��fduV�	����	Jv���U3ӵ��8��/�ћ�ʕh�?���S�u^/n��9zD�%1
��Mʋ����^L��rD&L�QO���d�34F�U(����+&���ፂ��L�X\H�a;��Ct��E$`���A},��]�����K�Z�\𻟆��o�UE�Ɣm����	2�*���~m���L5M����L�l��צ��L�C|ء�Z�wKb�uRs��{��Y��w�����ja:�!��F��b����}���Ȱ7��� h�̲�9�����������Y��z�p���q���}@���M��V<���;`�B!�V7J���C�|2����QI&H�R�Ϡ�����	�{��7�ޱ#� 0Ұ����yC� c��u�3�Vϟ�b?�&E�@5IF;h��d��	�v�1� e�Cm$��3Q\v+����n(1�ޣyX�����Ut�����M��l�+��j��w��XD�0��9�d���_V���v$,�έy$��Zѓ4�Oayo�X!T��9�A���Q+Z��+n J�����p�-��}^�����.�ݬv��vwgZ]��c��2,&o���Šgil�q,����0.l:������l��%\�O$��O�H��S�/�R�c�a�zH���Q��������4����J�d�l~���DԄ&�1��$�S#�9��Z���R�����b
�56���GX��jZ��N�d]%�Ź��E�Z5��^,1� ��׽�__j���M�.m��㵺۵$� �01Z�;��k�1�{&b#�y����fF��
P�])*�0��9?�Ό�XP��i <�©��$���M_#�ݺb����fm�J�wP�I�������Y�+���"���'�q��䕙�:=j*�Mv�u$�xq���E��X\�#	�$�Q�. �/4C���2�`+��������=�X���i������]��"�]w����[�xaf�z�_�9ΜN �6�PY�?3rmv
��f;�R�:�Kbz�Np\��s�j������lu� ���6J\���7G��G%��M���7%�]�Jz���n�R����j�Ν�&�*���%U T������v��#2s�V�b��m`��(:���+�0�Z7���L)m�|q|��$_;��G;A��oOq��Uƈ�-�0����h_, �K�oM��*��q(j��M�fu��"�9�w0�Q	ڗ�*�%/�e��v^,��D���m��)��I���tu�^T���Xz8Pk�m6�����Z���P�7�ƪR%���O�7_tX�~g��?��*9t �iJ�v�B-K��Fep�mއI)n�S�XSˇ@���  �)	Hd+�rcMJ�бL���K;m�RN��Z4�'�Ii�hyYǴ��v�����Q�����xq��
3�_�9|9NW��}����Р~\7@*���F'2m��$��7��	��z[�y��u!��M�{�JL:+K�<��1~���Tt,��j��6�Uˬu�=M��,�w�*��`VO��5��Ɏ�<c��l���,�d�8 N0N��k�o�ۜZ܉�����ZX����F��"�g	YqF͋}�l��c 6&*f��_ҥ�Ɯ	`C ]������p]�Z�c0���ڋ��C:��D�+�^<5Y:s��r������f��PZ�|T����R:%�%|�q
���~�_ �ntl�*Wp��c�����>���Q,@����B�7�qL�!��l^A��,�c�U�m�~W@���F)9qݞ�u.x ���8JGPO	^IA���["�/'�|���$q��ciA�`���c��/���x���E&���ү���%L��_i� ���J�r�q>��u�K�!���ע9���:���>��zJ=�4mе���~���T[)�kvT��l&�_��=C�s&���J�*S4�) ����{F��b�m��9����a�����XW���˳�Q|���A$Y�uN� ��6��L��7�����0o��c(�ӄ�Nn:���v�EЩ���`�O2keь������{�?T�u����&4���[�P��{Jz���'%g�d��(��5�8;�Ẻ�%�5R<��do���Tg|�h�=Y�q2���э�l���(-��KA�)�xu��>�<"IU!���qA`'�'XOef�×E|��4�:����*(���~פi�Xp@p�R�3pO��HJA���j�o���	q�����b:�8�G�R@+u� X��S�U؊$��}n�)zv��-Bff'7&C^�oɞ5&�|��N�-���~���}��CKِ�\-MF�T�M�_Q#I����bs�u(-� ��U��I�J�{���{��Yݯ����$gVh)K��4DB�w.'m v���b�aigOo�g:R�����i��������2�A��������;��s�Ga���ݣ��Ƹ��$�<�_p��ã����՗)�\e��!���>̚Z�v�goA�?b
ۮٽU �u�'َ�P����=�W����gwz�����"Y��0=(��%V����W5H�hA���e�ȧ��t�?'��w����ec0��a�JBH��N<{�����5)���[��Ӏ~��m�*>6��	��s�R�f�6]��B,c�`��k�Xɷ��&��������LF�C��c�@R���V�EPgT�$�7(а/�G^�N
���ž-<�SV�ǅ��Q��U]�$���� Z��ب�?m��`���m�8ȼby�c�	�!��/Y����؉51���g�2ɫ�l�;%{y� ����3o� Ns�箸�_�鸞ۻ}�z�4�-,�tn0�]%�Z���{����{�HO��3HT
u�bL(aqL3�z;��T�"?:J�+"ui���'�������\�S��B����7��4�0��;A�2#�9��li��x���fI��.c���I�
�۟���Ϣ�:M oMsFc��Kbޞ�f�ćXv%Ү��E��
"z�v�r��	1$ր�C��/@��
��䁓[ؾx��k�	e:���z�s|�N�ɶ�C�`�c�/��kH!����Vfg��F�p������ylL�+�)F8~��������)�Ĥ���n讵�Uq�,��'�U�$�wP$�$�b�b����D��O���w��ן@JPm�>�Ȅ�",!�i��H-۲�ڢ��f���F��E{�?=,�w��i�o �<��tB���)��k��pp3�J:@�%�<R*����(ܺM�w�����B����i��O��L�B�u�2��^$p�K5h�ș��.�T��>Kc�}m�ӗ?����+ٜ����1Dp�����LV�g��t�"W喇ŧF���+q�XQL�΁��,�,�j��7a�C,�v�;P%b��w:����(�w���	�������ps��
?�r1��]��r�0�+I7�aq��#j�R�˶��S��p|RP\NyYJY렞9�o�4�Q�	Eڎ�0G(qT��r&M��	 TQl��I�fՔ�\�{g�����5L�� ]
�v��T��5K���H���{^ۺ[��
�)��Q��g�"b����Qn%֤>m~�6u��jW�"�)Fכ��K#�v��r�F�̟p�Z�"RB��L�w�:�].V{�3�K�(�!<� �my|�'����g=V�߅3�]�[e���^�FRCu���qc�J��?�V4~�xrdP�%���׽L""g)�.{�=�|�S�p���!Q�>�qC)Ik�K���R@1n�z�k����fuc��i��yS��P���)Yg�Z�H���ّl�Rs���jMwv�=)�V[�2��Y�<�!�G`v��2�R{g�[��ĵ�	��M3/�V/�i�{�]E��(j*"�sb�l��*.4֘$��_X��w_8���� 
�	���J�����w��j't��- ޜN��M��.�^��Iʴ�j��ۧf�=|���sݙE�q���B|�
���hLUVP�1�V�I�ǜ�,S	|���Tu��/�æ���&0%�}r�R���G���9��i����S�޷!#�3�Gv����ז��kv�s:a�+�AZ�X8���[t��(n"u�e��4kTgR�8��>xa�m8�P�$���X�F��W<����.���D/]�H��rķx*�bøX����)q��P�&����~�ae��MF�!*S~�u���k�(������;�#��4��.ęJC��WS=O�򢘒�XW�W���e`K���Y�e�w?
���`��R������笲�%��U�r�'����P�I��#F�����~���������G-�̛���5ިi�@��t�3{W��
��M�.�dd4���A�4�G3�Q~�~10(�Tb�v\�)��������6t_��D�T�+�C���6�PD�?:�ɂ=�t�V�#��x�cT�"@ͼTѥ���bJ�@��l�1��N������6Fh-�I"�m����Ol�2�iR�HT���b� ��\I&h<��Z������)�Z�Hnm��Xfjn�r��!�.��ּI4��_!8W	�qn,����3�W���q��1琉�4P��n���Y���)K��h{Џ&�d�t��9�rG�[����#�K`'�]���%;KLw��H;�����air�+��LnР�٠5E�<�����{l]i��Kma�P�HT���eW u М>M����:}�cHP�qǛ[΢�������4�{�DB���`w�,��U�,MUp�V���Aj�ꅈ��Z��(26���2�4�o����֟���0�k�ҕո�0c��KbY�6|�21�wA�NMo^B'$���b��M9ƕ�c�+�d�j��~��a�[�EM휌��c���bKg+��ߘ���T��r��",6���ƞ���G��Nن�k�6f& �y�۹��]݉l+k� ������/ݵ�'�L_k�g��ن�?�}GK���}ee#����4�˴�����jFa���FcCJ�0�����̛��L�Gn/���4��5���l�h�����d��{T�yT����%���ɵ��,Eտ��8|�X��9_�d\,xY�%�P�O�Ҷ�{�r����c\�j����ZEy�ff=Ea� /����2�7�5�;�h�k��i�;P��R���6	�0Z�9y2�J�T��(��W+2�`��Zp�����^a�+�+/��;�E��t�b�������i>6������i��[�d�C�&0�/�	�g!��ǩ�)�|��`�	̝֣ż ?�ٞ����~��0�4���>�O:Mu;��i�P���<Xe?�{8����~�R�
��>�_P�=]��c��Yk��J�.�����!����8:p�t�ۏ����!�P0}^fC�eYI�x����UA��#���Q�������~H�>�	Tm�d�i7�P�ق׏E`��n=;��%�s�N
V��ҙ�ǵP@_�[O����~X�LJ�aD���i�z��U�:�떑^�J����Y)�(��
��1����>��Y?���~�Ѐ�H����c�?��3:������z$���ʜ��#�Z��6.F�+��y��0�:�X�K�b!%j�TM5oGͯ����ޜ1�+m���9b�[�5&z���$��hް�F�%��%���l(�H`u=n��q��� ���W���B�=��)�a �*���M�)u���āӫ�x�26�`Z7¸�:�I����w�dU<�Cs�+��Y�>�%��ܔ(H)�Ӻ�����F��8w�3J�)�PVݫ1^�-|t�+����ˏ1��Vz��pL��2�5�&寱�{o�����r&���=�b� �����xV��IA|!�v"D\X��>�S	�mb�?�]�̩I���]��n!�g/��q��*�'����7J�%��;1�V�P�-��^�!�7]�P=��_M���h��֨�m�<-g��h{O��Z�ߥ��V�4|�L�L���<���T1�}��ںϊ�t+T�\%�(�01�{�k�{VJ'�3����|&�� �e���*	T�_ߟx5v���;?��*K��{Ugep3���<)/sqKV��">�D�>1&�d+���o�$!�Pf��t,0�d�a�����!��O{a�q��*E����ɃSi@?Z~-�,�~ό�i�$�{¬"��UC;��T��sώZ�^��L6w(�6g)�N��[��e�ۤ����Z~�*x��~[bk}���`k��B��-�71+���q��U�䐓D�3��h���9wr���
X��-��a7W�:)�4Kk��V�@�Q@�)�~���J����:���n��J���e)՟kH����_�;I�%�ڱ��_���du�)�9�i8���.T~.4��}s���lK=h�$�I��ҟ�L�eK����SM�O7#��H��JKo^)�6U�� �y�ۇ��_�%�<�V�cr"j�Ա t�E�b���$뙨ߖ��phS{�r1~{0�4��)�
Fϐ1q��
U���p������)Ȫp5h�����9$��F�{��t�����d�9A��c#+R?0��1RO����z.��@P�'7�ǙA� ���<'��<�X[�/k�Mn4��}W�q�	/���<�I5��Y|ɾV�e�1���m ��=�P�q�ǋv�q^��g��o��}�.=���2�ԫ��4?|�Hཱུ�1G���G�����~5�
�sb�a�y�/�#:�j6�^$.����<;_�C������u�Ԙ�D�9���2�f���IK�g%.i�C��V)9��;����o��=�7�Z���%���?JZ��L>iM�|����ݶ"*�찏�{�ʒ�c���H:O0)�!����A�	�����S]�Eyxd�C��� û��l�fb/���	�y>����M����4v�r��\o������[lg�(�4�.�t�\�zD�<������Z�v�e��<߰Э�줮�s8�P ��i~���; n�.O/�?�[�Y�8��\�Z����E����E���z]��o���JL�ܐkzuڇ���ɰM�6�����|zS�OW�Y�i�Nw;�^�-���q;W�p�x�QZ��n6��Iq�j���#�;z �D�N&>�_NR��Ƚ�6�j�)�WM�� �4%29����H ;k�l�`l[u+]Lc�__���5B�	p�Z�mZ��Dj���G�lV
@�G�"���0$[^v!�0�r5���ܓ
5�I��u_:��XrE�
tG̅z/�N	�97�ѧ-
vkL���nPgc:���k'�s����X�$F�˦1�R a[D��[�� n�}��ͩ����a|�B�N%�!~"T�0gZM-�!_i�Ǜ�Vi�W����<�Z�U�S� ݵT`�,���$sR��eP=wK�kZ����|�!\0�Єſ݋�'���%oXg�b3j�zhޜ5SV0�Ɩ�
U/[���Z?v�����������砬�U9�b��S�m�J�M��N頙���qxs�y}�����*�d"��P��cj5�;��'�.����@��H4���E�� (�aN�n��k	4��sq�Fc�܃-T�J����6p��:q ��@���m�2�Zc|Z��z�[���^����g��F$�,4s���G�,q%,ԛj�cpzK|�JaS��<��A�B7}��0�5�HG�R���5�eq��Bq7��E���Q"|�Z�����"��O`di�kI�s���.��҂
X����R}p�R�ڸ�j�6H���@\���YC����NN�C��
Iw���?T�=ļ�4�FQc~]-I�0�=�K̴I�*hō-S��:���kp"�m�4�]��w�[��b�e'=UK���/
X��A���CX�����撢��3]4ă��Ya��Ik�8k}�a�&}e�q�%��:��V���.���l���A�
/�Ւ[�����.�:�R�0�d�v��M�m�H"�I1��7,�^+���4ʽƣ��?����W\�,��A���6����1t����s�$Ýi),o�6'�  lm�sB%͟l'�`���5S��c��S��4���Y5���O%�<H�aֳ��k�����7�������r=hP�
�U�"�'�
���o���ҽt����}Yc���#z�E�6���G-b?t��HPD��E�[�!0�:1����<k�ő�&�1�t��q�nW�������k�YT z%)�!�@��~�2-�*B�za��d��nl�~��9bV1(�������������G8��#�o��d��X���&�Z�PF(�W$����@b�i���P�,��)g�::Qd֚��k8P�/v����I���O�*"v�����4�ε��O5�����hd��o��N�r�۷��J(i�,�}6���:).��\�W�?L�H��bSQK�
+�˲�g�M�1Mc̬�����Mٍ"���0ez^C�l��k�S��XV�h"^���������s�E����{�>�	��Ӂ�	�����NȨ_�WXA�%��ni2{t��-���Xw�����_�܁Wz0w�Wa���o�n�gN�Wm%�?<B��}*���y���j ]�]��#.�B��Q��=x��
ֈK󷛵<��X�Âa{b���zseK �gE0DB���-S�2Beֱ#� �;�WJ�T}�ģ-O�o��)Du����qKZ(�}���� a�$m��s��%�?��z�*x@���n������0�v�Pr���0��YV�-f��vupo�x����K��/����6M�g+Y���[N3�F�MZ��������H�8���@Gn��Pd|���-���"���ٖ@���w2�i�������'���y���F�D=��r�8n<�L�f=>PY�{2rL��%�8_�Z�N����ce�~آe�/ť{�O�118B�}2>F���
ΰ�1�bV֯;u��a�a~؛������h����n!$����?y/ �
��`z�A����Pp�jXw���-����F�
�P����8}�$r����������Y��;m���$���1�jAj����zQ���R��M�&i����nrr$H�cNK�>��������B����E-n�+��uW��+��"���e{�l�W_��Q�y2�����\l�>� ���2�GZ|��f�9�}� [ ���{ʤ%����@1�i��z���� &5�D� ���E��0;���T�C�}҂�U�Ae!U�z੉fY'梠�uU��g�;�1�~��[��<��i�B�J�l����������$�E���zʩh7���W�K�(�3*��	�Mpr`0�Z���6l����6�Q���,�0�yRe3�Zm1
S�� ��K��C�M����1"�����ߕ�&�v�E)��3+'����(^�W,����x��<�-eg� 'E{�������%È�|�0����(����8 =`��b��j��<V0i��D�&W`��d�|�p�����Qg0D�{�X{�"���r�n	5N?}�,��ʦ-9���BDV�o�}s�zN1^!�����}�q���>F57��������WӒv�v��B�� �b����<3]�ᅯ��9���X-��@w���N��]��z���^5#�W� k �TT��w�)��{����@�e�u�A��H�j��^�X����A}��ʣ0b�ȧ�APO�mLnq�@�3�@�w���=�E��t��t߉e�����X�)��>$�'Rp�Ll'_�0z�p1Cx #����I_�������vq3�M:��oe�pt��K8G}ei4���P���p∵�h\����)֏��y��UI&���j��Ŕ:�ʉ��OW�x��hD��׈�Oc3�-�K��2�V3{�_���q���w�>Mɫ	�I��Ѡ@�����8��`ʋ��~z���#��ƻg��Xo�g���D�L�Z���`����6�ս��b�/h�r��Ř�d�ݔp" a���icq+�!����Gt�Ӛ�E1��%�`��.��4�wsP�?�/E�'�CYtc0��3h��"�}K<q5��|���gYc���֥-F�Le  NM%�z��PZ�tr�S(tn/ f81��f�F��j{ǶD��W��O-Oω�!G�%n��!�Ġo�pgh������-�q�A>�A���z���rFV ��7�*�T�{Sm<�Mb���;	�{�����v	�ut7O�Ƣ�3?���>���P�a��� �l<B�ƁU	�W�D��z��z9��2�a��!�\�I	��	u�|4ӎ�O�R�3b�1K;f�Ĩ���ww.�	���y��Ay�Pt15z��ܔڴ��K�uxh���.�cB��r͒��o��z!�ց�S���;����O��4`��L ���f����Se���7��
�Y8��LK'R�DpN ���xz�Y�V��L��DD�곴�����3��Ȉ�@�Ȏ�YMj��496L�7:���y�M�|k�i���j��]�	!�޻n5�/8�ŗ�������jn���������C`�4��U����A:5v|h
~��,?�3x�|o�S郂�#�g����������%�޴V����V,�b�V{�|Z����A�dZD�ayۻ�N���	��|��t�Xo����^H���g��S���)�P�d���f��,����A�2�g[=w���
&�)N��_ʬ�ݓ��f�-���g���YV��S������;YT��x�г/L�L�VR�ǂh�!2�Ú���*����2P�L-��F%�
8��� �������2�K�F?�05f�{l����Ò���UKn'��^m(��$i?�5�AU��k:z�Q�Lhg�el���N�ny�ڄ�[���� ~��%�|2��_��p<���c��.�c�I#��V�B�o��o7�������Yz4<���3,�*���t��Fž�/Z��T�hB�5��<-oU�\�Jβ����ߝ@n�z~�ȊV�H30B��Ҳ��14m`k�vl��X㥤Y�N�Q�,��և��Q��Z*I�+ED�K�F��3�P��p��d^�²U���?P���)��r�ix�<4];������Ȧ:�uG��.�$^t~�.��9v�ա��T��	~��,�쌞l��/aP�隶�h2��#$��0,c�%^�-���l�t���� �g�T���*��J���%�ę
���RO������ȮX��v��{��;T������z(f��Rs�G��負I!��~��=��n@?�%p������϶������p�k<2�?S�1k�j�����0lR+�0;Uka��|	�m��E�A�i�<Wa�A��i9��S����꒼#�^}n�>��Cb�~��:L�9�u�c՘�0�V�7/�n�D[�U��A�m��r@pO��,`NY=���-��*�@j�Q����t�R����e��f9��O��4��+�J=��C#̲Sm����5�����C�>ZԞ�c*��@��=;�2���z���{����W!�< l�h��Ⱦ �Z��RC�Meڇ��:�u59�Uޅ��ڦ�Wk��"AkaTjH�n����];�4�ʊoG��q���D��?�Ko�@��V�l��?�z��?�74V�߯"�3~�X������?�$��d���d�1`�U6��԰��A���lm,�Q3j���6�Lp�K���QbwRǗ8'�=�~�ښ�0�?�9��d�z6��?��k���a����h|��)o��d̜��T9M�;8ٗ��-�MoЮ��˧Q�����3a���[�Ħ͹�G��\����I<���bksz֊�(�~c�2�Q�*>��m
�n�,��|e~��e�.���)`�L�� $)z�Cޑ&	���os)0s\Ca$�Z�&��h��e���F��3]�FZ8n�sS�=�*�Z���� �n��{ᵭ&�3Ŏw]U�#mW]G_uV����`'8�E���l�ǈtS�m1ړ���eZA@A����ŎXu�ӣi�Of��7�R��Y4�Ս�m�F<9�$L�F
E�}�D���_ ����t{o[�I�4��C��ȡ�qÎr哑�!��\�nG%g!Ur�����T�9Ǣ��v��s-���Қ�ŭ�R���L����iNc�[�=�R!f���S�7�?y	!�w�ժF��4��|�^��EOU�|�b�%��%b���4�xZ�:d��tK|l"�f��<�H�f2H�$�Θ��We D7ϴ��k!�,���"�i�"�z:Ð	��8w~o�n+~j~m������˄�4-�r�N��̱��^�!�����^�t��P�Q��\�~$@}3�}tPy��K�a�AmDC�Ǯ
o����x��Ys�Y�sfڨ�9m旯��ۛ���P�+�r�2�a�:��)U.�oa��L����x2�o�7��glD���6똴�FR�5p��Ǟ�f����p$����&a��@���b�ng����Ui|��=� ��~��[2����G�;+�b�5�B)�	
a=
-!��rEԎ� ŋhX�������{vU�A%��s)����mZz}�dE�˚ވ�X>��-�C��t�������v u 6���*R�G ��}w�&BAo��;�zS:	W�`�j��Ұ�j��`3\����^P�8�7΁�lbh�#�@�o�䭎��j��� \�a.��x���0TB�)z��3��a7���xHZ�#^���qk��y`��&����7x6,��e󫮊�>ޠ-�h�J|�jY����0?�]O���OOL}���kO`��j�\ ����TX��-�LQݿ1̄�n�ԓ��� Q��*{�/�A�Lt0 �^f�#�����W�Ux��,��(�9���cMW	��1��x��e �!O���!��C�Zs ��l�>v`�)�'�
���$��f-	k^x����\~>j��[����09Or��3�tS��g��,J���'����f��$d��8pKd���O�*<I��Kucl�BH���!w�;3��}�ߔ�U_�y<�D%$c%f��[Ư�.fh�6���o��#���Z��X2���z����{�#�)��X�,�N]D;y�B���25lIgi��)�MI`Y��
�N�wX����������"�$��+=PE8o �w�
��Kw�v����fWc��H��҄ª$�jY��<�{�E!u����+���{Y$�,o���ǲW>���v� O��m��Dz,6��v���s�e�
6�������?I=v.�[[��-�L�?���kՀ，i�����J��7dr�X��ٍ`d�5rΧJ��ِ#(|��Ll��DP����`�?4��naũ�ۯp�ΒT1l`���o#��$����+����+mC�����e�8t����}��e щ���X�+k�	Ku^�/����h�z6:��	������}`��;��i@�lW3 ��Yi�t���	\l�.����II"�;ӖG�I��uE�<S3k��{�ciWIxU�e��&c�R �oq�?�"�K�)�\��dj��0���]���5Fx�������P� ��L���!<���3nuϱ�'N �_�H(@5��҄`N'�	��d9��*�N�K�n�����?ڙI;�V}�]D����-�Ri@��ě������������ĝ�S�B�ݶUyL��[����cIzd�L�ۢ�K%�+���lR�����!a'�
kx��x�U.���K�a�A�ׅ��#��<��������O��*��m���ty)Mc�_�g���H?#h�������uԈr$ܳ�kc1��p�W��
�f�3>�_���qE�����o]'�E#Ӽ����a��h�	��"$����tWVG��p}H��,1F1:�ٳe��x�I5]N	J��]n=�����ED��N5�#��8�����Ȥ��X��qt�1`h��ȡ��9/��6
�o��ui��+U1&ib�(W{B�CGe~��t���&7hk�~�S��%K@�`�:G��	�ba#V�;��7=��R��i��Jx�����$�p�"����N�TӪOKfŋ����NV�UK��8��/���ɤ7R2�Xԉ��VH�8����Vu�Rڑ5���'U��W�Z������Җ5y�jn�XQ��m�+�����o��mB�@��@]�06�-�:K����Y�t4G��`��n�e|�������nME�d]�z�$[�2�:_�z�ƙ�1��#��
>���fi�}��u@�G��θ؎�-�I����X�A��������+<�������Q�,�P1m�й�w���vkX���6��=�`�	������5c�NbTi_A���%��k<�kF�<<
���׷�-�\RNXw�/4ʆ=�Fŋ�aE��(s��FtCC�nD`M�y<u升O����-��b����y>��Qڳ�uL��)�l�N��`n��w܃���PP�vB�3�j�m����>���<"X�B|����1�h?K����O�M����m��wB>�l�.%�Eg/�|���_��Vs;]>�>Q���=��c¸z�wv�t�ʹ�w��͉.D����΋z���<��b>������+���k��,8Შ	|nY�Ke��Ke��ȘX��FO"�8!QͅH�ʥI��tJ�%��2z4#}V�^$�-m�1�-�w����^���9FH�OO� ��W���j6���M@���l��z�z/a�<���Z�޶<�:�L��M�A�%�����贔,��RAЇ�ku�����՚ܑEm�p#�O����X%����s�҂<֎+%ң�^����?�����V�u��,i�>q���RF_�<1�Ј܃a\�>�ʧԅ�N�H�ܷ;Xpѻ��a�$�{�@�xJW���Ͼ�E�3��6�L��Φ����u�P�M|`�=��#8\KQ�S�P#��U��C)�ՊXLf#��.���$j��*;���x���L1�L�g��Q�|b�"��L��1v���+y$9c�)
p���9Q�h����=��P��Xy�!wI���ץ���� D�*t�?��֘�h����o�X/��r�p{�H�mJx{�l'�Ǧ�|�?�����e���oD�\e37X�f_��?f���i������{�Cw�h&������)�;�S��5�S���6�!�M���Q�����v���g�(�U��&չ
e���9��
L(�ס�?��â������q��X�w���,F��q�����l�G˕�~b�K��h�:���i�83̠!b"�����	��e�� W���,������^ݙR�ㅡ*H:��2r�kMA�����붦T��0dS�=)N�r��i�
D�M�����X���&�f2l���#�ؿ��z�j�͜ǩ��7���K)��&�*C�QizcV�K9��q�Z��>ٌ\J[h416;\�����r�#�9�}��ᚌ[:�(��ݯy9I�*c_�o|`5,��4q�B��,@Ͳ�:����H�{���߶���A�àK'�z+5l��9$��lI"@�j�e��� �?���g��Fٳ�:6N҄XY�"�K�B��3f�/�'�Qģ�*�B���
�����Sm�خ�ƛ.��R�(�p8<�N21���1˘Fnlhm�^���|��{c ������p���|�b�ANye�:��%�'�����@����%u���a��=��}ؗ<�`w*N���5����a:�}��C�7���w�
�ʩ�y���Ēc�b|܇o�UQ�w�m��=d|��S'jݮ5q�~�I�ń�m�B�ѻ-"���s�\^�d¿|Le�Zİ�J`�VP�=%*$F�'�b�T�ᬺ iG�n���$��~9��[�����(H�{+,�	dwvy2��J釛Q6N���7J.��C� Ѷ�բ5>ܠ�-�Pei2�z�_�\X%oթ�񃆡���e	�4Ӊ� T�Ǆ�tƛ��8_C�C-t����iC*oO���\�ֽ��Tr)�b)�����l1�ĝP�^�ҍ��,�"�5�5���.Z���}^r��]q:_`w��=�<����U�3KXL���2����J�u��T��N���ը��c�"ݒ�_'��70�i���n��I$74���G�(��zL!�d /.tq��%f�|(�4_ӄ��6�/�%<8T��|e�j۬{T��Ț�a%.)�<��� ;�0�ٟ?u��k��d���H���������>�D��W[�b13:��u�o�<	�A"p��ď�(G�+(z�m�_u��I��J�������)�^JFnlL޶��kq�b%Ι��nH��e?)��(RC�6]Qp�p_�,��k���=�MiŽ1P�IEeW�����}�H����?�jvH�pa��8����"�]Q7o!���D��r|Ua�;���yrm�nr��竇����iF#e#6xP��΃t]]��[��yM�.�������H�����|~�F]z򧔋T�|�e}36h����b���Ē@ֿ�|0[�[�f���*Ǹ�AQ���$�}���Zl��I�k�MwXk޿S޵�z�����_n��6��
C�剑�{y_E�j��L����VT�YO�0�GR�D�HM�OI+�����K֔������>cV�`�6Ъ)ʽ��?XiV9�1҃�<���}���i��R��*҃�8Gm d�%�U��b�[{�MR�	ɋ�p�#C�DzG$���\���z��s�s!��I,���:�FiT��(k=����D��Q�]�w����[�|!�{����K�˘^�����!3o��lղ����]b8�>��'��rzY����_ �.U�F/������-W���^��aKZ����j�Q�]L
kx_�.�@F+}k��v���H+Ih�;�0����FZ����E�8ۆVg���iוJD��uG �p�8R��X16m�Ѷ��;zbݸZ�b�`��b��F�8
��!\��{<n	�0��2�bU���5O-M���_�`�.r��d��K2|~�����>�h�-^+�%Ċ0B�}��� �(��'�L�+�mRf��"�W�v��O�M�d ���͗Oc�>9����	�t���{[�K�9�}� ��݇t��$�F���`v퉇���<#m�~��Da]���������;��x5ZjU��U|#D'~JX"�RL��ˆ��+3���_&-����l�@J'l01X��~a[�}���3�#�>�=wʾ*�1�)=�mu���a*GX����]�>;��/��O��IU
�
{r��(��4:A�w��nF~fb�R������8�Sy���b�`߫���e�CI�Oy�g\� ﾏ#oRM�^A\r��PX~YE;z�U���$&���hy�ɭ�わ/e��s�yFD��+D�!&���R��j,���}�p�<%Ý$|;�\m��w�^�x\h���U���c�;7�E
b=tN��PP2�xβ G"8-��?�g�1)�1,t�"�O��=t�}5�Q�/�G��V�X"5Q�'�1��ɭZ�5��V���[ħK!�:ta�q�����#��P6��<�����6$����n��>�:�\G�����7y��=�xI-���¬�'#0�Ƨ�
)"������W�x/Qdj	�1ĭ�˹�<�4��5�[�y"+��.��R��dV�Hn�̥��֟*'��!�6�8���a�0�'��+M�׸��(x`�1���`�ä�������˜��[�=���;��s.g��ٓ!�la�9M ��� ;P�%���9�����h��M����%j�e��I�*=Ľc\���,�t ����=-���>��!��}c%5�����<<�I�]��)�lBy�hO$��C��g���)�b���HZ�������V�MC�Ə��MC�wVcv�651iL�q��7��]�89�hAA��dC��� ���l*Cyw�Z�\��do,d���*���i�i�e���xp,�/SN��\Sph+:N4�=�*� 9�]�׆W�,�M8e>I��2W�n֛8d��6d�������MH�p,ꪏ8�:�	�4��|���4+�$A�HW�Ɛ���&���$X��9ׂf���v[���}t�L"���,��0�M�J�A\����h��N��̟W��Ď�1S��-���e3��E4Fј�9\�W�fK��tQ��5qW=C�!K�.C�sh�G�{$ZS���-�A�C�̱�9��s&�I�- �
� �P]H��;-�D\���?�f�)��Σ�W�'�IpI������c������u{�4�G�������6��r�@��#m׶ZZѳ���ғu�Ë��Dx��&�Q�Ŏg*���L�c��F�=�Qȷ��ML���3�����f��;���V�):N4�2�6|@��h�s������o�]:]J[�u�x��}��H�أ0�� aW"��n��.��n���X|�� �(*���%w"�V�a[�&�_$Ċ�f�7��a�%�v���c2%m�a{���z�r���� ������n�lZ#�`��Qw���jݩa!d���y�S&���\�!����b89W�����	R�x���.�u� �	�V��I�8���2�ր�AC^$L�~sL^L�����ɉ��d?�.ܞ<�P�ۘ�K��q�q���"������O�H����ZS�!^�����%����2���O��NZ��A�ۺ0B�v౉��uv�pѷ[�/���<~�qˈ�Ol����p�2����!pb�{K*��d�f�St}��a�-���@�f7�+�F�&�7:g.�k���b-�d��E0
����1�I�׻5�^� ���a�m�ogY�?}�%4�uY�/)Ω*ݣ��n)�.'"�~����e'r`Ɉx0�W&�&VL�zO�Q'.Ŵ���A�Z콋a Ŵ�2��a���x��Ηw��	g���TV�N�:QD�eg ��O�$��0R�SW�Oޜ���G���%y};Ew8M�7]Er�<���U!s��S�����#C��⸺�[W�4�Va�LGB�q��s2�}8��'���1���sS�R>.�O�!I$��0��,��V%�z�D�z�c?!>�ľ~��q{��'�~fEw�J���>ݹ�덏�i����Z���35;����&m]���;��򭴧RH��Y���)ތӔn��V�3
g'�m�|��I��e>�ڗ!#�k|t� ��,�)�6
*
�h9;vh�K�wd,�o�=Qg��ؚ���BN�Sr�,���.��Z'8JI���ق�,�
�
��L��c6���K���ܶ���]������#�D[=8/4���5��[^�"�;�6�ן��ئ�M� q_�F�(G�R1]�cj��!��ź��mI*(OCz\k�����@�_g?Jq>�4$D؝g��Y�b��f�`���^&��a\�Q]�d�
m�ƙJz�H���c!;�=H!rcf]	sV3�W��p��@T}m��g�U٪�9�V-���{�F\�͒���s�$�������7*��b5�.^�b�Қ������"9fe�˕���#8��MW�M��aj,z�H,g�[�@��%��Z,�%g��A�[s2P�S,�~	�0��t��S����}fV��l�p1dRW3~�3���^J���=��-��!�l2J�F�t��z�Z��W:b�u}�1n�3szw��G��5r?�+��c���N�ՠڦ�	�HA��sQ��
)G{�?F��0��K�N�) Q��9��I�~��n��N�潖���V�z�Q_ރ�w?v����]�ֺq5EaK1��gs���`�r� �ߪ�:��IF.�������b�\��Ȗ�ؽ5/���Ff��Jѳ��g��&
}�r��m�9jU���<��'��SQѳ��� ���l<�c�:�j���&�(Qҁ����z��9
��'���]��N���C��I^$Q� �W�d(N��	CSK&@�ϥ�n?%���靮U3��W*��վ���Ӯrr��9�7�o��KQy��Q�����mA������vj)�8��l'+��:-&����|XQp8�f��)&}��4\9��A��ɮ��۾w�	��[X��]ѹ�x���j�������X��@xhLy�t������	�ի���e�x|(�OP�|^Ǻ:���a�HEq�������!!�ߣQ���[�Q �� ,�zO�T�e�Yx/�)��ߘ\%@��T�3~0@n"��o[Nھ�͍�F ���ӛ��7��1J�AY���%������/<���h_��#�9�< :�J§|�b�it�p@`=�χs��׹��?�.����I�d>C%�,j��g�m��Ȉ 
��I���t����<R>�O�%R�����6��0߯<փc������º��ѭ��"oob��q���;���#Ң |k����tV�����=��EGmwpr"�Ȁ;1kh�
�B]�,Ԣ��}�����}2?��`���L%�*3}��9���Ӝ�p[�B�+,"2yحeD��65���G@/'��+��]�~�4��X%Ц�h�UUNes'��<���>�'����t����2����"a';�����䇺�ʀ�ܠkD��!�z�e[P�s��Ӎ
�����������q)5��A�������h�K��� �X��Sx1O[(��r*^�zD�eg4M���.������x��ƹ��H�fj"4�h�Q��|ʯ���nݛIF�v�,0ž3\�R����w�#h�������T�{�&�m�t
�/��L-xv�{J��`�kBŎ��JJF��q�P�^z�([��(vKDNdm|�4�������:-͠���V���߿�	�^�^��?נ��u;#N0�O��ټu]�u�,�pM����ŵ��İ��Fk�E=c��[_u����-	��G�����#�"5��{(y@��T�������{d�Q�����v3�/W`� �}WЋ��\��[j.����*/�b�ZV���󁙒*M���kWQ�e_@4�)�����+=�4���^��( �{�/Vi��z�aӒ	� @�T��H�`���K�R��+;�շ���a���\ϗ֞b�W%�c�2��zDG��������k�}x�����П����u���������;��{��P^c�]{� ٪÷���At!C�7n�t��;�6IS��x�j5�P�C��Gd�����ZX�w�S�8�n3Þ��#/4�g�� &�mWA��A+�OJ#��QS*R u�j/媆[`���P�tU�x-a��u�ar�j�J'����mv�s�Q�鳞9�h��r�!|,��U�����0o�8��+�WD�/��ϱ�ڧ�d�����-����l����c��7~M���V�� [�� �	�,���<���B��J�=	��f�n�*���p�;ڇx��6�&���}N�`�g�� ;�s�o�vO���>����s�R{؎3�@t;��:�	�bR}���ƒ0���x���t���|X�� �0�萩n�0��v)e�� )Y����H�aY�.�K����Zx"�f��Bإ�}�11E�<./,� J��~��n��O���Z�6����N+wٸ��\����K��V�B�Q�m�����Ё�֟�&��W9[k�ڻ��M��	�Ȣmn�����O|b���K���J6v6�_��K�>�cCG������V�Z����ؠ�L�P+)��K���-�-��A$�N�k#�׋��&Ei��;F"�ɬ�Uk(k\YD��s�b�R��T}H>��'@xR�5����������u��<޳l$���{a��$����5_�'Q� ��9����J1�j�Y��c??6lO)��+*͌	��*
#�9��)��{D�rvMX�ƙ�]	Q;�L��菝g�Z�+�GF0{�OE�P��\u�Ee�[-}�m����}���]U����nQWy�}��f̊ l�I���3'�f��T��oX3��8����Cȩw�5+���M'U�V�OU~#1R&e��Z����s�[�88$���x#� �D`�M��ev���k��IvG9���1�����%��Ė�1
��q��E��U��P�[9(q7��o�.����įA��򂆦�5�jL{��)��<&:(��*-��>h�]	�s�nMZy�Ȕ��2-"UM%l��K���pՅz�vS��Y2'C�ʼ�j���s��3��Hz'��;b�C�%���e<Ӏ[z���yP܍
�.�,�xQ�
�Kw��,G2�x�f���c�5��~u5�?R
�Gr��Ɖ��d@�g(X��u�t�t	B��L��^�Va�+i��\� �E��
  cѠ(���@����v����Q|U�⚽���N
��s�����d�����'�z\�z��J-4��6I@"�M�K�������%c��91\z6U��4v�*S�Ȯ�&����%��E��ԏ	�KJ�������0J�KG��6��!Z��&ӄ"��pO(�%��6:�Wٸd-�"\��R�.o���(�ty���F*j���o(�������}�9�����S9W��Q��!t��>({4=.�Lv-����X .О�w:�Q~�󫡇s���cs�	��6��nLA��T��㨤��)�!�z5 ��N�)�Bx]���`1
[g#��I��L���+����.S��;�3q��|b1>T�ɴ��`2��UX����?����a$e�% Sy@_2����I�����9N�2��-��s��a^q53{$�{ZC΄�}T����f�w0�$a�LV'}׾r�*�r��l�z�$X=� �C�1�`-�4CX��ŒP/�hm)���&�m�!�J�?�Bh��N� :6a��"Z�L1��,?/�Z ;��!"���H���ҬJ�f��P�{ދf}� ��`2�o&�r���,"f�:<^[�{���j�@6.9�,I��3s|pk�W�x~�^�/#V;���j2�K���?s��\S���fA	)nn���L�` 0�c	G�� �(��4L=gd#�=��F����3'B����i{i�b(�'�o�?�^��@?ծ=u�Z�xET\������(����?��Q,�	�ӏ�?�Aj�!��4)��|E���N��?��҈�GMq����W��5K����w+h�� ���z ��F9��߈�V��d���zaL�lj�j��ub���B�X�w���v�;\�����W'�P���J�$B3�.�q�zjL#�g��)�B�j���J+^⦣9���y1JeF#w*JN^
�aF�~��WY��(�`h3�H��E�5�̝OMb�v+�h;�V֫�� �0Ͷsކ�)����/�#�zI��-�Q���|>��g�ڂz48�f��;�\F���K,��?H~f�+�b>C�*Hm��4���3�N�M5���� ���^R|�P�;O}�����ؙ(}O�|���n���\�\a�M1.���p[�݈៻m-\�YE��gEt˔�XG�v�x�f�ӳ�ۯ�NR>}9�g�Sv-�!T��p�Yr����,e�A�,�G����� e����W��!���r
����[�
��+#Z����ںz��F��d���CH�[ܯ�Dʯ+�~����N��p�V#M��W��K���[���x�₞*�m�Оd����|P�pV��<��|Z�C�|H�\�J��������;�V%�)J� ��nA�ӽX����[ͽ1fɱ��;{�dE���yY1���gX�~����u�#�������zo݀��R2z�WhM)Eq
�6����F.��@�:�	"93V��K�}��:�ݯ8Y����C- !�As��m�����oeW!�c�.|q!�cUJ2�Űu�Η����~��4�>.���� O��xUq�de ��'�8� _1P��F����:�<rҝ0�&wS���?S�_�7+0��.[�b����P1oY9��@��&y#0��cjtz+��K�HF�̞Ȟ7���7��<6h�����~�.v����P	�'H�^�A��H/���Ca��uX����K�����䌰[ݹ�j~Q�FSk4_��Ņ>ë�ew�|����i�9t)�g��u��w�-��^��YP��j�,o�nK��az`� ��(o��l}ND��R��D_!���	>��
�|5gLEr]����.�t�A��X�ѯ>aO"ӊ=3�ʎ�N��g.�0�u��ҝ���ʑ8E�Q;����s����UN�\���u��q���̘����`��LӢ�KT\@ǶQ�ckg|��՚����a#��	7��]r�"P8CS<����%ڬ�&#YF�:� �C�+J�s�CV��POf	U�Q{H܈S͙�
r��EO���?��gQ�
z I�|��#�ǼU��N�v���2��v���_�!l]XQp�M���[����s�t���#��qx�	O򃳊�ݤ�-nd�l�,'	�/��^�'������*�P���o a��Rۊ��V�8������^��E���\�Jl|S��a�kܯ�n{�	*4�n��)a��GM�n��|q�N����F><K ���˹p��{�J?���\������A�Gs��o��"�� �����h	B=PI��5A�$@� e���������K7�����ٝC3a1
�1(��B�^�����,Z�\n��X���'��R0w2��|�Q�l"Qj�Zk�bj��ַ	�V���M�g{�
�Yk��ԣ���$�Z��|C�ɽ��|.(6��Y�Y�]�q$��J���'�������Q�,���{�%���l'4̓ZG<�;F��&���>�4���@	�|�?�.��	8ц=��>m����4���I��Ba�ۚ:PՔڑ��ʫ��9���`P=����2&ŊF�����6�YgY����Ԍ���\�,��"�` ���.���mq5mLPq}3x&^;$��*���hl
�����������t�)X���K2�:�Q�Ä�M��0�-��z�(���E� }�ز�n���挗��Ȫ��kP�O��eam��� �m~����Ʀ��?25�e�*��.)��)xs����\ے��Ҁ��!��|6җú3� ��H��Å�˅;��;�#��]�6����e|C��k����DՃ� Ѧ"��I�ž�nN���4��g��rE�e�ז�
Ґ��,�:s<� �cdL��ݾ���ףo�`,�,�� �G���>�{ _1Y2���#��F�P�iu�O@;cz?y�2
�Tؿ¯�D�5��P��+�jM}�?~���u=�|&S�}��t�$��^n��V�3�Z.���T�^a��/�L�uȃu��cbʯ�yI���*�S��J$k^����P�8����d��-ZG1tVLMPC�.R<$��B֫G �(9s�Ɖ|�#Q<Z:�f�r�#�!�%>v�0���M\����d.�P24g�ύ��)~G1VF���� � �~<ײ�R�&KF�������m#,���4h���1v.���-��~N��O���>'X���Ԥ/��O�:��4;C���;�����٘����Jṱ�N�'��T�J�f�D'�����N�#9ݞ��8��õ-5���ѧÃk���㙐���pWֺxg`/��!A���ݬ]��Jlӭӄ�.��Kg���z>y�MH�1�جƸ���|g�cS	JZ�.�h�SǪ*���9ē��D�2����VY��p�l��K�iW	"'U$snm:g�'	����s�0B�OEB[.ɻ&nT�šF����Pq�s/y�T�O�-y}z�5nw����떽G�$n2�qިX��~���W��ọ
�G<c�~]^yD|f_Wv�c��c��o)�bo3^�?���SV/�z��0Q�^��a#Ӳ0U/s�3V u ����M��X�g=M�"(� rŧƑݣy���9Pv�����v`[��il�i��;��+���5O]@�pw��y��;�c�������x������9[��"�����N`g�8 �]��e�A�V!���z*ս� &ZwDk�ajV���*i�4��A՜%pn�ϩUk9�8z��{�����Z��}�ɮ����l�*�>�h����+�����V��9ђ\�~oW��u]S'�8=��@�LII�Ĩ��� $��5Q/o{��e���$�#��7�[�,�d�.��]�v���]_P��t���O���B �J2��XB�7�ʍ��<�2�:�{az"�0��7n|O�����3�V7�\���$Ժ�=h��/t��5|3oC�W����<d�e�_��O� �_.|�-��5��h���k@�R����(�������8��&̓q�q1�qR�,�q-�G�8��1�z�͜C�x��@��K;GFf{5��7X��[�{.`E�����;s�x�`��9�d��7Y.�x|��w�\���0�,�j�ՌᏅh��� ����E�� <�G�?��y+	c ��|��A�j�Z�D�H����)�Tc�WY_/G��_mp��W���I���SZ�YL��8� ��<�K|e��2M��kג�(:�"z����տ�p�[VCd<GpiۉI�]Eta����t�i���.�ZK�ls�s�����!�^5��G2�Ww��t��D�[����p����Lم�eF�9D�og�Ɉ�Y7mQ�:s����¨���]9U�WG�%<�3�)���>F �,M��k�wC��W�V6U��͏48e~���qƂ�?�6&Q�����[ϸ�4؀l�T��X�t�v�I�G �!-˨1�l� ��� U"I��²��3�ȿ����:R⎹�����7��WeB������Ts��A���	�Nnp�%������ek��4�:�Rk�<;))UF����?k�}�Z�kC`���ؒ#�{����G����v$�њ{��`��weP��p�o�=s -3E���Jڃ��B$��$N�W�܄����l��հr���h���kGG�U��R���-
�Ӎ���M�؃LՀ�ۯsTz������u��1�
s�G��z�$�E(�
��L�,�F�b6:�aD��:���P�JT�W���`�WP�s��.�r���k�0O#"��(�!|�=C�0#e=�RRI.�Tȵ�[���hh���Pf�ݬ\� �#�������k�rPc�����sX\��;��mե�x��2�/Q&�ܞ*�o�9�N��%�
L%�!�ωK��(d0@	J��-����Tr����$��o%˸6��$,�VT�	F��!ۇ2�=]��&o{��(��Y���d���|�;�u���ެC���.|��D�`Ӛxd{,?
�4����b�e.�V��D����g� ?m��;^���P)�KY�U�yƺ����~ �[�ozv��,լKq���\^ Kmo�;�a��̺��O���g�"����n�!���1j߻�K�l)A���v��x�S�/�:-����4Q=ϫk�֟������2@����޿US�Z�m�y���Og͐x�c���-�$�6� ~��
`|��U�^��+z!.���Wa�'������������zo��S��5N���@hm��0���M�H����R4�uܓ�@.M�`YĂ�H>
�����ʔ��ZM1|�t���V��M� �ԯe�fΤR�����Oq����T ~���B�ܞ��5�}�4� ���������Qs����$�4yXv�z�M��`��%�b5��i͒���m�Q�YYEP��pT9��$��Қ f0���~�]-��	�D-Y����!w��؛(����x�$	M�����)�*�߇gЄ�K�����|>;����T�	���NO�Ǖ^�t�XD�Iܚ�^>��(�q�J��:G��S��mn4J��Н0�K��E ���Et>�_��@~x���y�܊+Clg!����TX�������P54���ɡ�_}&Ɇ\��5P7~� �X_�܏~��S�D�m u"	�B�̔���t�|9ߣ�Oz� �B�!A$R��&(;�v,$��s��n(���,�]W��伓ʤb�[Ž�Ba��)�`�X鰢U%o񒆁!�j(��_h	��;��M7B�`^=�X�jL�Yغ��"���_�q<�n��x�"�������'^�䴴�� F��p���3N���^�M6,p�s;G.�>mC~!���D���h��ċ�h�8��۶K{�ְdf®q���p�ߊ�	�"%5ϡ�嶣�B;/eYL���qqF���jסc�$!��b�p�4�c�� O���B$L�f*"3(�m���6�B�&�������T:�>�S#K�hQo�')Ol�p�$z�W�!�>� �&=�f���
Je���
R .�N�\g�cO��T��O]�6�� }�(B�*Q�[��L���ֵ���<�a^�I0*k�,�b*�3^�R3��=���Y��z'���:�qeS�B7��s.Jf"[�=�xt/�{�8��{�@�bލ�:5;�6�7qgV&��EXe[e�~�9� ��~WʔM{Q��}���}C�5���(��,���Yc�p��t�8or�3}�P56�q�b���_�4��5r���9"�Q�8}�����b���?۟�y%[	���h1�2gXZ)�3���28�� �t������g,n5����WQI�R@/������Q�l(��z�Q,����~���I�hF��5
;���D��@��u�)q�X|P �P�r�V_{"�����ev1: лhA��4$��H�
C�K��L�&� �S��M�B�>�1����\�������7�~F{\�����"݉�1��y���n��"�[c�N����������Ƙ��vJ��(r�	��ɗ�$'T8?\��U
�Y�>��X�xqG�[��sB�ӳ||����Rk4���L�aЫ�p�D���'~Zop�Kn��Yb�ך�#'� ��1,D��4G��e�2��s��"@;A+.��~�vS��V5�̰U�"P��0W��]�i�<�2	��_�(t��\�S�U��^��6[�QH��}�}��l�Wj0��LW����R��n񵒍��'eh6�	��o�a����=@�˯�����V6)#_t���*�O���c�
�gl���q
���	F��|��V[֦�lO�����V�95�yuƶ������l�Z�m���A7�h9>I�qF�FL�ӱ~�)��#�6$�C�j�|�K�~����1^�f"1�qĚ�)���/�b!Cx6TZ�7��U��I����C���uu����&@�����͟\��.i}:e:8���>6�e�sBZO��Fj��x�,B�
��<@j���)���fN��5bȈsIK���֥�Y��*u:b��DZWp9()zY�h]��S�iA
0)}%�HC�J�U �D��Dt�[8����65m8)�M� o
7B�����H��3���C�sO��|6��{Q�a���vy���RS�+-�o����6��8�ዛ�V�´�9�Q�'�tڂD��~KP����ןq�3Y��4�N����YM���
�Ĭ��3/0*=H�׶K^'����,�JT� eB�*�qϠ��!�oA�����zgF
%�P)��m*ߏ%�td�������Cd���Tn#�l�������E�@*ͬ�[��gATQx,�`����q��3�T~H+\�� *��|d�t!t�0�3c���-��a�� �3��B�'�K�̼�!d)�d������$#Y����Pm�NkƤ�K��䴮���@ܕ�����T�$���[��B� R�6�]�S3Ϋ��1C�e�79���$��Q*G���0�1���y�:deE�� ��ͼY�i�V��/VBC�R]<��,ڷn=��V�QEC����6t	~"M&-���P+�<�:9f�'-WNA]UP�E��ǽ%�{�H�-ĥ5o��y����J����G���Ƌ�$0�$=�F�����
���|AڽG�r���!�W�wM�\�Өf��
��绹��|��>�g����|'LT���~�N�m�������|��ϱm8�v/�Je+��>`Y��	������,Ca�?ֿ��.;6d��
E�A�Y�`�
(��<��j�u8�.I�^
��6	�6���-@�+{qX{E�˒�A�r�[�v�,
��L���V�;�b�,�Ijʩ0r�<�6�,�n��F���ɍP�]�n�r�?6`K�:�H���U�S1$��Mz,�]\U��໚yQPT�Dkn	B��gz�s;���:KVg�l
��i����?��1�IRG��#V9��>�e��@�؜�*޼ק;��R^%L�l�G֠B�TljM��NQdf�O���CL�7��ך�?̣1@��,NS�_|���e�?��R����BV�d���u�d�^�tf�Q�g��0,4��x^7��L��v��dQӝ�9�r�&<�d_�G�;�MA�<k�iկ|�P��tw̖��@�R�N|Z3E� [-e8gF6���
�F�&9z*n�TC�٩Q{�'�{���AF5��ԗM���;��آ/M���W���#QVH��I��IG�p�g�!;-es����
#��p�w�Gƛ-_���;������N���޾��-���D!���Qm"v�G�����(����F
W��&�f~>c
cTÉV��l�O8��I߀��`�����,$�1ث�9��u3���T!�����b���5�w�^l/�dds�.��}!�M2��<��Y���A�+0�dI��U`�f�Vɦ��Kj���ɳf6��`��0�L-�0��ΞX*7�M�-�	�z6�.CŢ�eEGN��q#�dR����#F�2�����ӡ{4�l,���E��E���ڟ�CD���^f�z/~C^U�9d�o?�no�O��m�l�XRI�?>Л�gNf8=٥��c��)zp�n���)�ޒ��/���e�e�d��T��6cMg��դ����a4����&���h��]�z��h��o��w�(�g��OL8`�uÊb�h�A�W����"~�a�3LSlm"���i*��k��y�@��]%C�q��D���Fs��1�YD	��������T��d_?�g����0�-39p���(�1%���G�d(Լ���j$!���1���LMȻ?��s�j�6�����˘��*O�IQ$�}�����oaK�Id֧]��-d�p���b�,ل�DQ
t�-�ȇ������!e�@<�PH?\o]|�-��̇@��V���'��4����Ⱥ�	'�S;{���5��G�����������th��ݢU�?�D�-VG�����FI�S�f,��NDYӃ�͌�]tg��٦�`��R���d���-]��~^�\Zځ�7�8"=��}��|�0�L+� [Yn����`�y��`��+�o1`��T���B��S4�X�$��|J~�C��As��d����K�B��<���H���G5��ak��Q���S�'=l]!�7ù/D!˚P5�Mv�3_|֜\Y>�&]��8�Qʡ�m�/6����|�	�M��Ҹ��ֆBt�$f���_Tm ��37�h���,ҤC�b���W(�ß���t�>��%)ggڤ����j�<4�9k���0˂�/���BZ<��I�r2���$����Ɖ���OZ?�6Op�������N�ڿ��5CFt�o�'��յ/�A�u����r#���L~�$=Ǻ��ثqrE���Ys��\�����L��Q�|0(�p��sC�]�� �{�S�=�%l�Ln����ڵu����J� �t�p���d�3��G����Q���	^�Ŋ��)����� @� ��v=�vc��܌
��<��fz�&��@�����	��1�s���j�ڻ/����*摦޶C6����s N��6�؝6�U���7T'��<����W״aTV�g��n~Ԩ�em(|�!���B`��^n��� m�牓=�ntr9��:7)b�(�G ��o:6�>CG�d�G�^J��Q��\L��?P�u�a�.�t����օ9�$T�2�q��OL�gvd���B�㽣�s�N{�L!@m��b��n-�N	G��!���<dV��F��όS�B*NҴ�a6l�W���$�'Q��9����#N����<�����,�(PD��4<�v���vvk�aL�MN��Ur	�l4���TW"�fnE�Ҹ�2}��Ki�F�`�0�$�(�����L���~T�y!ا|E��R�quma��vnY����\Y�=�2ϲ���N:������sDj� k��_	�VB��ѭ'#S��Q"�9����=�d\��Zt2����0ֵ}F߃D.y��zm�h�ķ �{���K\=J�$!��_����(���*��'	�?��9��G"��บ���]Q��K��Z
��b��S+N\bzA
����Y����(J7T
76>霾��"ɖl�Ӳ3P��rSPʯ,(X��;1f�TlI��j�7���Ij%Z�sm �	��{�s����]�Ż�ä��qd�
\�U�x��\4�*�Z��Ф���'QI�����C�o��-Y��o�:�Z�|�NI�fДit�T�ܾF�j�{��;���R]�<	�����)�nH�ch#�8���(��ف���[w�۬y����{Br�����c�E�E���^���K��o�OĊT�ݷ2���4.���'l���<Y�r��g
�[��R���h�$� Az��$�|�1�hޘ�R&$�O�n2w��]�+��Z,H�����;k��!�Q.�XA�&ɮ��]�j��]���}������͢)�>q]�S�*�7��]1RD �(jE(��nC�8���'؞>M=,;�C���X_Մ���wq�s��3�쎎Ɍ6M5��h��\�'*Ä�USWZ��z�2���3�rgJ��'�R���6E�E�tB
�����LQyb�z��/��(�>X�A�u�.dy�EB
r�����eea�]-��Q�a5S�iW�ϧ|��{�ہ���R��D>;���4x6�
i�jj�����]��⇬�y`��۾��h4�2���T��]x(
����'$�xÀ�1�B�LpdO�SEI�~T)$E�P����$�G��W�_�JU��{�N=�dc����T�0Z�/��0��-�_�H5��;�v�́2~!���������)N�/������wڐռ\�����J�A���&wzp.]�b)�X}�}f�D�r��]=�>�E5�5�%�����z��w�<b� ���H�h���]�������uʰ�r��FEB�dB�p%ŧ!u�x3��|�>�jv߅m6���"��F�����p�m�v���3��|�b9؜�)�.X,[Mp�@�W�\��N�V�T�Z���g/kq��}/��c�u7��\Sul��5K��z�mR��W���r+�	7�'��s=T#[�+�k(�4W�k��m�j����8�	9
3�s�I�V��|��G2o�T�$�7=c�j5q(���&�6�8�0F>y"���~j*�0�nw�%U%��I.�Uh����)��L�fd2'�������8�w=�C�z5�xZU�z~I�N8LC���?��Ϝ"�p����_����WnBo${��˼|����!u�{Vf�o3_��D�ȯ	 d&M��p��� 2ܺ���{**w���y�ʠSH�B�iR��je��M\n��Ag�w�J���Z[��3�z%���Oꬬ�p�*D�7��i��ĉ��3=2�F��4*�#�O�������L���R�L���8��R$IjM���ސ۱������P����>u6����_G��Эm��;�Pr�{e��$�xkw��Au��h�6�h�b�E�*	�Q�%�$o�0s�҉�|i7�M�b�^�E��_S� ��%����j������D�:D�u�����c3�5hP����V����_t�'�x.%���� rY��>�Y�x�P��9+�C�L%��vb�*7Y�C�C�6��e�FB��ů��0be����j���A�'�0�X�"��A��_��T[��QP��>��=eDYd��!?��W����Q�t�I��u�]�9U�=�
�!/wa���Yf��)�+`��W�ު����Rf���<�[��@��rF��a��f�k�8?m���V\��xM����*�����G�wI�ӂ:�uVMۣhS��h�|�k-�������a3iz��$���txy��Q�={�o>�7QL�%'յ���{�dʛ��ѐ)ҪYV��S�&���/��-DD6����tH���հj�\]��w5�<��"T��9�(=ku�77��J��ۮ�,�,��	��E��,u44jZ����I,[���R;�K�լ�v��0����ޕ�lM�(�3�)!ȋI����)J��VV8�a|�����5c�EXZN�Q�Ci���g~�%�F���)�����J�ܔ3B�goT`��V�'D{��-Y%n�`�$p6^���8�)���v���	���]���|�'��t��wj���~�q�|�4�,y3��u�72Ww2	���/¶g�K�R	���L�:���cہ�hGGa�v�~�~q�uň����_O���!q�v���=G�@�J��s�4Y���i�'ʛ�6J:s�w �M��6������HQ@�����]�PK�s���r�`��(I<�.��$�������ya��c�	p-�������zF
;�����m�;���q�ț/��;��q{���c��iW�2v�A��`
|���ȷ�U،czny�=q ���Mx �4ݪ�p"!�������P/�_��Q�G���d��#�Z���C9�W-#���'{���'OG��Y���Lz!S�x�Dd1mf����A�v/�j@T�jxެJ����+(��$��&�BA:&�)P�y��c�6��Sz��Wƽ��`x�<U�۾Q�Q�+/R�U�qJ��ȉ* 7wwGq���)׿�&�F���A����jx�����咊��'����~|d��f��/�^���ľ�+�vO��.a��"��rj[U
���'��°ۈ�Ze�s��{f�\n����P��[�Ζ��?ʗ�@���0��$�
?��7U��"��5�S�U9�-X~��w��ߐ���.p�n	��,r���e�ie!�V����
Nj]Z�.��������ط��o�IYk&���E���Z��K���>Ɯ���V/�"�^������C)��r� �$�,�)�~�H��V��sR�Om���m���l��Y�Ɛ�؈~ �hSK�,�/1lʋ��9�ˠ](}JW.��<�Z�=l��1`���&>�T�� )�Q8�N_2�Ay�!:���{I3k	���>��o��E�$�C��i��Ь8�}Hź�U�jBX�

���>���иW*��ǔ@��u�=XM�7�uH��X�@�?p���:�K��3o�e���=u~�-�f��x]G���.��[�\�ӿkc�$��o��X-��	|��ƞ*CI�T9�-T����c�֮wQ%s^���u��W)�Ǟ��[T8],}��$y�;Ql����;�/���2��R�NY�&L:��D�����s� ��i5��&ʐL�)+�g�c\㐯`�^�� ���N����*��s��fP�
��1#X5#~Q�工�*%xZd�}�����d�!9��0�k�����m��ڱH�\{��>�����$R����/ �˜�g�T��s��^��z��#��r`����$ϵ����jyY��q����֊ys3��g,�(@dh��,��e�1;���m���.�dˡY��Hd���9������j�g��S7~��_�O�� ��ϐfP��m�=F�X@�t��D,�j�H���yM..�|�nJ�#�7
{g87��Q*�g�X�W��T�ƙ@�X����v��z.d�Ǧ�E��)u �]_�K�+_Ӡ����ǃ���Pٻ���j��2f��f���3m�]`}U�0hX�kI�D$Q�%fp�ނ�w!t��Q)�
v2t&D��!�E130���F�Ub]}!mɣ)�(ˏ&��z��=��wye#�:�UJ�-���N�ݑ:��O�|��#��X���f�m���f�m����h�bB��r�����Z�*���$�m��������!��B������$��&��=��y<��|��
����r�>Ǔ����ҽ_��֬�dg���P��@�*yF���:�ܘ@�.'sC ��'V�Z�"���"?l�j�M����%���]���:���p��vC��{�岘�M[���J#�L���:q�Ҩt�v���������"Y{W=�}յ4H���sP>X�л#��X�_+!���A��[	!W��Zgc>3��*�U�+���Fx>�|S���,��R�
V���pY���av�z>���LL�{�q~XҫBI�5���������)FFD4��9��6�1.ay�nۂ��L�*�y�������
y -���w.	�ٛ���o҄���TN��_��Y. ��,�,3��!S��?Ԉ�bεl��ɆA	��1Y-�%6-��5/#�)��
`�9�<K$k�" ����ˀ?�!O�4���1s"��$^�:(�b�*����� ���0���Tv�U��m�8�JjW�"��%���T�D���q��� Vs��37��ɇ���8�KZ�Q�W�*Q׮��~�HXz�ך
	pI9|4̸�sn�k����$K�Y�X ��ے@@EP���7�m�����T��_3��/D@����b���8�B�ܠ8JE!�r�!�*����Ǵ�G�֗rv��O���Qp�s,&�҅,h����	��v�ϒ`^�|�ٻW[�0�{���r�Y���s�#5��&�z�Ο�6�JK|s��)>4�XnI[��#���Қ#e������'�O�LJ=*EW�y�3ͱi�:��g��sL.O9p>��??��6s��PC�;���u������G�@{>]CMs_Z�+�����
S�O���j�⤐%H^=4-9���T�-���U*�U1�!Y,�S>�aХ� ΐ�u�N0��"w�m��{ZD��P���s#�����H1��YU2�L��P#T�;|�n`C皊jٴm��A󟑩�k�$�l��DlGJ-w�Z�t!GlE @r�~l]
+���-�>������Ά��Wd"g,�����w�uJ���<amr`��Hc��Ѳ0r��Q��#�>sj�]��		Ǡ���צ��`5�"�#�+u_�{h�� 	p���v�#�-�o�X�~���d;
�#Q$�1�p4��-t��6~6�����l�P����Ň T�G	�E���f��S��b�q���ۢ4��	�������t5+x̊�p�gX�����޽�BeE:����I�{�T��D����U��((ǘ�w�3GR;k�hrt�Kn�����C"��:�kO+�7CZT�#�C�����lO[����v�7[B���A�_]�u]�Z����_a��z����C���0�M�i ~XA���nuY��smX#N=�Ԣb���W@�xa�ӵ"r��������0ϏJT�m-�� �*P���ϗ*,P4	�#����a�VJ��`b���ޮl������i�J���֤.�p1��Z81�0Y���y���}b^�R�a���ɞ��D�9h�n��w/˄w�0^. ҧm���/��Z�h̍[��]�)F[�ƅg��{�-�ыUV���������:Z�.K[�g��P������[2~k��Ϫ���p���)�����]���̒"`z�1.^]�;A��T�Ix\�����}�|ebR��,9���vQ]�\�4a{K-M}a��zZ�FM�L���G�gQ���`�Ոߟ]�4!j�\�3d?N�� 3hDn�ٵ��;,DC]��u����i��1���>P��tbh,ޯ<����1в�i�QOB�S�B���\	������˧�$H6g]�V<��~'�>�	Q�Ng��ʭ���=;9���jd_�!�x9��2������ui}O�*���M<�:d�A&�  �e��U�^z�6�4]�j>7��p�gL��ld��������[���q�&4Hꗙkt��_+�5�j�L�H����||9S����pK�U���P����9d�L�q�_d��8��K+�̲s�k��ݛTp�yk|�16����_8�"����E�'ri�N@q���L�ǯ�,k����T�q�v���X5k�x�D�݃�R���{�;�4��$��\����'�G�7�c�_�� �GD���E� ʽ��5�gRc���)g��[��z��`�Ф�ץ��E1� U����=��c�%s�ʞ�y�[������_�Ó��`a���̐eu���h�ݺ~�������5e��J���]v���@u(~c�v9b������ %����?ח��BlE�>�{����	��o*�sO�pY��m�yJ��̌),:��-h֓v
_�7?�����΃t�]����ĭ,+
���"�*a�|�D�>;��FV�3w
�Oy���׫��.q���4}��2����T�0:+�������{��j�n8�3nN�F�J��#�2���+��d)#�c�@1���K݇��q Α����(��9�Un����»��B1��!�+�� ��h���7�eՆk6�u q��ъ�&,�[�ն�H�RAQ��¿f�	�<D옫��a�4�ݞ�͉ �T߼��K-�C�>ux��~��1� �[��� J�Jcwq��XJ�F�f_e�:��87H��[�DEڗa�.itΨ�%�#d�1��P�Jk%��w6����b:���ͧ{�B����k�I9%8Y�$>�� Ӈ��X��VN���F�I�7���m�Z���߳��蜰�WՆG���ާXJ�t���l�l���Tuɣ���S�P�O������xK�$���ItV]G�RxE�B�� W^@3ţ��좊N�O��QO�p|��ƅ�W��$rHׅ)(�;�+�;w��ﵩ���E^cw7�!�gb>���{f��iF�I/���n?U��ؾ�3U�h{j���(��𗾖|�}a]W���5c+�[h�c[�E�VU�3&'�I����I�R���p
|?G�-����'����Ny[C�]#�p��<O���5�s|��g�UV����5�`���q{� i{�:�`u'E��wt�
�3͚x%2�7�~��bЃ����d.��/�G��)J-��<=E{a�fΎ��p^�H3jD���m`i��
��ap�"dΒ
�Y�19�SE�U2Os4d)�m/���e�\��p�~���F��,N�A��p����[
���׎v��eH�6�iT�ܛoc�@,��NZ�?����#8#,H�5n1W�U�%w��������!t�i��I���Ј$�:"B-�=0A���g��qVQ�~t	 ����<p?�$�{�:���p�b��KAV���J����U߲@�Di~ɬ���n���d�Kz�I���9%��wm���u�L�׵Ԧۧ�,�-��a@�� L���#k,�	凃��`偨V�����X�����M��[yeE�P�;E��\n5�'�#T��<���}�'�V:x�p��=��(��9��D��D1>п�3=�#Z����9��W�� ����{�+����T������:��}��]��|�t,����
ձ�F��/D9h�Hd�����T^�����;�߫�қ��_�p�(;�lz,}�v�e��.��6+����n��;[����@{�ę�J�
Vp����pӖ���,�!¬kL*J��#��O�?5܎������s��7|,(��`�5��5 �
?l�$pR%ܭ|��u��*ߚ�1�|�����lj��� ��T���6Y�9��qSg&]���I��D�k[m���V�z]�ʙ���C4ls]��8���+&�y�$�y��}���q�*QP�7m_�烥Ccu�B3fgUE���5j|aw^��1Q�zSu	V�V1�l&��
i�f�?�ƈ	��ExH���^Fy����ȩ����U �?�<�fo�ErT#�������؅`�DS�,rx?C�
ӫO?��Lq��|?t�����燨��FY����ñ��9�Y�`�Y�Z��a�p�'"�@�B�2�\�R܅���t�R�k�ʋ�L�����(�b_
�,�$Ʋ�N2ӛ�|E>t*`�n��a*�RԥkL�n&%�"-�lQ^Q��K?RF�2�W�,"}�r���Z�Sc{h5TxJl\��f�z��>ΉWv�ZR��I
��
��t���Q[#S�.����}>|D�s��ҿg�E�
Á�+t�20׊�����n��0V�s�E���(S�Z�f&
n7.#R�q-�ag!����̫G��~��V\��]��Ю�Xtsܨ��-�X����>c�S �J���(�ǚ"wy���#��6����V��ԃ�+<z��q�y��vs�7YC�7�<���6;��',�|�݉=�}V�<�w�4Ӈ�ΨIД�ޤ��T.���@�t�	`D�M�e{��%�˱%M�_K�c}�t�u^h��=�IL�Ζ/���0��x�=�`�*:��<X�<�39�v�}�>o��a���xCE�䞱�Z�v	����o���l�D�Ј�^F����J ����p���+�����@Q3�׈;g~d����Y�����h��U�Ǭ��|�����{Ʈ�$v�BB�H��I��t$��W\Ϣb�}�L�\��(�敒
R�Y����" ��GyKc^����� �VI�������He�Q(�e&/%��w�lZ��X�F�FTn�@��L3���]�F�Ǉ2{�m��t)��{29�T�����m�c;�5�Ƥ�Cl��˺.|ۆ�\�@.a��� O$,E�Wl����Qm��������$:K�H���i����X�M�`ɋ�ldb����8�si.[�;���ܲ�:s�;�Պ`zsUP�/S����a�@-%�#�/p1js;R�ÅQߌg��&ąf�}�#J�;L:�I��������T���o{qJ�0��z^f�IU�/�a��\8ǢZ�)��!�{���>=�J[P��������."�
厚 ):ޟ������J+d���?�ԇ�r����Ze� �B���wI~�P��"en$S�o���*䁴�?�6����%��M.���y.�eH����D�9�8���mI�'۠!.�S[��J4��v�0kZTO�����MhJ�h.�I�R߳]\��$�6��b�|I(��]M��~�G]?�t䏟ڲ��:,^�m���Ǐ?О4����"�eȋ�Ő���Cc|$�*J�ߵ�K�&��W�h��]ƹ��S�=䟻t�V�B�/X��m�O�>��r!4��<�Zb,����2��w,a\�^�%]â��f�>vZ����l~�k�y9۰	�&�WV�Z@�*�M�����U�G+����)=ɰ��:k�'�����1�� ;�4L���]A`�j�
\�� +ӊ��_#�I�	g���E��<i2iOR�סE��;6#]O��H{p����{_Sʂr6B�v'���as�0Ėr�e#�\��v���E'3�,'M?��Z��\�]>n��&HS4f�[�bR���q�Q����8W�B��ܒ������4;͐�PYƃ7�^缇j�y�b�;*�)��b+�9���n!۾O������� �v�8�/݄�6��p�X��۴.@*Z�i�g�V0	31�m�,Έ�u[^x�Ԡ����b��cY'��@k�_����r^I�B*��~����r0c�e��>fx[��޿�i_�ӥS��1&�Gb�`�ߤæp\�W��LB _˽�T\�����y'�;3�d�����L�j?t�w�!�ՙk�O0޳��*��4s=�� �ր$�jz�J�ȋ`�!+�P|>c(ߒ)C;�'�Ri�[k�����l����l𰅡g9W���?go'Q�ʄ(w���2�����V$�6/�O"^f�MO-JdF!bw���w�S�C�1���"w`e����]J����a3:J�v�ԣ�@��:܉Թ�E~j69}�f�Ԅ�+ܓ`L����(�{�J�iQ��#�����L쟧��	 &��0������2�ݫ������\Q�[9<�.��Q-K�HU]G>:�@�ը��e�X�����"��A۟ai��o#$�Q;E��=�PS���4�ߕ_ժ�He���+���g��ٽ߉�C$�x�>�@�2�@�����a���'8*> k�R�r��1>�U����x�	�Bt����%-Q�Uˬ�g�I*e���
Mo�P�ywRf�rl���_��}�����0���	�H+�D��/y�|<dI6�;�f5H=H��Aϒ�+��@% �Hޮ޶�����a�`4঩Q7�ӱ���Ѥ�:Ϥ��XB~���}k������B<��t��gY--��cK]�ժ�e�6�MPc=��_�T�ȷ	��(~jl�cVb�v\�bIr�/b���;�_~p�R��'����`�0����t婰��VmR�-�S�R��qam��Q�/�[z�7{��C�N(" ���8���U����5��I@]���w�rY� �6���Q0^M0V}�X@��������'��8��i���c9�[N�&%��k?�� �Ďs�@·N'�k���B/�ߛ�Nk�ҟ�^_B�w@���u�F���V�W�\��F,tŸ�4H�G�����q{�Z�)>�������0wE��P^��{0�&tӜ�y=��>�8 Z�h����G����L��Mu�LE��χӬ|0=E�yYā�Jj�+���0n�:@�.Ci�_E��:i�"&�b�8��xb���� �HF�a�;%4��-���`�ex~xa��9o����K��$�i�Goܵ�_����� Z�,�Z!��z���K��E<�K��˒+3W Sm?=�-�������n88�-iM�sC�~Q�"�U�w����G�ty̨�MW�*|��5A������tM����VP>��$F�� ��.��ľ{�*��t��.��b|���ˠ�*����-[��d1��˾߉[��N�yX*�e}�����_��#T����%�1��Wo���1T��$�J���Y�¬���'��4����Ov��#kn���E2*���l�b2�}�G��|	M���頄��Z^ž�#w�i0,�7}�;�VE�/Zx���e��.=�+�k(z[�op5|�f���Ihn;�����2���uR�Ωqjt�,�<��t�S�^}.�_�3�#d��˱�(�a
?io�9�f��"<���J�l;���'M$}<A��m5��L��7��f�e�5�T�G_})�w0Vz��J�.�iCo{��DY���%�C��<���i�^�9�*�v�Wk���-,�@�z�������
���o�'a|���\`������ˁ�M�khR[����O�]9D�^�Ԃ�=n��$�uro����veK�zT�B�0�l&��;�<	-5��gGe���X��w�i	O+��_"<Ԑ{��nՏ�uv�@�d.Sݯ�c`���,d�K�fAb��B3�X���jbS�= U!���*7��J10xB/!!�Z\H����ѴŁ�sf�&Y���@7�c߃���"{d��J���^��Wx{��@W�2/i���nct(%�^�y��W[�D��F���q��m�-����,�/M>��w\�'�<��d̀�(fw�/����{a���*�x2�G$5�s@������T���^����w��~�w��y_`��j��6<�]�G�읁�B���=ME��Iq���Λ�N?˔bD]<J��G�D�٥D���l�A��<�v Y�q��1�����Jj_�8���o['�anz��N��ųϖ�Ɔ	��4׿iA�V˘k���z���Lf ��ni{����&��bŤ�� ^]��0�Ż�_�8~��<m@���@+|0U�o(��b ��]�t��4��q�;�m�����@Z	���Kڥ:���_�3�z����v(�i> �#�����Юy&�~���-�$�X�����o܋M�&i���L�������{��n�b`"Qʱ:t�ܱ��,�����|G����u���b(A 0�I�V!��;:�!c@-�>���.ZE�3�JsB}5��)w�B�,��.a1`�/���޺R����l2�e�s��"��5#�W�������dh��k��\�V�F�B
%�!�[5=?�oW�d�Z�K�o������a��?�B
��4��^jQ}�	�7H��t��ߝfQ�N]��Y�09r��g�;IuH4 ��ёIWߎ�!���e,P�*���wLe	A�3q������y��d�j?�"�4�l�33[(xv�46$��n�"7�\�
��5㊜�1_�O0���_�=�>bAn`y��7�a��2�`0��Ne4 �ҁ�\f�ȋ�/
l^ژՍ�X����g�������W|�
Ԝ���&f .�/��@Z��CC.s��˟�<�-�pk�����y-�C,*?ϽM��W_?SUΔ�K�t�j��E��E�c�K�-�Wbs8_Q3���ᑃ��࠵3(L�K�YF�Dm;�Gd-)a��|oyҀQ[R�5/ ��ru�E�q�/�Hr�,��LԺ�(4?��Z��֯oV@����Lu��O��x�Et|T2�2��A��N5��T��X�݄�﷬�	.��}T�l3q{��w�0Y�`iNC�8E��>5��o+��r\�Ix�b�?P����uŶ%a�Q�����o]��\L5�doe���p��B����h�QW���g��g��&�mL�U~/�왑�����r]!Nf��Tk� S�I�+`r��d(;�֐�w`���^��n5�,�K�/��={`�{C=�*��'�Q�2B4�f��+p��C���d��a$���5u��0?��������J�H{��> 5�c��dܼv�,�NQm��j��f���2��G�7�)��bM�-���]�l34���B9����H�M�Bi�-�.��!\ە	�N�^�/b������ɡ��S��a(����ln�c��.��$����\"i���
�`6(2H���H�p�ұ����h��#Ũ�����֢	��깞"�'h;�,��uIM*c���A�1a��L�
<n�u��X#W�����m_�NÆ?h|��&�-�kݶW�[�~�E�
��*�rT�b��Z(�D��ŀ����׊Xws�����pPҟ�!�S�����H���f^�y0���q�vV�f��_��9� )ג��N���+�̪;ރ�{�J��tґ^����пP�>��
�ZwY~f�j��f�lC����Т��-�K�
-���1X�
E�8���O�L��M��w�L,�QmY�t�7XlrV���G<��٧�A-��4�J�6��`�����}m�?�}`\QuF�v{xl��-��U�u ���2]�v��-/�dom�4���ɨ)_�JM(S^-�"`����Wٜ0:y�T��|O���-���%Z),��a;~ܸ!�WS����n��#������6d�|BjD�l:��fd���9�O-�[�lVkl���!8�[t8Z�IU���yA������x�s��˹W4\Ȕ��<5j�HU�2�Fo։|�C��F�R#�.Al��B��4�&K�b�����j[�}O\B��
C^z��)I��кK �*��V�F��R��&r�m��M(��;�s�{A��Zׅps.I4�Z��Rw��0��5
W.t��)��Q՜�n��9V�n�_�)|Ǟ��Lϯ�qyz�����Q��X��Ex��;��-�1U�:�:wL���q���.A�6�<���֐�	tQ�[��:�W=%@|B��"7wi��o���nTO(����-�")�}^t[繆�ԡ�Z��F���J1�1Qv:ϧ!�Z9��tG�܅�	, 2�o\m���!z�OcG�m��G���܍����V��]��w�+�o���4����W$�׌e)��U�mɉ�~#�@��.Z˅"12.x�"B��8�s
t��]�:OL��e:'(r(]������f�3K���÷�+_E�.-N��*x��,7&i"0.(R75v�wH����?�uX�T�!i�[n����<��YE��Y'���c �y7�<�~� ��=�_��$E �,#�mo �p#JM���7=H���fݦ|)O��N�nG����8��C��xH�M�[Y���j��D��@v�g�T��ě@G�4lҁ���*�R����Ĵ���y��[t�B�@xi֪=��Y7�S3�?H�����T�q�ۇ��p�δK2G~ɘ?���|��3bc���3��~K��	��d�J4d��K����+L)Ջ����H�<�2'=����¾�� ����h���vWR<C����1�?G��8	���a��J�b�ٖ��=s��[s]E~�>J}�2�1}�&�̇�����T�ƹ���o��q���HPx ���\�ʹ#�pm{���Z�`[Q��/�%��٦���7�.��{������<�e<ٖl�  ��pό�@
�)�Ȗ�DB����X9���,2I��#��x�'['���{]-���g4R��vL��n�<�T���K����،���to/�a��pO��6��ݱ�|�������.�`gv�jn����H�4vq�,8f��Q�>�g���R�zL�� �u�E��^ں��-��n��:�����
#�Պ��R`��/����`n	�K�19�S��U� Ow�Q*�I ��^��u�\��dQ�$�0�W�7���C_^s�ifW��gm���f�"��i}ǑڧJ���Q�1)�����;n8��yj/��i���[�a�5A����c��\��\�h nF��C�R̘a��r_#E����|vB\Q�ї��a�AT�E5���ʎ�N��[��7�|���n
�@�ީm������]S��<��OG�\� �o��n!�7M�D�pl^�Po�w/�������i�uK5�CRa`���=��y��M�������h�e|��<��^�{�=�*�|���c�s;t��y1Bg����sћ��K��NR�P����eWWK$.�g�pdS��}U�����s~~};�B�fc�Ds�s��1�6���d�'�ŁN���P@]𖑩q�F
�mla �+��{R�#�.Hю��J��P�f������O�he<?xғ%�J���Kta�P�Rn��J�9jp��v�['LϺǫ��@�Χ�F`1Q�U�<}p������S���عg޺�����igl�K	h�Vz"�t�}�>�c�e�� =���� W^�bM��&T�ߠD?���(?�E���M������Υ��]Q��̷�P�+���7ˤqb>�<��H�Y���s� y"@5��M��P��C"ؾ����nO��iBA�����Pp�	�۬��7�O/sk��Z��{��sc��WsT����0��E冧a������Iqh�K���f���%��I6����i��YB��Ț-Y_9Q;N���vF~��
ەe�����x@��ʀ"<��F�l�\Sv�Ǜ���y��}4.����_��ڮ� �:����g,����k)��f��`(9�s�#k�ɯ�<i
j�Ȩ��<p�����"�ݑ���/�Dj,Ƶxnn�7���n���8K%���B�q�S�c�V�d� x���c��!�ᒙN�>��n��w�ϪG<�o���<(z����LE��sC���{�s*T��f�w�lZ��Ta�ộ'�X�a�B6k�A^V*�t��k�%�	��w��rt�7e"��xi��u�ؠ��{d�u���:�N�)��,�t^�n,~�M��֭��}��Gc7Ũf�q mQ�6�{#k޿[P�[ɀC;��&��Lr&��Nag�ǜ���[�7b݉S���� @�n��z
�k��z6�%�K�S�V�g���F��*<
&�#{��~���i8���x�&��R>Ҏ��D{��+�
Ж��H1`Eq�ڬt>!�Ct/Ag��o��9�y�c1)c�%�Et�?lM|�_���B��U��zǛ�;d�E�5���2�i��L+�ͳF���4g����/����j�ŮW�Q+�w	+�ʢַl�|Nؕci�؏Z۷+�v�z�*b�Y��Qo�Y��Ҁ�8Dy�2�~^��5�w�Z�]����m�X�{�c7��5��^(��ݾ�������� �ex�ig&�y��,9^�VN4䱔�
Z�G��w���5@zA�I��h��tAOѵ�U�̽v17spq��I�;(����h�Z��d��N��|U�P�>I�-=!�Gؤ�5�$�jx���w6،*�"�~9x3�$|�,�Q�"�C5�����8n�P��
*N��4��5�&jjdbV	��]^f[,~ɂ��C�����\bRZ�G#�^�9�Z���u�WC�6��{��	I�X��+�� �KM��"����+N�5���Vg�����p͌f�04���������m�EAo-A�ଧ�!��7��z���g4Tn$��j��ᠤ�`��95/��|Y&Xй�����/�E��A,����{K�1~}��S]G�Y��V�q�#C�' Xz�M�[`�������bS�';�����O�����2���+G\��2��',wO)Mq����>�;U������&m�?�J�P+��Ԕ6=I���j)s��)m[��S��moĜ�F=&�쎽��
��/�{��p8ô"����uUdgB�����=��rs}T���!U��I�hj]4�d�Q�&)�ѧ Z�I
���N�s���VL���w9{:�}�9�?;y��o<5Ԫ,�F̦�~v��L�|E����M�7˴nkY�T=�0�kˆJu��	��H����$r(�K��Vɫe1vx6Z��گ�z�Zo���6�F>�2wuB9�����r��N\e_؇� ��3�7���·n�,S%�q:
gDt�k��%��������\hU���҇ƐA�\d��4�9��$�N�
���a~|��B�J �I���>R�/�E��,"l����:��p���V�*�����`��������5�C������r�+�*����l���k��Q�"cU�V�͂%=�K��1����h�AB�y��.*�W��㛓�sں�rkd@������e-9K�;�Ҷ	�47���Ѷ�$���+��Se�+�m�.��}�_D� H��1)��~�x�2�h_=���6�������菒���)B��cf�6�Qm���D��7�Z�������f�G����2SjX�=z��N-m����Q�����fBj����e�ϘO�D�;:���s�qГ��$���߇Ts?�x"C��ɗ���=�-SA���j�r=���(j�6�o�5 �K,�/4����֫D�����}�D�ײL�Ǫ~F.��D�Gt���.;޷��vA9_�E+T���@ �N:&��n����i�>�Fa�" 	�!��l�j$�_� ��{-6#��n�|��(�3	�����Z�c':� �᫃���e޸1C�3 �;lӘ�`-Wh�J��L�>��4v�����\6!�ܤp���u���?l ,ʗ�>�� Ͳ,�'�Z!ӵ�$
09ҮZH��%�P�%<_�K��	d����� Nz���Ma���@:.�r�z7��u���^5۽���7�y`�d��N�$m1o��5����Gɪ�n��ӎM�,�l�����2��Zu�U�"H]�D*���p��J$�!�T���mqⳤ�2qi��7
��v��`}	�k&�b�@��w�~)��0��e�7�I�0�C5U׿��,��
������AE�.�9,��qv�\�Bi����S���J��݅&���bگ@���z������gKo%�P~�ʁ;>T���@��v2�{`�L�����h���;����w����(F�Fۖ7m8p�(t	���>ؖBs���T��*\���%��ܧ2��IMmV@@�4�� ߝ�68*��SeN�K�o\$?����������5S�xm� �ӣ�:,,��
�մ��';¿I�$RLH�0��n��K
U֪BCv�Z���<�d)p�LN Х�O�k��� I�"�oDG���L�Y}����i��]!�O�"KM���NE�axv/�� #�B�	�e6��Yb��k�p���a�R�@�[sӽ3�b�\�paka���d@�%���>?7�0�U�ݲ��$����촷(����rn��z]������bN*a�g9��Iᅑ�A�Ng���
6�;�!�U5#��{M��U�����}Ǖ6�s��谎P��C�{�]�-�/x䁘�;rnM�����D��P��A�ƃ��/#�����6.̹�C�)a%6��4�1�w�B��۴���~g�H�Ѕ�m�s��P����-�&�nK�ɼ{\���O�.T�pw�Aw;E���Kծ���؎Ѱ���YjZM���8%Ң�/���S��;D������~��y5~(%�x�5�S��w�Ȯ��y���@���琮����d�\LY|��Sb`Uԣ�u]��tMRs�7g�W�1�~���#��
G�&e!�����Z[���r�6REϩ?7�r�u
��;�@�&qf���=1
BP��^F���5�Ps��S�w��ca�t���Y���� d=n�j.Nu��@�6���z]{�[vDFl��'��!�)N^hC]�6�s�� )*�=/���F�D����Q
6�M'���c�Ts�����}S��:�cx�H*�t_4e��X��%r���	�-@��N͖�o�������i������0g��B�3�D�ɵ�ֱ}�y��l�7�4B����I��(Fw�R��{�]��nJ*����&op_P�	lj8O����`=g�C��me�3���>gvO�$j�uܧlp�q��U�tCU:i
uX|�b�Ӛ'_���(t}j�F����s<��M�����̛�4��o� $Պj|C��]��
Ot�z*��8duq!�i6.n�6Kd䰂1�F�`��>���\���`?y�~Ї���6 o���p��릲�f@x�p�d�
���������z3�,_�M�oRk���k�V�	�6u8�)*�"�Ģ>-�� �P|m�-���)7 6�/���*=X�(���!-߯eÒ�n(t)8o��]����-�K����hL�f��ܻ�N��-�1ްq|�Ar1�sdg���X�]�j��(�ϐ(��h�%249"?Uؔ�8�ח�+P�v��Ro���,��S�!����lw_���aoynj�1�wԋ(AE�l�7T�e]����P5&+k�� ���I����\=Y]����hN0��	�
:�ۣ�46�4��(ָ����o��e%z_ލ����I���̤v�[zGk>�ӳ�`��CF��u�e�؊�8��m��t6Sׯ�7�]C�;_�K���i�� f����@xHռ��W�Ќ�ܱ���0o�N,䊐`o��{��}8���Mp.6���z�0@��a�wDa�����)~f�^�Eꜞ��U$P�!���:	��
@Q����M	s_Q��-c��f;��gLY��P���L6��o����B=vs"��A�đ;V�e��LTV��j��ӮD u!�)�}��p�<�o-��m]���$�>��FWc?U�����Kh��9Q��ho��+1$�r'�*K��@~C�>�	��;��y eD�	y
��.6ev��vh��e���Y�5(��^����i/����$�d���5�a�{�һ��w�L��T��J;4 �t�:���C�E"�v@I�3�8K}��~�xW��߄��5$V����+� � y���$�|r�U�v�"_γ5��B�׷D�}�����,����o0���q-�W��������9\#��.Чv"�T�]9�B�d��x󌡊��#K��w3L�׍ ��{�f@�����M�_�ZzI���B!���w@�����f?tL/2�3	���Tnh�:*#@� A�ـW�X u$ăNf�.�k�Qf�Z��Uz�XU���C`�
�ª���#a7bJ
���G����/B����eS�7��K�N	?�:o|�{��#肑��e`���2�=��	k�����	l���ʫ.Ѕ��F����� ��buW�"j{��i*��
q���t��܂�Î�[����j)tS��z�ʐ�����v��0�H+Z�;��ҌZ��)Qi`h�E�.�M�1*���o3�B$�hJ���͢�o���n��"eHR�:2���/�:�
��ֳ�	�SA����Y�� �M��]���)�˃�TCZ�Os��� ֌0b��O���or��������d�(���Ϳ\ �o	����X�{1�R��x�%���t�j;��>6�rJZ4�.텧nif�%���ߓޡ����n�*B��R��u�C���g��8���#y ��alԞ��g��Zm\(��$��4|�&��2��1�;�\��n6��CH8)��S�(!��"�f(#�i� 
�!��w5�����d�R�Pg�Rl��g�5��#h$�1��|4 b���@e���@B`(�3R�H͔jo����F�ь�O5�5�"�%׍�2���b���}R~���c������e�M�o�1��挵�X�lM	�E�VO�'U
�#�
	��vϣr¦�/��埛n2_�ؗ�֑ǈV~ܕ��׎.5L �Go��/p\��d��&��5�Dy�0O?��yv�P�L�Y�����<�3w�	�
V���J��bH���!�����7_,�T����m��dY��xgi�!�!)�C��D�?a��-�[a��y����o�FW3�mf�xͅ3'�Tt��E�fG�q����i��d�u�l>�1/A�ok�.�L�^%ܹ&�w()
������F�^�qwYh���Lv*�V6Z��W ���Eq�1ʡ�N���-��;�蠁6�3$ս����� zWKӮ.�#�v\;ҤU�P�w��,�d�0⃬�>��*�{�?�|�n��m=j>%����]%1�rLv���:���0���+|ٽ˭�o��9I��a�{���W��2��S����L`����Mu��^��άJ:�k�Y3��!��6�UN�vE���형�\.�j����D��Z��D��Pѱ�1U�T�/�<��@<�B>���%��eE�$���\.�E�������!#��G���L�~A�*YHxd���|
�p3uADK&�\|��>�;<��� ďz��\(�q/�Qz貰-��t�60y�*���k B> ���-|U�6�s�8��j�
�f�[��c@��#T�z>�Һ.���s]��w��O��2s����Ɖ�c�j�^�M�u#������"��$3h�	y���K��|��FZ�^{����5��:>�?e�_1�s|�R{�)XE��rTD����-ً��_	!��>q��싨 
4ɰL�g�<Z�[����i�z��Ϫ<z�!�d7\-���?�3ђ,��?c��so>1qZ_c�K?�hYR�f�!�'�ݚ�m��������1�@͒)mn HlΡ׸�e�}C��a��n=�DVt�2��%�)�9]ʰ�L��Ѓa�Y��
a�	�W�Y�u睅{�?��� �N�0�}�Q���2���`�	/4��w� *|:����Zx����l7vS/�w{Xr�#�v���z*���̇�p��/�^�C�f~4 HIǁ�bЕX��M�_O�u�BꞹX���\�v�<����A����a�hI^p�^T���89,����(� ��4��������M�����&Б¦ϟj�4,ɁRo�<)�&����%<�e �:����r4@t���(�V����է�fM�܇��Ƹ�Z�+�[�.l ���=����Ú�aCE�ٰ:�>pRTn�� ��|˟ƍ7C�t����%�P�{��\���AȨ�WE�W����Do]x.���Y@?��¿��ƍ���-!�8!�Y�֠�Z������R�qM��PfӂʣP4ګ��R#jfOA��,���OL���?]��π�&����c�x�4�kz��l�9�,��n�cn ��!�����֥�/���f�qH����Z���c�&'7 �,�_�V����8��O�x�Z�r��v��P��M#c��N:��N��co�����[�8S˺��4�����
B2���o�V�Ș��{|�Gdk q�;�b��-^Ki8g�aw�~�u�N��GC�%��[d�n�	s-���@�>TO�2a����:ђ�nK�b�����֫N���}.�p�vK�-�m�T�[G�}��Q?o �|nM�_��_�RBTh�Q�ܿ���h?y��������
��c����
�[p�.��v��#�%O�W��������T�����9U8�c	8o?~2��ڜT1D=��tY>g�+� �GFh�L�g(��>�I�K�<��L�zX�,D�b`d�ǥjwyD���2�CSM�+��{�\���e�����Lt]����4'���]	���r�[����l��/�65i�n����o&���۠������n���4����TV攐+��v��N�,��:{܄��Hü���P���3#�H`8�4������7�ߘ�:
Z ����Å5��7��T�F�i��������Ů|C��8�V*����K�*hz s��K���<��ǜ��"#�D�<�`��]�Ċ}�7�VQ�����HHKV��Ʒ$c�隞S�t�y�����yb+�Un
E7���@ i_=_)��O:%u�He|;yA9t���Ђ�f`�|D�I�q�� ���m5�P�[�!�9��%Wv��]���:��)��*�"�-����3�����w�Nc�R� �;�`\'�MZI|�!�m�Z���3�3��fo�3�lx�����)�IF���g��}�ú���<먑��zB��m ���i=@�19��.3ի8��Dx�2�*q?��U��c��=����Ի�`V�C��n�3E��.T�%�9q|Ѥ���U��P��߸��;r�H　A3�Mo؃ڕa�<J^��*|e��H��Q�n���-~�F�t�|im3αJ�.IIA_{hYS��gxG��448��ש1�[�����70L!����2Pu��k�����x�lDj��L����uJD3I�P�QFW'��6q���� ��$�g��̂z�-r��)/s�39( �F%�֑��PwC�v[�tL�Ky�Xa�ĥ����(Jj��!� ��%+�UL�#����!�"`�C���nv�3�41s��Ϛ�s���_��o�w���x�bO_tב�ߠ<�"Dă���a�!#��T2ɾ�u��Hݳ�!ߤ����>ɭT���5����%�5��J��*њ�M�`��=ڗM=X��F���;_��YvK��5����	��&v�[��HAګ���D�Wj�%3�uz��;(�wk�-�J&ŝk]�����4#;�d�, :�"H����OD*�3��$�	Ckf?�w��x���y���5`��W�!�K>��1���3�	�c�-�mť/�5)��Ͱ����͠"��xaZ��c�ci���3w�f� G ���,�ZG�Y2[<E*�{�����uUf���X(�
��z��%�3��U� �PSm��WId����� �=��H�{��NϘ�)�7=��
���ۑ���X�w��3/��� 6��a.���K橩L�SR*j��`J���$uC�N���Wڠ��P��l5�%���I�k���v�� �R�E�B����'`�Kt�GM��gv�]��f mIb�7�a����� vRF����0>M�4�<��#O(�c;+b!�H�Q{�6UG�O X�'K�8Mq��
C����yl�쫜�7E{%�2��"
�G�L�	���N]�	�ǃ{ɈÐ��ɁE�4J���l��Gd� 0D�HA��7�WU@jj��+C�3(�G1�\t�Y�F{�huY{J��c@��~�1�u��
q!p����M��d�P@����}e�������k��*X� ����߇���iY�B5�k@R̒�X�,�U�2J��1����y�ؑ��D�6";]�r�)�Z�o�ˁ���� ���k�'$�+J�pz=�'Z���L❅ ���"�,�`��ּq-�gT�B)9��M�EW�FKP������V*�Ц����2C�g��]8E�^!� ���F���`G��߅��M��������;��s��`��$�K�	���+�e.ց'�@�O>T������`q�(ۤ/=��o`����X�)�=&$�vB�M+um�����	�R���|PIj�	,�z"3i�X�>��C#|�ӓ���u�Ӂ@�=r.�5p�v|7N7Sl(�zQ�����=�P�i�%Uk���BJ���p�{����]�>�?$��M#��#P,7r��܌����ͤ��N�������(Q��}r�OAZ�[�����'��\���+�#�0[�R��]��vp����#���@E�4D��:�a�n�F�=t�"�Yӊ_�f��_Z�ug�+/A묬���!?{���O�r7�!8Y�:Z���"Qs.�jr�_�8�[j���6M�������|V��V�ϸ�p� �XS��P������Oړ�3';��@���� %�1�]R��_�����PuK�Yې��[����Ա������ �Bz�Ȣ*��t(v�<�hJ�^���B��[K/��q���]��,�j�zfwc^6��ұ��A�HI�4����tz��s�K�*Go��(_i��Ժ_L��\}KC�F����Pռn$�Bt%7�`^���o!~���i�`Uݼ�����I����)M�3�'a�g�eC]�;���/E#�>�����Lr�`�0FI!�*@ld���L��+�d �S��E�_��E�ğ��G�ވ��!��XjC�_U�l����fYT�� �����u�2��Ͷ��^n>��;S���7��cba�=��6݌L�@�x�
����S���W�_��\���=l���-�LlE����&=<I�\��T�T���Up��'u�j�oXE�H�������v{K�D7�b(;�3�3J̫2�@��	зl��V�jzɖ�˜ԞV~�"D�D����\Ş��cN���C~hڣ�>�5��k�Pe��-k�)���)P�n�)l��� �X�,�~���kM�k{;%�Rg=􆊺7�T(�8'#.�?��Z��c$W�4�,v��=JG�S?_��0=�x_��0��,�sD��M��/d
�K���c�ɰV�@�������.dDv��=�La�]�fp�x�)��$9�l�$�Hє������Q�Kf*���%��.�ϭ��ѻ�7 ���^�����g��k�>[��;��/�X���W����y"rX}Nu�������M|u�~�["���
�A�����tOڅ]uxĸ�r�eϕ������\����ۓ�x�b*E�7F�c� \��f8C��r��ҴY��� *����E�[�װ�'
�JMb����^t[��^s�B��kuZ��0X1ep���q{t����8�Կ���'=p���7:�X��L�c\ҥ����e�Qa��x�"9�e��ɣ~Db�fc��\c����'H�!/a�N)'�CHo#XJ
&xfQ�ڌ��^e�|V����vin���XL� ��y�UO��]�.�xc_��$���d������I��k��sB�S,����H�0��^��bJ�����Y��ǀ]Y"Zt9�����{.���}]�v� 5X^(�`}I6^�5���:��b�4��2����#���{�o:}زl�z]s(�s���!�x��V�Ng�8�jI��ݚ^_=��L)E/	9>zMZ�5�l�s���^F4��d �-�5��Z�b��6}���T��h �_��x�`ȿ]H�i�O�E�;�#y&�	S5��x0�	Ye���ف�*��I�^`�t�qU�s��Q�H�07�1Vio��D��D�@]a�ozlw�q�Q.K�7J���:�nP�%�E���:l�[P�0�:�-���f�{ppb��˧�lr#��d<��S'^��dTD�������ï�m��*���/���pم�R�ͱ�{���BU�%�ֽ먡\�uw����ĝ�\O;^H�_���(�B0w��S$���MQ�`\��~'g�;��K��՝����#����[ٺ��ɬ��ER���5����6z�,�#����v�Zm�X�2��J	��R��Tv�:b>ߺ!�ڹ���V��?��S,>aܳ���m�gD��ĜI�q���9��E���lMI��>��M<���OP��[J��!��@-���� �ȩ��ϝ5��ע_��%6����$)�j�~��Jq�*H�eZ�')78)]� �%� �CD��G�Q�0H}5ԺW�|�v�/x%���**$�t�jb���b3��Ђ&�k٦2g�s�0���P~8e������;L�b�	+�I�1�OO��s����K@���
j�_{���R���as��8
P�V����Or��%��fÆ/S�,n^���h}46�_̍���2t#�L?�E�������!��F�J�{�M*��'�<�� $;u�
'�����ҧ����d;�,�E�d&����Mهt�����L�S�����#X�����f!>O�lr�?P�QPF0���T���&��A3hS�M%�Wm��tp��{[�/W�:�Rw�M��� Y(tM�0�G�l�xxIn̔>i�ʕlD�)���>{_��Y����b_� GQ��������l�tfKS�?�Z�w�>�Y"b����<v��"�1>�u���ٝ6e���a��̶W�m�V�hƌ�%�~՝�k��]�M�ј�t��>߷3������&�ڶc��Ԗ03��򹄌�ޡN��71�ȰvMAl_�nua��Ub���]`���n�%��waEq���o^�@�߫ù� ����C�;L�œ|{-&��}��rCۀ�5��m$��� \��܃ɶ���ft�7�Z+��d��!/c�kϋ���'���pk1�(j�nQ2�+���ؕn����7��f�9]ea/W�E
��Y�yae��߈����v^*|�}�9����h^���G����j��$H��I�C��o��M膧����'�&�Dd�s(��%�ȧc�]�����s]OpR�py+}�}�^9��?49��H�����D�,�^�	��� ��7�<�����A��G9-HJs���#ʎ�ס��s��w�碶ݑT5� �83X=��o��9�B�{ c|"����;[��i������x����ᒜNjJ��Vs��s<�-�-\��,�?8���a��Z
�d��X޸�d]d��%-�*su�h���E���T�P²T^��WH��*�g:�Ic��ɟ��=t������F���W�$g�!� �|�Va�jF
<�2F2�O�� �@�nr� �����l�O���%w��8h����u�Jh=.��KȦ���?f�|�B�c~���~'B�3$���H/7� G�F�����s���\�{㕏&��x�-�֑��B����a�Z$�e���c�^�����oUҝ���	��6�$F�n�����RZ�bp�]5�R��E���~�?�d����3�=�/�ȳ�7x>J�X�� ����߯�9}ok8ب�u'$Y2�5�DH�����%�	t���:H �@k����lu��m�Z�![���y��&�ר1�%��Ȇ����wRa�j�>�e��Q;t�c���8�N�`Sm��:P ����eت���^�M*�"̸��4���[�f�#�bf?>�:��30�˫��fĻ�?�%��S(�n�l�Ub���ӯ�|O�
/>w�I�.��6p��<?4v��Pd]��Vl ���!{e��F��if`�^��a��ۉe����/��6�y��f��Gu�-R��M�����I/- �ɑ�k1�p��U��+M�y�Σ��~)�v�+]������9�љuOt�a<G�aC3�ڪ���f�_� ��H=/?@����'�=�>�U��̺>��ҌRf:F���h�85���/���_*?�na���-�Ї�|%�Zfn;)�ąt������')�9y�Ҹt��&��
TR�v��$V3H����S-�����w�3T |�l6��/g�����3���K���}g?��۬2��9akJ)[�U�nq^%����a��q�K��ꟾ���N�,Oo��~ޑ�%��=:B~�?x�4ȇ/��(�M3�a\��qf��R��m�`��4%�@�ɐYM�/��:�Pi�&k�C�L[��[Ha�i���]qGz�Uq-�)n���P��ҡ��R#�^}�4t�Lŷm��>��>�ɇ��C���,��9D�Tm�����Ѧ����؉���3nG��~��"�&i��~��z��`<���;�ƛ��|��:q'g��$�)�b��D�´O.>�C�fY���������V�9��?;�X���2A�!e�����#�{#Dd4*(����=�B%��Qs3�jc|�}�����r:s��s�|Gk���$��̵��9�x,��o��e_�LZ}���xk`e���_X��~Z����vcP�-����J[,$�Tg&�A�켟��Z��!�R�x.��ꅃd�T?���V�5ͻr�C��|;^��- 3�nZ:��7f��|Y�%��� d-�Y�q\��g�������lW�HD�Z���I2O9L�p��T��bȇ��	�9X9:9�o���.�	g���?�+=�Jߤl�X�^���WX>��դ?}E%?��+!	,m���AO�9X��?-�|�o˾�4���~�P#��'8?i�"J�����W�#����m5�A�*��iƈ_+�/���~}���+N��P�]P��l�9-���=e=?��P9���-�������C��Y��$�_�lEGC�\�I�z�u��7� ��RqtX��-|g��D����:/�{K��Ѐo1�9�&%�~�#I��~��G��.��;�9J ���3�SzWQ���j���E/�L��#7i?�Z�hf.��|M�E#޾S��ʳLEY2~]%�hq)��xέ�K�@��HhKF�WDQ���n�S]m��Z:���#9���!��/����͓G�xc�=���%���&a�_xE6U�UO�c�N8�M�W9�"���r�^sc��48,Ip�W����-D�5���3�%1�,��JDW�/�U��&ȯ�I��\�G`1�!��J����+6�I���bʡ��3�涢�
"�5pHQ]<�2mm��S�
 t�hC\s?c"����6��#'pD�
;�����1_>���h�8hUKyG9��_t�aFZ}6bER9c�c�:���Y�L���f���[�(��N�5g:WWБ�܃�Iv�����"�x�߷0����e���v�+��ѣ�B�� �E޵J�J���q7lx�� u���a#	�K�5G���[S�
5��_�u�E���
�P:F���(5�����h��n.�#@��(t���EP?�;E�Kg�攊��))ԀΞ2��ۓ����䷂��wKf��R�XX�������}w���9����"������Y��!}9�E���ZUW��	,*�Ĕ�6������̟�/��2%�5t��j}��z��d��qu�H�?GOkK��/}w�z��&�o���PO�M��-���((�e�����V�1��$��jf3F|���1ے[ǵk��tܽ�$�SEqH��:��_��_Xv���{C`�k'�$�T�ܹ��<����"� S|��b1.Z���烛o�Ki32�(���I�@�����(��#C����Cưl�66hI&�j�����3O��2�L��m�/��
�P�f>�񂝼,�G�(��y�����$��[nOq1d�N�ç6#9�}h��92�Y�`�1����Ƥ1H��u'�����1���W���;I��"#>���h��M���Y\d� �"��.K�XŎX,���_��n�f{�:�V�:�����X܇�P/	V�0M���9]�������g�����[nz.𺡕����/d���H��bp�?�"8p���U�:�X���"��D�F���������lm�: a��BR�A�g�?1�/�)�nw/G�G�s��Pn���:����7\���sL��4f~��r����$I6D[
�)��ցA9Wz-�Z����'<A��e���F�Rf�ʹ!����u&�vHpQd�p�:�P�wQ���T+��5�݅��Ax�rN��Y�z�����̓����#�B$��ۂ�[P=-��Z�;Є�S7k�D�yW᪃����qlQ�o2ej虂�t�]�D�}x�/.����XI,�|O��Zcb�ύ��'է�HY�)��
zMY�#�����,��%[� ��q���:K�nW���|�?:n<ݟ\9>���_�]*wc��E��5��-f+��O�����X��p�t�0a�'�s=���Es��u�r�P;B���2�F�!hh���Ð�;wU�֫����%Ԝ���\�>��"��e�Zb>a
<L[�>��'�B�I��`S��$ͧ��\��L���u�)���Mp�w�C꒮~��j�(!���8��2X ��ll��Q�i��q������ѕSv�I�z|�P(����Uq*d=x�o���G9�G��p��S\��n3�A�}�R/I&6K�0,}t��^I�.L��@���W�9R�7B3�k�����ħ��r��!{�<w�1�|�0q8kq�+��Cw$$^5�DT��r�\��0_����c�;��G�i)�x��z��	l��n�]/{A��P����^폓�S����h�r��̩�K�_������/ApP�w���"]@�F�|�/�-�;
.s%��$d��^��;]�����gG���xE�x�'���'0�Y��;�cJ:��$x�A4g/�D��r�#� �+���#�(y���Y7
Iqv�+���]H��� $���Br��./�s���wR`�����my!-���U��"�����xҠ�t����6*���s��e�����`|'�g��XOP���?�u[�ʪ�-�p#'�;�V���aߕ���U%��ק��6��x�_�Vܦr�Ab0�(g��7X[͎G�4pdϳ �I�� �����o��9_������<�7��]����k�����^�i�kc.��
-��P/!p|�G��f��o��ڗN���)�BI�6��3����(p����tH��ڍ�1/����؇�?�"���$�!:���C� P~a��cA��+��Jѿ����!h���8�ʬ�M�Qê1ER�_'�)Um^�ڦl�,�ᯀ#��QfWk��zEs��\�+��T��Q���t��KϨ]�q^uFt����e����sz{0�ȏ�|�oV��#�y7+c���u���ޤ��61� �4k������g����/�*	0[�)�@S�;D���� 'X��j�Z�GW:F핶'SOխ������,��Ї�A!�B���{H���W�	�5��U�Ϭ#��Sj& .���a��?������q�k���U�1~�6k՛�Ǯ�@E~:�6m��uֆxD��ǒ��C�լ�xiWW\Ś����p`�b�eae�e�4�0΃dr�ڝ���+�ͷc�g0�O�+��Z�fu|aH$���Q�+_�����<+���+�cV�[3em�Hn�M�2�^�=öv�-8���.2���r��M���M��s��A�q�r �M�7^O�����z�#?~�_�i1�pG!.]��D���{5�#������G;ɜ�_�F���>o��֍�5{ny���ȣ����j �h|�3��+�%�W�q8�ɞ����i*��P�"��h�����Z#Ti���@#7H�D$��_���Fp�:��bg�c��Ny���.D�Ji�.Xq&H�⧯�ϯ�3%w���P�
,*T��q.8��>�РX�Y��	e:��n��K;h���a�d>}�(�w|�W_�Z"�xdM}f�`mג�������/9�1�~�?��l�]���듥Y�&��21�Ln�1��
�Nb������hu�j]*Y�q�gT�wPPQ�x�xH�Vj�N|*�!U8�@p?C�A�JL�����l^b�h�r�M}4D+��N�K�ª{���{���C�c#�c�F����=^�߹7A�K���`�&�����Ű�	m|]H���20BWi��J��HavLw�/��	�4�[�_^����(���p�K�c݁�08_�S
7K�k���ۉkR�r��P�z�U�߮�j�5�Ţ�����T#W��T��|D~NW�DG+I�(h�����3|��y���WV�js�:���&C_#@L���_��u�6	�(QOLV#IE�1�'���\�O�^ژ�x^��s��W'ə6�o��p�5� ����_�v����N��&>-��57��d��S7Y�50|�6b*xp}S��)�Y���23�>���I$�Ʊ�0�
?����4k����/?���s�X�6�nl����%�H�y�E�&)�_u�ʨ�=��z�,�Cz۩{�M)�0l;IV��U���&��o3'��B[�][Q?�^:0��>��GA���5T��IB	�����$�c9P�-mi�G�ƺAN�?(���_p�8�$�ɓکY�j�|N��T�@���?��M��m��k�aCK�d�א�P��3�F]�P[}�N�����ђQ�w\��w����/w
|��S�`�@#H�/��y���Xj�;�e�Ao9�C�+�����XzP�d�kN���@]�%����6�m^6�g�6��-s�LژM Jf�j.�(�8Z^Z=�	�	[]���WL�䐽�M�_F�"|������F�U�����Q�I�!-��\�5�㏐B5�лz��.�3K���_�Lؖ���Q�l(�3J����ɳ y���>����>����z0���8BB*��|�.��9.˸�Bp��U��Rӆ��B��o$�I�]�@��]9�\�}���������?d�Dpa.�H��3������$�"��-�e4��n����QBHp�A�"mER�r���oܞ�wk�3�8��H��E��L��7�\��?�b¶6UB��5����B�U�b��y��#���ShT
��͛t�(<��a��.m��c� ����pXu�<��Hw������l��d�Y3���rK;� ���~ꊨ[ �N^
���,��0��O _�W/�����!D:��B�&0{��%�]ufq��'�.�R�jƺ�
~�h�1����!��?��Wŀ����Rmb8S��E$������T�M�M�{�~<��§���MihiyΡ���?����ʍܩVPR��yo2Y�4̅T5֙Y:;�vPCX����`�PĐ �Yr9�Z�y ��wD��g�1�agM��2�?��F�������+��u�2��;�)C$c
�e�E�P���ar4wV����^���*,$�!0�q|�{(���B��t���Y���7IʩK���������^�h�n�YRe}�!���sDt�۫ͣ�7*ס�+� �p�b\
��%!�7�Śv;��5x�iq3AYL-q�%�Z|�f���u4G��܂���K�H��+Sa�Foj���@*ʔ�TW�IB$d�%N8]T���l ��m�F��k�9}ۘ�˭�����{���H��_V�T�9;h/x�\��V��4��50 y��g$[��sR�M5U<>:�Q�:&�jLY�U��5��]�1�~��LDGe�:���|"G#�Z�$����П��t���S�:˙�>]#qp���J/���9,�f�J��Ĭ��? �q����ȕx��,��7�o�W8�Ζ���XM
�T"o��NaǗ[�}�g0�����LY+N��1.�����9=_9L�����>x������ &S�[�����[�o�IY��6�*�~�)���?J��m4�5��8�f��K5ߺ�pG�LN�I�����b��>�L}��Q�'�8���YEu��t2�L�o,Q@�yk�:e���C�]�h,GZu��W�w�i��ɻ�M����F����]ݮ:��o���
�E��AͻA=�-�0� <�a�80��-a�/�S�������G43H��M@4؉D �b�4~���~x�t�_��wn���{��ËĀ��N�.N+W:�����{�= n�fP�-��?:=�HR4����:�\Dw��^U �:�9���/Y�!����ŭ(s��Y�y��so���Է��חZiXs*֔ ��&#7t���u���-��bY�,�%�3>je��p	�-�~���p	�%����6%p��i����#��A��ȫR$ˠ�+ڏ��rn�p�!@�Ϲ��2"c�Sw�
x�18n���EC� l $�K ��3�0�0�ja( Yc�_&+��5X)0ՔOqE�(�_�4��o�1i��H�B���L"r�B�7������>/��*�`����50j�9jL�QS�w���~Q��EB�$�O��.��:\cT�k�`u��)
�r�>��e�3���$l�{H15�Q�78���Mײ֢Ɠd���ԠQ_E=b�FW�dF���dʏY�ˇ���_��U���2͚�� ���0�A��M*���ȟsދ	�E:�[i��T�ǽD���Z�l@�:ܵ�`�?��U�7�{�l��+J2�����_.���2�V�8����p,�1|�)F��ؗP��!�ܠ��\V8�0����~lm���pz�Y.��١𒛚����Ȯ�{1i4���#!�?���
��,���Z(@	�g��s\��L�[��܊3��������+�0��ț���VՑ�����p�f��h������S�4�@��^��ϛR$<u;�G��z�!@zl���L�	<D#(v��x:k4�7������y)�4�`EϹ(���ӝ���@sgQ(]������>D���;<ۋ �N,N{r��P�����A��� ��������PX�uV���`�v+�XѧB�e:���M�E��P�@޹��N�3�[_G��w�����V|�[m$�������0B�t�
�c��._.ό��NT��k�����
5����A��2�M�D�r�a�tJ�r�����s�����d�DD�t�s����]иd�;����m+�b���A��u�\�[�W����Y�8.�+s9%NXq�%e�Y#FG�}'����	X;5����ă����05 9\+ˠV2Ƒ��@�S�:Th9���(�܍��:{�I��o�	q�Bj�%lK�\�ڗ%&Kn��@��Ӗw�]�J�tݐ���?+E[��O�q�m!��M�&o@bb��� ��R�!�ov-v}�|DA����i��!.<�sZ�I��M5�*��sH��B:�a�wd�ߍl�xJ=�V�Z\���4w)�I�Vhi��t}�GB�K;mx������"y�٘��>�-6���[�\3�J*,��v	Ы��e�ϯ���{L��5	T�r�E��a9��`��Zq��	.�Z#���	`jBj���x6)g�[Z�m�iyug�z�ו�d�Qm&t��B��D��s8iN'�� �<IO�[U�C�C�C��Tݶ����6lْZ��}ƾ0x�7�0Ѓ���<�I�"-�y@���5�{�_��~��J�7�S�6�i��d�����#ҢB��`KY���H���� 2@���_C8r�T��Q����+$z��.�o�뾿ٰF���{8jy�+]|3��>�C��Z`<����YF$�&^X[���-���Ҟ��(�+��^��˷(�NB�Ih��Q��X��pZcåBl����ptG�_y�Gܙ�l��~�)+�m2*�?�T�2���Y��8�������̒�"
O���&w�aT)qt�� U��o5
���~L����������!K���)^	d����1U��ǯ,�ʊ>��嶣��<�����y�z���ca=��%�������Q�}6/��G}};P��E�N�-4^Zo��ң����fC��o��O��K�F���::�mQS�`��%v�����D�x.3�XHEg��Y�'I�R�;'w)i�r�� i�� )[�b�奸�����^�t���B����*��M
Q- B,�vW~a��N2{��a��,���N��2�� p29�FNcQ'�gS��zm��*���,��A*�:�"��VI�������o�Q>#��&��Bh���t�\e�)�x��1�Y^9���@��^�5�M���)�^O�a[�u{�]2F/�K����˥*^H��n�
IV��-sg]H����`vъ>NVrX�D�j7���\�R���=-��q�brZ�5`r�4��@ߧ�����l����s��,�\��0Բx��dP��1�� �W��aL�K�������y�b�3DS���UY����|�1.�X`>G8��|��rmU�CQ>"�R*���Ǘ{���/��$�A�8pt�'{�F��/������l���@���w��J���sN?��OL2�-�����!Y�GTO���B�Q�ꔑ�?x�gE� �
lh���ܳ`�T���;l�մc�avl��d�Ŧq��-�V!yƯ�!`Px+Q0u��S�5
�ر@�Fҿ�n���z�K��k��i\���x�:8�ؔ�?�©��0�����H��t�d��nRa�<�~�ŭ�� S�"�[����~�s{��5��az(߄̖3R���Ћ4��������|����u| ը@�l�����w_%�?�!t}��!�V�okU��5�����3�Ρ�Y��_pN�'�c���0vc%�k>�YJ�t�ӻ/y��
ӎ������W*���V�m`���yI��7�$��S}����l���ݐ�ţ��du�ĆO1`LH��ɾ%)ToR��J�AU ���N�{s�"�n�� Xo��8��]r�o<q	���q[䧎&�a��5�0�v�Ā��/t�W�,�� ��.[�Lc�tGj�l+�Dx��#���`���W��4Կ�T�&@=\�mrk'{g�`���^/�^����w��u2�6k
=��������d`He5-��JJ>�ۉ]�a[�x�0�2P)�{���e�ruz�����a)��gZ�u�*#~B�r��C��9�^L�ܔ��!���|~�BRA���mW��5���=�����R����6��f2N]������� �Wi�?��6�$�i��H�^���nJ�����N��aL�����x..�X�8�I�����eUn�=���'����j,�Tj�CW�|��M,�;��5���]U�:��J�&耡�EU18I���E���jڨ�(�k+M̑���n��BK�\U�ҳ�wVȓ�w�@4�_L�`�2¸, ǾoK���/f�U�(�y��=��O� Edk�N�����o!��G�������;�>Vt�57�e7���偔	��q:�o����p�^U�6M��c�u0z�7�L�!
;��2����ӽ�=1��HC+E���1�ޯ��ԩG�'j8т���H�j�tI ,�]|�4��]w���JG�
g,%��#}��T�vS�'���&{$��C^��q�ߏ��� ��P�KC���ۙoԇ#���ַ��(��!��֯�\B���_�T6�0�͑(���NyR�:l��hTP��)C߄�����1�݌-�wc��^�"��Co�<G�q�����E�H{v����z�VB�\LJs4��Mr�[�O��f������4����w������E��fx��v��r�z_0E�P�c�bm	Æ��h��52� a �����U�ٳR�}Dr�vnq�DyaR�·]����QQӏQ�v�X|)�`hpK��-є�����<�Sq�Jִ	m���`���1�i�K���A��/R�/�t"��E�5�I�\��EVu���_;lMB���RvE��to�M9���W�8>ٕ[�����L�[{������]��쪻B���G���~R��#j�:��ZS�WDE��p{�4�h��9���9K�\S�&��*��F�"� �7#	=�'�u.���_��l��ym$������H3? E��Ѯ�a��R�T=��B�b���^�3N�?��B����_�zn��z"�����4"gY�cmd�bEX�M�=Ov��8C1Bc�\�s��NɶE�[�a&��-����F�����v@U��w���Rq*)4��ȝZ��\؞O�ۥ�KJ�Şـr*�h���"�H�)-��9�C7&�}.�\����u�O�����.��g�� ���/K�-���l�*�D-x��L��4�IɇuyԢ��1�T"�CGg��-k[EӢp�"Z2E�I{Wl��Ja���ss*��i�\螜����6���4�ڰi�CꞽVqX��t�0W낼r9�~*��ZQ��Q�?��`������� fz��zg�C?�7�Q^��WNӄۋ�߀q�N���/�v�#Iy&�2����꾬t��<�a 3�<o�L��s柿�j�6Z�%{�ْ�Z��̘��=:�%B�%��)ՌP͜�ӏp�t����5Ɵ1+3����Ԛ?H
~*C�n����V���3�(� ��7T��Y 	R�Vٷ}x=h�E������+k.rE�C���Z��n'�	ƚ��� �P�r��{�Ɵ�cb�5�¥����}���K��l�q��Z ����7|��5�w�$P�D�<q�&����8ꩰ���a�G珱�4���2f�k�]u��Z��Κ,�1>��TШN^��\��p�%D2�Q�貏r�y7��w��v�>! �gL�F`���1u�(�Ί�t�Do�am�98�F�c+��!�څu1p�BTH�c0]\X�Z�K���{�
���1�	s~���O�'��OryOL����QS'��Qԭ��hxX��������ĳ=�t�'�֗�v����ͫ+����̂n��ԁ�_��A�W��pӛ�>y�yT�1UV��J
��o��E�cܰ�M���}U�]MM�����p�ls�A2�D3�r����M�םv����V2 !2{��W��a;~���3僘���ž]�ϻ＿܂�n^I��-��v�!+�y�nZJ%�ɇcJ�̓���L�@SO��^|0���Գ��ޮn�Jzef,��>V8�@��W�
9~�����;�Ҟ���J'�U��*�<�����%��3��'A��g�������`���S�I>j�ͪC�F:U�hNV^�gD:vhv�Q?�����P�(F(qH*�ty�c^�&���>�)���2/�=-?�E�egr�A�1���R��1�<b�2�Z�g�b��ɭb�lx�1�
�:\�\QY��� �V��%|��`z5�W�<7/QT�&8T�(�q�^��x-E0p��ܽQ5�Ӟ�vva��x��sd�@ԀJ�Wv�7䏠�}E#z&¤�Q`��O]��c�1��3m~�f����>�7QS`^:����q��E�n�b�\�A�]�U�Q7����w?-#q���)9�n����>$���Y"Ֆh���KC��r>��������v���A�\\�u�v��[�^�Uoё&S��US����_썴��R�\�1��Y�&��c�C��Z}���,�b��.����1>MAQ�jZ�x��ĢQ���*�-
2d굱nNѨy�q���]��B�`��Rn�����C1]��5��a�ąo�"���(i�e�3��K�HB�7�E��*��n��?��8�����ָ�+
�]n�p�~�s��#��\0dK2ߖU5W��0�[��+�'ƣ��_���9]�����~�S� �o}if��x�3B6#hT�L&� ��c@F�$�"F�8L:�������Pa�P)��$����Fk��m���h��&&��0�$�d��0?�FU��E��_��ݐ[L���� �,|��<������w�[��N��`�b���zI �z����oZ�&��s��|�mP�K#��:b	�M���5�L��K"Kj�+�34�`��X�����{�n�P�@�u CEHMꊶI�H���|yٻ��Rv�2����E�B5�7��k�ٙ��۱�d]^B�s?-^��g����a�_��r�u��,?l>h�%�ޭ2�W����󵰦��Z>0�#k�`�l0��I�_�� >�LU
����N�ҩj��r/4z
�@�w�f�d~<4���XY�_k-�M[rW$Ä��T��_�l�)����4x�	+��:��B�g��"7��e�4\y��i�`d�\pʲ|?<��F����cQ<�Ͳ�M�#R�6�%�c>�&�	&�8����;_��(
�b�<���>ZR��G�\C����h׆�� �?촠TdQes����M�4�u�OO���1\�q�W�Uq�Yv�.V��pE��|4�
��#�"�xُ�%�R�/�4�On�Ӻ����3���UMu&��b�yt��z_\��E�M�\�lP v�T8N�#�����W/'��u8���2˃;��GO�$m#�{E��m�K2f�W��J��wCr��I_Tf	�}Ī;��eH!�q�U�*��R�L�
�D[k�V{��3P�B���x��2�B�1w��:�7�ਛ��|^�ܱ<-��}2W*q$Kmo6.١F���%�w;5_�S������f�wD��fMԨI����JB���ưn"�Ro[g����trF�
��1`�1����_���*��s�5����0���A�z��tP�y@�F"A���Oe�;�4���ŵ�٭3������g����*�w��7h����%�Έ���;
0N,�]gJ���ܤ�h���Is�H��J�VW��j�u9�cQu��u+;-�!�s*�"��M$9�-� O���
�J'��Q17K����h��4�I%����P��׬�Ɨ^m�X(F%u�`�hQI����r����ey���[��5\���~�����t�/����p&@���M�0�n���Ձz�p�/���r�A
��䴆�ŉ]v�����5�M�t����V
��Ty��g͒8�R�2s t?`�4���\&�e Q���,}���{�锔�s�3}-�o��c��p|B��C��E�s��CrS8�O��6.Xa�ҥ�|s��F\m��|��W�9#Z���z� V:|=�*��+�p��Nr�BY�?��r�'���]EN�)�����ﶛ�Z5Q�cD�e]�p���ی�u@5�7���erIf�c��V�� iMYt1.|�	N�^x�-K�������O �A����O��=BR����ə���"�����99�**{m����C ѷ���b���6T�X��G~�}B�������B�+L �X*%����b��F����Yյ�c=�p��%��ۻF����c|)�({��	eC���V>
��1��|I�c[���Lcӿ�d���'i�Uc*�@�oo^�j����I��-��.0n�O�=�}��X�
EU�ϙ�y��\�7��x^�&�-H�?9�����9lu+�]��iI�<��Ya�w�cڻL�3�]Ԩ���Ɠ=��!�m��1�J��t�9�m���W*�і�Jf�>�?���E��r�9,Z-��zl�l�����yVh���3���C #��|��&�K�^Nç
q��l���Z,��񣧻���Kx���!0[{�6(#��|�X?���5�EV�p��<q���%�Km��k0ӺC��������EP�F�/퐅�w%"6y�4 �(�e+�.?JtI`L��` �C��(�y^7y�@�D��S�~h�c܂�k&5��0}�%E���cρLs+U�1�g=W�wj�*�tV�K��-��f�m��q�X��P�t~-o�
qW�Xyzx3*&Q�@�9�R�k�*la����`-O���IM�
%��7�ۨGN��N�_6���*�HXN��ɬk�F�g��?���(���I��޷P21�y��R�pAzt̾	DG޳���MmKt����&�`�١�YČ�u�Nh��(Р����Zb1�j�m2�"/A�[w`'�a�����S�iD��`9�7%8�ua��ܿ��Q������XU�km����ƾ���_�j� ��c�\4>蠬最|�{>���-������H�������߰Ћ$@�����YY戓�:q���ѵQ�u��z�$�I:���Q7�ކn�[���<˿h��yk�Q4���eܛgh'��Cxv>2�ӶeSxu~�Y���W���Ǣ���*m�!����l����){j-�t����	n��+��؎�*K�z�g���Mb����<x�ϯC��r��7�(��N�v;�$-�0�)��3b_M��I��[D��ڢ���8~Z�<�[�Z{Vʽ�+�X�*M�t#��Xy��_
N7��k�ٵb�S ��KXj]�tZI�w����1�=G:���4��g�Bm\9i=�C"#��N�@�V��]�r#@SQ��PI�=��٬z�GS!p)},4i�|�z|�+�T���n� �w��{0_��)�Cm�cw!2�]Y��jX��"Ј�uvhwU�^��I%��������rl�R3�P?&#h7�u�}��"��J��ԕ�&��޳��b�8Ƴ 8�xP��,�3�ݺv;�6j�3(C�6�aR��b��uh���2/���z�%��9�<���2*7����"5��ׯ:5Í��M�JN�[�j���*�0!�>�z��v]N�D�6td; {6'���K���fmcѦ/B�S��h�b	P��=4�j]�s�Op+:no��G���٨���u$�ns���Rَ�����Jw8�>C��lk�E�\��� ���]h�ko�ڷa�t#E�Q#km,��c���FEz�W��O �	
�]�2*���Sǝ�s��e��\WKaO�C�s4�2�4��L�}m�P�]�G�K�-,�h���	(��-ژ��u9�x/)���皻��Lțy�H�&�h�q���t�	�qmZ�m!���K_���d٠8_q����87l<3)�Q��˥��a���J߷���hIr�3��w�؞��ٱׯ�02�ЀG_B�w��gS�Ӓ.�h['$<I�*���?�N�-�#�YWǘ�������������a巴,#�
g*1_x�P��*Cn�ਅB{�	�S���nET���T�VX�o���q� �[S�j
�s��L*�y�S��yy6��B�1�5ۣ��o��Tj���ɾO������3g"�L��%	�͏��]!t�����n����hvo�����m�~����'�##a�Վ�;yE�jC/�k9QI��jv�X�����SF���J�{�9\V����enl���yV�Ϯl�"2����ݰ��-!���c-��,m��{Ϝ�y	�Qc���a�Q:���"��=�
�]���*���ڶG����؀b,�]�0�}:�j�P7(��b�P�#�&��D��o�n��$:Ů�ߖ����Lz1���B�������$lh���,����}mިbW|ȯ$�d��#E�K���� |mQ�Y�:�%e���'�s�滰a۠�wU��nA���P�K��%9dHd��ğpC�^[�de���1e\��l�W+���D��!�;0b0����Dy�/T0�&����e^��	S�^�E�.���Y+���:A���ei4���FP6ކ��.{3�z
�4 }ú��<gWKwf��:k���K���a���I�5�4��cv�Q��e��rf�C��#x2[ن� 2�P�	ng#��h
�Tά(N*��/Z;�"��/�/�,͏4J@'�7�z,p�j�
ze�t}`Bj(�K]��i�č9j�\� ��4rU���6�I�֑c�z��,�wF:Pf��>O�����m���H�lN8��}dҒ��%N��-�v$��}�W���1������"-׋��Jp�P����b�"�ki����������*�*A�jj�5nE�4RJi��pzUD�'˖@����Z��N���3]��.ǎ�Q�*�3h_�F���	�B�Y_{���pl��D��;�c��͎}$�����!�8<!!�w���Z����T�Bm7��X���.�9�T����iX�Xu���а��<P\PD�R�]�<i�p��a���^[��焍�%S��r���-a��Y�f���P�E��dr�UWr�]c�Kie�m�Yf�L��]B���$ˆ�U��h]�!����*P�y�w4M��X�+z�!p��ek��:o�e-���N�Z�1�
��A{c3���!��y�N�3ۀ�e��_C��5���ӝs�
|��i�FMP�/wo�4���i�B] x�6�W8s���AWC���[��ļޒz�r��2���7�(��u�g���D?��C��o��D���IL�ۖs�@Y�e���#r��o/�DSSs�;����D�����ӳ<��RF�;/���O�8��61����%s���AQe�f�`}������e6.]i� o���c$��é>��2����+����J�����3���I�ño���kG�V��5$��uA���D��=T���b���)0o�y����Ė)�B�y��k�'���S=�����;<�5!����z��'=[,3Չn������i�S�|�����h� >���~a�~�]>'�H������������#�`��1x�pk�c�$"�/��D���D3��C�cK ���a,J1/E�X��QmPl�Q QvK�DER�	�Rȸ���5-Ў��b���=s>�sd�!~����#,��"��k-ѿu i�D x֛4����`ɖ�ݖ뎄�O&)<�㪛���S���(��5����hŖ1s���(����A���1��p'$[m�2=g8RɑB�o,���DC�ͥDF�O�E#��࠶�퉔�f�i�5�"p��k��Wȶ6��唓�Ih�:��҄b�����!�V�|���������j>:oY�3�����L��;���%��sB���d�#\���]��k�ۙa�0�N����RǻA@,���k\#b�-�@�^+39��;����(|�G�(���`n������կ�ݓ���^���6�_1볳��'K']���ܐ"��4�� M��������V���Xq4j[҉q^���,>d�fvo6yŮ�U�Ӌ+��܏�n(4)����d{ @jV���r��n�Q��2�uE2j��U0��ʗs�T���%�|:�	QJ��,�3��m�P���Ī��S�A
w� D}�Os?�eơ@l:m������܂vv�CJ��Z�}5��d�NC��~F�\�ѳJ�;�\&?�N����oz�#�s���1���2׮���Z���J�!h_vg ����h��>~ {;_��}�B�p������YW���
c?˖�g��s�>�l����1Z�ŉ��A�$8{A䁲�eɕYc,��������Fb=���帐q#;���=��CJ�=N�ӝ!ƻ��,����:f6�U�H��n� ����}��~^���Dm�Gpp��uK����3����^	���ud�8��^�=��o�	q���&�����5��:h�Byw��1Ls�OM�h-�ܓ䕂���y#j�v�}VL|��[I*��:o
��v��	l���Rz�ߥ����PT�C��?�	���+r�I��������K<���^��5/��1��?Q�21���H�qOq��dϞ8�d*�B�(��z����:��f2:r�k>�k)ƌr��j�G
Z���A��� >��~⣻�Df��B�;�&�FD�	�1x,o���O\�	�a��>�EFeJǎ��ؑ��?��>�c���|3�J�w|��pM�zK��r�.�C���%a���a�鏧��ں������ �NH'Ƽ� c� vxZH�h���X��}.Y�#��Y����^�ΎC=���
}�[_KE�$(f�&dy��������#���*�qἔ���F�� |wb�V����@+#�.�N(��`��B��uEv�Ԏ �"5H��O	�S��M5^�ξ[g,�X6��;O5�	������:�1�(���<��Zz�x�,��d��E�!"R���_��2١�����w*��{�$���w��*�a����1>[�;��l�H�%��(��k+�˪h"݈˳E�ro�_���`�o|R?�Zm��ˡ�Q'6�D�;1x�d���_%����isi��̃;E�xy����n"��eͲ�6�}DV߷�ؤM�3�
Oԝ������h����}?�q�j7��k��q�@sRXݪu%]�)c6��RT�#��1��;��ͨ�����H�߁�(`����:�� ��\�dQ�}fh��B��#x\�i�M���c�;X��C	 U�K��asMc������0�p@5*7��(7���wJ�`�������6���X���ԝ���.�@�� .�:��h##f�$�rR��Ρ�xb��캋}��p�	5ۤ�%vˌo��v��p1|��X��1��f-s�@��I�s0I�?6������@z������="�Gַ�=��U��2T��܋9���ޘ��"YP�O��"��?�Q�:�l����e�x0�&R���j�#���&ߊ2�<7'�6�C.=�5�0��(%q �,_�V$o]�����hHË��?���a�$V�;����3|�
�tK[5[��o3�i���<μ�����+r'�u��g���A���Zf��ۘ��[w|���wYO#$���?���T��~��F%�kp����~�jS��$�j���q7�x���=J�S[-�j<�5p��&Q�,��g ������q�\ �l���� �~1�$W�2W��ƚJ��	ς�$8 fo���a�ɿ���=��~U��$��Z֐0��"((�q��z|	hf *�䕚T���FSOy�q��n�cX�i/TR^%��
������Y��H^D�:K6����<>���Ol��N���t�*V�,�i^�dM����W��+���Y��d����ެ������d!��WYf�D����aq�M�P��ra$�ᵄ�Q#o����wG�]�G���J���A�D��;o����;���r���t6Ci1ȍB=%z�H��&�P�[ɑ(�P�w9��9���%�i�����"g�@���<�ɕ�3w[C2>������`c��'Id8�mZwVCh��l�S]��忰<��.~��	>v��P=�I��ѯWy�Q�����F�Pt�B���>�X����a8�r��1" ��gÙ
)��u��M�gY_Yq��z����h=��1���pp�h�2����\ `%k �����xF�V�*"{�V �
6Z(�*Y����2���m6Ɉ��N���V��Pr��ĳ ����\�	�Us�X_+x�S@�ò'c��8����`�T1G�u�%\��+���k��{��7�M��0"�M����g=*���)��Ӂb�=EA���R�ŝ��;�b9��
_v�\?�w��Naa���D�Q@�V��$k@�G�a�j���u���tI�/˽&7S�\�ͿL*����*�>м��J*���ٽj��=�V��SG,�:�QU���J@�sZa\�Ж���1��'!ٗ�r��� �5bp+���n�sj�ِa]G�be�}y?�eV�`۔1ǰ��I��ctV�Ч52��M� �M�j�B������*w���ǩ�n[m��>���zϸ�� �>�RcF	���[87cPZ1G��ja���Z�b�0�-������JE��j�,�zu�b߁ƕ�s���-z'0P���4jm���_`%��(-�ܳ���^�i���*���y�Y��Ϗ4bx��l�F|��7r��Y�	S+IN�8��JnS��3hHn@z�a��������gy�2�T	Z �<�V�s����^�R?0�$ދ�U��K�y�c��[�a�ڹ�o��6�J�m>�GY�U����)q���v�(�2r����L���
���'I��4���	�av��j����U��oF��ד�%��"�j
�Z���)�#�"=�8��8= �c���ě�6�`�M�@ZH�Ћ����č�]�4��]��r�\�[��UO1�f�=i,����_@0�o*F+�����&�4z�bL�_��8��
�e�����Д�vE�]ֶ��1�'sv�"Χ\^�cx��O�,�c�������,7p]�=�CaF�s�ݢ��xpw��!l�HU�1���{4+koߠ� �h�dM�˄>�k��@�~뛛���T�-@��.ٺá��w���ſ@�pJ���2�>3)iD��ઋ�E�&�'/m���oǍ���3����1�����H�#B�Y�
��Ҷɞ>h�
�?w�sI"�����k����o�����D;U/�rx�� �#FP�d�� ��>O]�d����l�4c�s��6���;���s��,x1�`bG���?c[����E:fͤ�ߛ��@���� �@�EIV��sY������z T�*a������P{ж���_���gʡdl���R��3�����2�N!���<�Hő����#*��Q?��Dc�چ�g�����/8��J?@<�8C�����fG/�}3�N"6���$�R�AK�1����)�;#Cb:���W�RRT�g�ygq,e�Sf0������EaR����J|��J��t/��ޟ�р�~�v��3�8m���C�.��T���!`4����fibn M�wϤ\c)�kao�[���b�	x���P	1y�#�\V¿�I�v��(�l^�v��=��� g��o����T6.����j/&��o�/�6�(z��%��6�I���_�a"d��
���#�{��H�)�ճ�v�4x
�_�- x`m%:���"��!)�\1�Ht��=�oѼ������E�k\�(
%p�\�Z'��J�8rg�� ��ˊ�C[J��?'iTV���+;�ޞ>s�[\�d���c�%�RM����Z�(���t�p��7P�q{_��7�Ȃ5P�]끩��JY�Q��PJ�(�'���P�o(�ڲ��;m.�ca���<FE���zY��d���o*�cEH��`V���Qg��+���ݛ 楨� ��F�<1K��<�xF�f��7Xq�Ad5��ٞh^���T���v�a.vb��P:nQ�i�5�!��b~�����17T_������͛�r����n�� wk-���y����Tx�m���W��0���	&9o	�N���7n�
��a&�l8ї�w��u�A�(&5U5+�������oB�t��=�wɗ��:S�5� b���&��DU�Js�Pf��q%� �'��̆my����h��ܰx��r���Gg��x!D���ާ�w�jIv�S�	tnQ�R!޻ý~��[�^͙4���	�=D R��0Lό"�(k�OMl!Sxs,�L�V�@F����]���͑�+���ݚ�67�y���\��F!�Ly�0�֘.~���K[xYӟ����]�iePY?��u���A88��h_f$��fa`���,�4n�\]Hy�o�v̲��DM$�"�i�ٷgo��0�ȓ�z�&�A�ĥ#4;%���?56`e%Q��2GI֟���7���Cp���Lg�^���b�<S&ߠx���E)��?�a On�o�`J�q��n���#T[��c�!��l}Rv�Ě��`�8��_��M��k�+/�$�Nj_��L��`I��K���A�+B7[��CT
{P� ��X�@)�"�:Q
!8?0�(+췿SЇ��!B�$Q[�M �e
���v�V��:�3>�]��!f
ʆHb��"��^��v����g=�=�_=�{�����Db�o�:�jvL %K�8�OA�`-�����&��˒O���゘9Z�0�n|3mE~��*Z��x C��L��G&fu�sǰJ|�@�U��ؖlo#������\d4k���Y@C ���f�ґ:ٟP���OVF�t��y"!��/�y#I�� aCٕ�n�uH���`ap�n�(5�|5�{�'SX&��5ݎ������Uh3.�/����pao/釁D(\�J�iW����`
�Dg�y���t��k�t�xKq�4��-�v�̑�{tՀ�f=�=`������U\[~i�6�gf�����PoMcLb�^�������ؓE����lV�Y�ۛ�
�����3�r����?'%��z�Z���h[�0���1Vj��q�ux���aaٍ��!3�	w�5��4 ܧ�w�i�?^�^a�]���[;��[R���,��j͛�n&&�|����K�P���2���tFmz�V��8ߪ�^�V�/���J�S�t���5���(]����<*��b�h��NNQV��	P�1�h	y�\dA��W�_Z]e��1��j�G��o�yH#��1d�2��
ZC�؊��3���ٜ�X�hݨ?[W���Ji����!�+(�t���f�ϲj��R>����ۻ��=��ө��U���d�v"oΊ~�5���-��A����G�=v�>Tq	��t�5�LM(�_[F�>c�(����l T�;�A
/*�+
Q�Ј$���tt�����{i��p捴�^�t|_��4_�l�2�65�iB�'�P��_��6�#��A#��,_�b���UH���{q{ ���_�:T��+���?U�L5N���.��G��>Q�m�G�ۛ&~��õ,O5�E�q[�tԈ4.щ�����g�=HLW��*�Ǔ(�z����V�/��͈��@���a�@��,�xrY����p�.�e+�AV�����_�ג��J��A�f�R��xg^b����f��>�-96�%Hn�%��{̣�=�v�~�ƺ#g*3�������}���as�Q��Gw0��nI�ooKG��E�k-�����Z�a;�M�)� ��h����7���K��G�C4��kЪ��j�g���0
�|b��a·�?����q˪#|q�n��"��j4�q�K#��^I��J/���O�~�� �4k�=4���n��_d`��PXn��tP�7rvo��g����&�X���V�yO'E4���4�}Rtl�T��*I�-na�Ф�`��`�>�y7:,o�K$OT���" 6-��TXY������
h��D��.�]��R-�7$dJ^��Q�*4aV#�-ٗ��n@�ݝe׊� ���:���W�u/�\nGR6�e��O�K�hMIK��v�r��ϑi���`�u�)�)=Gâ3��0�o̳�����FM>����UiSCL��|�4���i���O�b�Y�a֒���,_i4q Y��XAC���,!�n�c�q4��7�7����T�GTаz6':	�Y3Ȍ^@�Y"���C��I�K���q�c^�L �f@��3���d�R]�������XA�m��|X�<����?S��} �5KL�Ȉୣ"�8�2ձ�b}��p���@��9ī�Y��	G�ǉmC ����J�Dk���&ER�Q"%�vu��ח�z܍��3؉0���k�,ra�n�f��5e"�!�N\+�~�(_Gi��EY� �6��� H^�����hKX�I�v$jS�� ���^�v~�x�u+��`�:�Z0����>;v5Z~o�}R���6��N���;����	�Aײ��+�JrZ�c�J}xĄ�2���ky��t%�Ms	2��u���OOcW!*7#^�m-�|���]i���?�����v_˚ˊ��rG��r�AK���7X��fq\E	�.r��O�r��}p�9�S�R��[�7�l��2��D:"q$kD��}� dO�1�;��[���|p�t�{�>]��b.���MW�?��@�O�	�,?G!��ta��Ҭ�]�А4A;��a`Ps��#��K2���YA�u_Q�ts&z:����1�� SɃoƵ������I�ƍE��qZ˶Eu�>���Ҳ��{:��v���4F�Gf��\Җw�~���L� ar ���h��`^���I�܊Nm�x-�IEe��h	qK�ܕx� �����'���;�g�=�8�af�3e��wj��&A��Q�K�w�yQ��7&��ڪ��MS?@��(�JV)�DWj��l�c��^:�9�W���A|S}�W����.�lk�vzΏ���������_�]�D\s8�[���v��}��h�eUc��
��bℱB�3e�'L���/����4)�b�6,K�0b��Q�{��U�k��idFV31�fF�X��A�!.��T 	�Cl�ңF��S�['�<���d��LY�tҜc+׊q[�bO��;٢C��ZP��^�{�D��k��@��v�t�*s��q��	V��>�(���L�Ea1�yf�Ca�=B���(�UD'B�̛-������3�v��J����␬�_�H{�~?)-��}��KoЁ���f���"Tfњ��pG��It�m-'B�GLݸ]�Pۊ��8g�tWv��'�У��y B�_uMHM���Y@Q[?3VJ�Wk8$	��LœT��,�]�#i/���t_�-���as�_�x�Q��Y���g��v�Ѩ>��3���L�w�8Ix�������Ѷ���� _���A��A�[��S-=���G~rV�Ҕ�� ����҂j��t��o�M*����6ʉʌ��Q��J 4�ؠx�'dNѠ�	����R6��4��L���u�����D�r=R�$oWhD8�^���PXYƴp�d@��Qg���r��Է-�*�8����m�^Y]
0S��hʷ��r:��ҭ�E�1���o@�b�BL�d�z\��iW���)˓$WIJy���h ��,VD{^W�0^q%����ȔXF���۸{�_V��O�!��T��
9R8&���.�q���as��h]���x̦6����{p�R���]_��
��`��mʃ�&o�XѢ�/{����JܒrL�=��6��z�
�w�I��&|p8Wpϕ����C)J#�Dr�c}0
W� OW �+���2>��`1h��q�LԿ�T�.��t4J��9�X��Ƭ����P��|�)y�.��Rb6j��A����(1N���ƭ��rS�����H��r������O$Xܶ�N��/`'~���Y|�4�ȘH&�=| tKm7��ɢh��?�4�	T"ruQ&��mu��e�<WՔ���&*mvE��g� @O�o��E��v@[��89W/@z�Ł��+�σ�+/D&��#�V}���#@�_�Z�z����*W��*�P�_��Yzw���E�t�]�S.�ޙ�!k��^VfLx�Ͳ�ֵ";�G��@�ϐ����=�M�����9��V����0�Է�,�`�!��%��*��$���Z�I�e'[|��;P:�?7�oE!��@����_��ں��Z�w�����6��R�ʎ�k�Ň=2��Xޏ�B$e��j�Ä�^/����90�Kv���D�
��L�N�l ���� n5	���ʹK�G��iE������a�I��S�~a&�X���:��˖ق@
�,i�F���:�\�x�Ͼn�&�2�F�vպAl�x�Y�].W��m�V3/�[+���b���]���W%��@�?9��q5��>uH�z�|�C��]]�o���Lg��a��y���=��>B�`jH'�?�PNN�N;=��C?H��U�vǨP,|N�P��,��@-���[����|f�	М�Ԥh���ˀA�.��������d(7&�y���X����4���}�Z����	3g�Z�x�du� ������X���4��K�.sxL��%ԯ�bn~p����{vs���ȓ���5Q;�2�'VdB�x�k��sE*���p|� �"�1J�j_�]�2b�Qn��T�ԑ��]?�_���u0����4���<�UT��s��ԙ�3����"�B| <����'V[c���B�K��r��M��6482խ !�P.*�Λ9�"R6Y�x,�������dpg�e�1V'8��x����$�|O��B�u1v|��f���������,���䩩�7�.D# $l��{�I�F�A�
��d+��!v����b��I�'s���?p�����{�D�CjI���e�z�3�6r�}�JҶ������bt�WH�1�����Ծ��6��V!�9�(ik̘{�c���ZA�d���f31�˂ˆ��T����Hu��`q�1��.���H�,h�h�XIϣQ�p?d�)�'��4��O�j�}�뿴Y���Gǵ ]#S���T{̑��S��K��&;��iv�6��T̮��H�W���6�������;Kȶ�;��4"��:��L#��"�����ήF�
,��h�t�	�[ǒ_�v�[���s��c_c�
F�\[A���[�!�3/?d�ݗN��5�N�f<,z����Уn�������w\�+�I���|��֛b_ƭ]ZVf2	�����p���	:w@1�B��������Tu��,�/�JDv9�*!���Rٯǧ�t���}och���NM�.}�.@� ���]��I�zz�.��~Xcm'`�G���;ϫ����l����A���ݟ�P���l���%�ɹ|�6��FU^�*�r�X�ـ�B��:�x��?;*��%81�C��S� ����f9�����#�z{�(�m�����2�+*��! mL$Ѳ��Akݪ�EEYea'�� �����	֨6Y?=��G"pF��׋>���.T�ê�׎.��?7>�� -��o��%��@/B�1��\b���v�j)\�L��}v�_v��^��	y�,*:�G��c���-�9OA��s�8���Z����^�Ҁ�l���`k �Qm�'�񦬶��o�f
��������p�B��o���Xs�k��(�e�����f�#=�Ze����ɻ���~SXw0C�w^��B'�#�Jq���b/4s1����H�^�q�Vc���F�E�a�W� 9�������+h~���R({�M���V1�|�z�恽�>` �]�D!��*�>̉(0���N LAҢ�H5>�1�zOb���Ou�\���i�yiQv�A
�)d��2�K�+0vэ�hz0���*���7a��FN�.�b"ɥ'�[Nx�+n��f��\�o�p@�`��7�@���\�^�/��5�^X�{�_Ya
���s�n�8��*'�KkPb��KJ��Ng	����H0��AK��4v�VJ�KΥ�B.u`>O}��?��O��\a0׳夌��Y�������wQ6:{�qv�$b��r�x0�����*3X�M��h�J��V�܅��u	�O*�x��?��S��:�X���e|��{?b�84�٨���3�#Y��!�t����c���+:q��^�%����a>���xߝA73:吏r�x���@��UD�]�A��$^;�&���H8���х�؄`���`?9!�c�X
���t�����;�;�7�(Iw��&�]��,V3è`FC]���m� #�X�+��5Be60!5�͖ک����S�T���ا���FZ��r��Ɣ�;��AOFvzF`%xLI4(��GE��D�>�#��ڎ7��JxB�&���_ˣ�dYlm9B`Ÿ�Mb�'��n�X��N����}��]���|e�T�+l;c8���?m�� a�V�G�G�α�K-K=,ً����'	� ��*
y���N�P\��)�`���->y��ܥ	�O�|8~
���JZ���g����.)R'�m)���&�&l.4Zk[TI	��>��0$���'-'����疺ڛQ�U�~}D���> �8:��[��"������xm"A*�l����-��WT��l�J��b-��Z��ȝ�
���u��K��J���0��+����n:d�|�������7�B���훾�Bim���_E��ԧM����з��s��p-E���>�z!�y��4#%_摠��x�4;(��R��T*���mi�1��������|��K�d�ȟ�Cj�W�	�KI�`Y�s�W鯉�L <Y�_�l/�HJ�Z������]�dU<\�Qq���.;w�زy�U�MG(�?��ox�qꎔ��H��#��O�DtQ�����1X���G��T'�\H�"J��k`Yl,��Hu �rW�?�xl�_f*�qڔN������v"�fM���J^��Ɵ�r�˟B�0��G��f��_����$�ꨐz��愐&O��\>�E/*<.D��hS�T�X{�C������ ')w���e$PZ�Ж���s40#�0U~Jw�k��~Yx�(�B&���e"\<��d6��� "}X��FI����!����.ì`$���_�C@��s��:v?m+��Z=Y����:��A�Ā���=3vd�u���.�R�U�솆�͆��tM�>��>]t�K�����d��Ð;�>��np��}w4�Y�U!QϠ/:
�m�Qf�lK����:���J��=42�݌��1(Ca�N��]�����C'����� f��h4r�f\�E}���W#x��������ߙ��K��"p�s����qn~;�U����6?��R�b��0fl��"�(
p�?5��8�����_�eҰ����
���1�L�c�B.��uKȵ��ޤ=�Zn�!K��1{�>��͖�������8�筛M]6��|K�D�-Us3H��3��:�A�e ��`� �\5�"[�>�~����&�B����,��R����8�4��&I�3����kmE��YO6�����?��ƣ�F��WL��>|g�ߕ���$��ø�������W�_R��-"�����T��J�*yGj�u:)���nJ���+�]Z��W�Orؕgy.�I�5�E[��&r��V�����3��_���$b�z����= .ے���_�n<g	(�������
�}M�آ���J��C~Fp��D���o�c�o��1-J αE��4׀���}��	����A��P�or�8w7�}l&��iIZ�*�P�1La1����͆��E��!3�t���S_��Vb��T1�k�n�g�n
���䶾י._j��2�'͇t֞Qcj�;�Q��<�%r��eY�w�e�������]��y��:���\���>X��m)���p;�C}u��#��ׯ��d!��2a��e��
cP:�:�2�3߮<�,��jUƎ��s�<i��'�t��+[`��lV�R�C�M�mnD��k3D�%�D���]�o���T6��J�Đ��S�KB�p��\DH?�4�6�KKg�6'#��5S!��j�����wY�)�oU-o�*䇺����`��_Sޟk�w��{[z��������Pwb��*3Y����gy&��zrW��*�����2w`Q��z:+�|+X��Y��\ �Tu�[�I2��'b9�o9���Kࡀ�������VQqy����oS��(~.=G9eY��Bh���&���1�.30X9����/:���I����0��F���h�����50m���5>�~�{l=T\�����T"I$zHnK�t�ڿY�(�"�W�ÁA��B .fdm��~R�QIs�g���U�a�5�������I�e�MR�@�46� �Z&�6�Ԅ	a�)ã�^|��
s�y=�h�ϙ�Rzu=�+K�f�
9x�9P��L\W��N\��1a����;�V����x=*@������I��Fޔ�c]yP�9EwM�h � �+�x�0� ׼�h����i/�dK�SY��Et��P�\2+M��#p�$C��P�Gv�Z���?��v�n�������g}�_*���-��L&��N���'X�&��gD��-�Dp�Rl�c�lMŦ(���%��N�{pZ�A^zi��I���3�?ul2ޙ��vh�7^������ʕ湸�'��
L�=�\��k���^d|�v�F �Z�l��7cgisWzalv�QG���Y?�d�b���!�x� ㋳��xa��'����C �7�Rao�2��w#��J��I�0 ��&��KvY����������/}�Y�+��1"F'�XAQc4�(�t�*��W�/ *��� �Ք������Z��{�owIx�Y���giK�|_�zub ��x`-�!�ߋ�bC�`����~�(�F4 ��~��#��ܜ�^�q}��y6�H�b�TD!OփE	�"�����׌=��ǢGmbt��jL�]�V!Q�����cg�O����P�n���ꡑlt��ヺxO�ԍ_oU�VXRb��v�#�c�EY��y;��q�K�2\�_�q�_�w���G��%��G��E���_��9X"6�Z��D>7�Hڈ�� �O$�y�Ki���������V�bZ�L��ƙ?bM#���!qs~�/�J���ݞ��^��$�!�ŕˁu�<�N�
�	]��>=��*%i��o
9��1���"
�|�氬7)���y�
���źhw��TΟ8�2���?���>��� ���,\� �^a����h#M،�������A^LUjO�/a4�B���Ҝ�dm��Y$<U�	�b#gW�=�[�z��@W7���ة]K`�y�Z"�sz�
�e�m<{Z�4��o���-�i��+-4�*�g$_f�o���1�~�)��Y��1���}[0����a�'��ժږR �A����:�YF��Gp̝��$@�:]e�T�z9 Z9[���R�Ȃ�?d��b��"o�8x�����)#���d�\o��N�?� J��h匝���F0��{��R(9��G��ua�LZ.�R>l��樣��<���%T��|�����h�v����?���5#�o�s;`I�Ey4����y.{�x�;�.�5J�����vn���	~�d���i,�P؀��,�%W������}�	
�~�	��߉h�<��e����`#�Ͳ�^�L�V��1c�*V�I��,� ��G�a�P��=����Ȗ�}`�+U�R�&]�.�����V�+�>��Ę��A��~5v�� �q�.���������5f��6R-��D�i	��v���1 ���D��y����ߞ�2�.*���n
�`�Z7�=ƞX�cd�pW����΃���/�����sւ�j�&\�s51�z	��WER/f�m����U��i:�����%N����NH�(�t5��AD'4�l����B3�v�2�S�$����o��Y�嫯�MSJ�  `"z�]j�a�(r�uU��Ģ�vb,	|�(�B-M�@�a��ΰ�	K	I�)T��,g�����$MP�Ud]�#2����}=n�'����`{�J�Lu�.��DLk���a8'�)�c��%ѼE�ls��E�4`��q[�f���}%3�9��5M�ޮ?G�%��Up}x���	T����������Ƿ[ajMy��$�B�t�6�P��I-�c;G������p�m�n�T��t5��ytycB�a��U%��?��Xb�}�6vd02�I��{9��v1`�UHY���dS���ؑd��p?��hV���{"`n�*�3w�~{�w1���m�:9����'E3�>�ն/�tm��:p�=���DږتN@��b��Y��:���[��j����إ�_/��kr	r5A�Xrsٍ��*��cF���j&ٶ�����Z��*e��~2��=R^^	<wt���A�x�p�3��w{�ӫ:��e��7E�S��GD��t��^���)��
�8ܮ�E	��� ,0��A��)|D�M�ոC�|�ez�CQ��<����䭅��J��@�Wm��ͣ2�񫲌)�n�F�c�~#FI1�]P��44����p��{j-���A��J��+�]���EVjO�$��8n��r�D�}����0(䐮����ѲC'��y�k��jv�F��>RF�׿`�D5�4P�� �3��h.�G^e��4fY�Ń��m�P���
�c�W��Ɖ��� pݮ�ع����D����ܞ�YZ15�{B�h��)�P�ҥ<�A�}g� �FZ�/&�M8-�4kS*[j��3��V�o������1���O֢`�ٟv����m�F7����q6����pb�p&*J���Ǳ2��Q��X�Vf0��%���	���6x�Ó��)&t����U���ЬD�.��JA�>�Ũ
�훮�kp����6�u�k蝪��U�_�d�yL���.�E
C��E�F��d�ג^7�͎:��Xꘃ�<�Ћ��)��L�ـqB�<�@T϶�������Cm��:ل}��X� ��/����G�5�]W˃ƹӌ�e��Y�V���P������sb������w�ۃ)3����G:V�8���봋�p 
>JU���&+)r�5*�ۂGQZE��ϛ>A�Z"�o}>�rV�K&Gs64�Â��@(���o����u�t����>D�m�16���~�d��L'T�1͆+gn0�9��v���F�����X�ԇ�A'�)1X�M��k4�ff��۸0SW}��Y�o��qC���cCJ�wOVbc�ZP4TiG�.���c����MSl,��5�3����F�x�Y<�'��ЭO¸I[���:��0E5+kJ�b��Z�:Z)���ֈ���5�Є�1�Ӊ���)�����9�ۯc��m{`�1Jv�^!}�f�f2^I��sy>g;fI����W䊗!ѠĽb�'܅#`�.��]��
�F�-dV܇�I�c���|7�wl4��3)�����!��|_��zn��� ��}3�bp��\��v���^'x�>�u@ �����Od$��D��	�.@�X�����"�݈�v�'��5�ƝZUHc�r/I��s�d��-�˙������yT�͒[��[E�B�P�%/�)�߰��=�	���q�]��O�� �I��e�BG�~��5�*�l�M2�C��H��Z^"�3ښ�	 6���;搆�j�S^ǆ�l�����5b��*?g��3�>�UT�p�%��F=Y6��*'���dZ��7.츍�U��6K�y��o�P0��KQ}	�4��^�y4H-���
�A:���r�?�?������K��)N�w�	�`Q�ͣ��y���=�)<r
gsdg�������w��#��_��Fv�ɭ'%���C�♹<��Q=ڭ�c�b��vpf�N�v��*�T@���n�w]M�2}�+h���sO��p >"���ۍ�22����Po�{d�kK�ƴ_)R�]ӫ�ZT;P/_�W2�&��#�\z��C'�efcp�������x]�o����?1S�r;���S@���k�T9S���?���I+�m��&t����|ׯ�cO�i�a��z�;(ǵO�^�����Y����r"IN�z������uF���
&"�p���r(i�����2J{"��i.m���N}3lz��Q�V�V�Ro��Gf��r���;^:h�3��>)W�2%_՘}]�i�J�ȇ	���M\��w�S���ɀ�z����ti�~���8����"�d�.�SږNse;6��?�� ,��#�{�!��xP���nFG$���u����w�+��9�m�k'�}�=�4vn�:K��$aR�6�Խ�E?����2;TNL�4�J���sL�	�� ���sf��#�ԢEꒂ�/�|�)x�+.[�Q�)>�/�4����E.5\��nL��jk��h]��ۃ�����o������ʟg�n���e!�ͽ~���xi�̶⣊����[��z��U߹�[Sΰr�g��K�7LY�D����I>��S�&C,([c\����T��o�����O}�Dy���Ղ>ۖ©q �*�8(�����6+��^Hn�i�3�y���t��5g��M&�!o��{~ٽ��/�#	��(�F��6Ib݅��9�NU��9A^�&�ߵJ�6����~2@˥�8=<Iw�{�CG�g
6@=�V׃r�����&+�k�ő��G\������".Ѥ��eg-��x�?����O)�1�7�Ԇ�/jL�w]�M�ͧ�9K��i��oE
� �����6&� ��Cz�UO �N�{Mʸ�)!�L7$DKӢ1��q��%,�a2_���tZ�^1�%�eA�{�K��\d�T�}Lx{A�<��d�b��֖�Wjd��|]-��62m�.��^g�J�h����iMP$W?,#��xZ��f�����j��� ,�Q��5&2�#8Qݠ�y��'w(�q�����9iJ�,�����0��]3�z�O��\���ޛ��G�Ө���Zi�-Mj�A`܇��eD0�N��&�c�i#&.S��{������h���Į;v!�
+�ͯ$Y8��=�"������)_��n�.�ͅ2�y����v�̛WkU��:6=�	�1B�>1&�'$E$
�����:>������Mӵ��6euV�q[�u���&�_<u��Eb�*Il��5�΅�J��ؗ��uM��.��1�sBA�Z[4���	K�Cw�&Y��6����Mޟ���Atʚ�Vy3/�c�6[�aWS��|�ဃ!�@ ;,��Q�7yUB�f$��Y���"��䂲�8-�5�{�9�בFo����褧5�T�o�XxjN4�לj-<��#���:C���i�a+���{�r�$�3��&_5�����õ+}��Z�RF�k�I�����eVw�H�R?vc���Bl�Pd������3��/��sq�����#TI,������IwF$��PG �/��h���W���/{ӯ��������]"���f�af<�C��~�'�n[�QN��7�B�j�5g��e	��~���ġCL�-���{�}C��o;����pnS!N/��r�^fUT��TM�oR爱��+�@s>֠�tq�ڜ�����4�6<�J�e]� �¸�ls-�(��]�%�1K�<�x�%*W��:0��l���[�P��?����q���z�`�$��7s<�_����CZ���Z�E�F��Pp@~{��4���o��:�䍛���l#�R6<:�b�">7ƽ�f���䄥R�,�aW�2����-Y��_�������i=�b8+K�Q��R�����{��ӌW���N�I;�:X4r8x.J,&��ۆ�8�j�RI���&WX�:�����ɥ���.��Ll�BI�3��(=D΀�G�L�t�t?����JF19O�q6�H�Wa徨C��Ni�]��ӳ _rT(V������O���s�&P�S��YJ+�1� ����W����drRA�c��+p�����'
K��y~�+�Q{%6gE�fi�[�5c��Q�]D�^�λ�Iq.�#	����p�Xaikŧ�7�l���%8QQ�8F��F3>�`@�^�̡w�br_t[� �j'��p�)_r�씰��U�,T-AT�}(����o�(Utl�zL�hp�8CC>�x�??D�=���K��VJ����_�#�黁���l�7K&���<���Ӎ�_���۱. T�&L��ybft���aK�_7)��3�s�c*��F���g���], ��7j����^���]}��3�
����̙���И�E)R\��U�זK	�t�{�Ɏ��hPs��@S`������u��&��p�ϥM�Adf��F�H2�!d��5�%߭j�ꪮ(��'m�<䚗ӧ�1������-�
d^��2����o���*����^8%;Ѽ����h�@���f����F�*�D�ը�a�ڮ�b�p�]�cXn3�98<�~0$	�x��b���R��k�h��3.^�]�b�G�U���M�O���12-j�Q_+�\��)<L]>��?��:�J&1/U��V�Xqѯ��|/9g������eύ�y���sO������v�蕵@��(�ct�o�ǅ"~�1N~���*%�\��H�f;�0�K�h(L�\����9q�eB H�`$��	�9�f�a6���-�]� =�ӵ#��ɾ�<G�8��f=P�|�I̴�3��8
�c²)�Z�f�����N��Db�>�����dy�j��j~�w�?>"��6�)Gq �o�6N,M/ʂD; �3���l8;����,�+\���O��a���U/J��`���RI��E�5^�f�C�JD=�6H�� A�`T��O�9[����r�ٹ##g�꧷?��?"��elI25�̙���������� [$L�y%���A��ߺ������k�x�"�IL�	��W��CY��ӟ�h�Z"bXQv���c>��l���zQ�1;B���+/�Գ��ʨz���5S#5>�IН�x뎩rc����3%Z&�*�;Q��S\�嶖�E����X��_	���}�IdC�@�t�x؟-9�2�O5�}r�=n�-vG��t� ��� ���E����V4_�4����>QW�5��ke;I�])�Ι�İ�8�F�5u]�h3Ƅ�Nd�8�D�c��+��}I���g�F�0��&c�k�S��++�>�����ֱO���V�f���y�K<�wk��@�,}��3ڊ��`����\�,r*�C7>���h��(�BI}�����N�{2gh���r��WX
�~�����i�t?%������d����z�Bj�M�3������K��
)�n&\��9ag����J����+J��9n�#�ݯ��H8�ۘcd�#Y��
���$��Nt
�Q���Y>s��2����z UtjHː0K���j{�ie�Oŗ�a�oĦ�J��u�y�$o^�5�3gV� Z	��,Ч<W�&�(CJc_$�p��\���J ��
��
�ʧ[e���A�*�%a��(�m���F]o���z}-I��*�>���\��G�^;��s�� (dsb��M4R)p�)@̡�%K�+_���`ط4�� +:.���:<�A���o�o�T�۽�#pF�\q}	p��}Pw���VS�V���U�n����VL�E��{��G)X���4쾕\�@>����ndn��s�N�ԟ�=��%�z���;��Ga��� q����m����=NjB���3dCH4�g��j�'2\�Ml�f��J��93��n;���(E�Z����`���S��cQ��ãZ��v����v���4xxZWC��n{b�D�l�M[��=��1+�ې5� �󚐘��~K�����	�9���������
kn�s�4;��jc�q�e���9�r⺯�r����vkd1s᫿�=ZB��)&���c3r���נzq������5�^�X���0-��j^�c0�/���=���n�e{�+]�I��.�]�vB���7@����#L!\�<���oH�X�'�A��Gf��(78�%Sb(�<�wm8�r�x���`�ѿtׇ ֥`��(�p���e䏴����V���H;7��ָⶦVܪ��b�X��l�	3������]A�@N �"���^�%�}.�����ڬ��\�PC �f�S��Ke��E�X&���7#ȗY�G��@=қ���4�����7Ub5r8�uY�13dz��P�V9GT[L��7�K� ـN�8�Z�.u�%� �}X3��s��݅�kH��5x^T�nI���?����Dt,������ͦ��Soץ�g��o�Nܺؿ�}N�,�y��P��%8�fa�:"��y�N��0� ��L�����ĺ�ȅ�:�2�~�xU��w�uƠN��RG�������sy���l��ܕ��|ܐ
��HɾZ��"�Y���+��I�J�.ؿY��[;��j͌���"l1P]c�b�o��d�/ɀ��EfԆW��+w����+鋦����3����_רڮ�-ɭ��<���<�[��TAP����{a���Y�pA�s��������$�'5$�
�ǃ�t�)�����z���7�oߌ��U�z[��\��*?WIMu�NЅ�����x���7��Ey`�v���:����6���kr0��P�5`קz,�*>(
~Y�3�L�Z�M#d�W�s�mc3�jH�M�o��5=�g7��b����gլT����2��?�S`��&��$��	�����4wS>	ƴ�Q1=�S�=@~P�2蚉�u9�Y	���s��<���Ջ�qt4�9Y�����qn�][�YB2��{5��v6��v��P�i��7�Z��BO������S�Էe���]����`��q̭_���-�O�4�9	����&���B\��|L�`�̝���U19y!�� �`,B���/D���I�!��r΂h[���M�������/��8a����d�h R|貧6V���H�H�=a�����]��.=ԤJa���	�K)*�W��B�H(���L�8?�/;�7��1��7��;��>\���>�6��Bp�b��\��Q�k_��E~���Z���j����O���A%zHf�~1.ǚJQ+��j���0L���_����m7�r̳յ))\@�yl�&Y��oS	Ś�;��v���%��'���8���kN�q�7�^m>�Da�;ZH�qx�?W%DpG�+��)�>=�F,y��!����⨜��W݄�ʶ���72Ʈ"&γ-v4��ː��N�!R;=͑���bmp�����^������9�d⠁��i��/8v'-�ŉ���/��۴�*�����7a��.?;��V�y�H�1�$��LТ���r:u[}�E&���8�x�N�c�eo�XQ�'��|h��cw̻�<%�֝ ;�l�e�u���2
��쁜+}�cʽ���н�ӏܚ+�ߠʫm٦oy�°� �/���kD�Sk�v��<?ѹ!5xM�a~���G��|��
�'��� ��r��D����,�99רzz�!|I�A@��α�q?@���L 5 �_�w,�����=�w� ��>��8�C)�
U�W�X�ц�{���m�͹N<Ԛ>����3��Tw�:��9>��a~�@v?q(\�4�W9�>�����$�-l�J+���8UT��"�Wh���=[v%�?�`b�ҡ[�A��؉�'���LI,K5oy�1�"��z�ln�޿�K����'�g������|�`X[w�s��2�ּc���	���v|�����.��36_�uI{�������辙6Σql�Q��(S_�l���E�B��Y%�+���x���S��li����B�PjM���xn[�]�:��Y�׍)mY×x+3�&%�/F|jD(��rצi�_ƙ�Q��q+_H��>8nW2�rL\�,HJ�b��]�F�c�^Ui��6�\�>��SǠ�@}:��f�^�V��@�^ں��X�5��A��%��|��S�����3�kr:� }[�b iw��|z�ic{�B9�ݻǌ��Q?�C� ��y	�+?�Ҁ2u��m8b�y�S���'!�d����T���|N1p��r��%��27mAE���Y�ٍ���������V�1���'�y�D������xZ󄜭�uF<`%*^�$��ewf�ڕ�+�@ ��s"
x{�6����z�)�u�hE�m��1P����E�O�PL:]���4I�	�	�d�@O�v��K�~1&D��v��J~p�%T�ο�b��m��h���~�[��n��ߤ��*
6�j�D=�/�V� �f݈����G�z�=�V
{5��J�NnkX�i�g�� .Y����`�ڈ;̢VO�g�K���%kn��C��;~a׎��HFZ|�zPLP��3oR�chBˌ�[�@k��2�5�'1f[���O^z�J�GlM���(�2Ѥ�y&� HơM�!#��u��y#���,�l�UA9h������EJ8��̓��;���快i�|<�9}׆��g�&��>��,#xT9J��G"���XA�dX:7��q��[t��;�G�n�9^�\Q�#U�84�z��0���j�D��aw,M�ћ0�������&2'�vN�\���E A��~�V�;sXM �Yω.)�T-V�JK6|�+����ǲyX�D��g~���&��>Ʒ0�9�߀ Љ��ٜl�Z�%��\�'��s�%$��T��jo��*�WQ ��ss�;�2UAW�|w�c@OO--�+�A/gX�[���hbL=�S9lW��p-K�:���-�ͭ� lK4.M���٥H3\
˵b��+���s"���c3�ZT�T��*\&bB',|^�_�%Lp�1����"P�&�2��F� J��u!�(BP>xċ��6��C%�ʣXa���H���!xŸm`��P�t�'M�?��n����o(W}����~�R=
�
o@�!X ��m���=�C\�˶I�(�ۣK��,�W1�tr�Sݟ��;p�ŕ.��2M�1D;]�q^i��nc{b3H*M|_��:�@�T��,�CFQk�6������B�-��AK]���)���p_�Y�;�}�_ %�t����n^m���&���\eG��ơ���	W�%J+��`�[]�g�e�%H��0��'n�^�櫱(� �e1	ޖ�޴�V��h��o��j�o��Jg�cR�r\��z�1��f��/ ������
M}CQl��Nc�v���ޑI�PQ��UR	��N��x+�,ֱ�>�'dt}��c�hx�T%�\{���1F�X������_y�%�D�����6�Ŭ��!m���E*T��~�J@S�xl���t 
����J2���;&|�])g�hiD��M ��:�e�[ĜR�,����"����=�.9E᱉����٢�9�.�9�����	�e��W0]�qh 	�5�24{є���Š!��Cq�DTl(L��ùU"����]�s�C���X>�5,��:F��F�r�W�lҶ��
��5�����{��<h(w�9�_�A�KqV�(I�����$��n|잸mx+"�x�S@�x��E�e��d�Z�i�����ֶ	� ������#q@?�����3�������G=a"豰�:��"�a|��A��	��zY�1YL1	 M��u]¨�(���а��U�P �xL��;ʌ'^�� a�ث �<��F��J�o�A��#%	�|
��u�����~Bg*��%��&���u�͑;�3A�e�yCb*�HN�ѱ�ᵓieGO7'�r�H��cq����,.q��w���l�TK�x���iޥ�B(Ur�?	�ǿ}�Z�/{�o+��/�A��,��\L:����G�a$L4VĦ >�(EL֘���N�D
K��:t�x{2��#b7����,?\�"b�� ��L"0`��ᢣ����������GO,4�<�g�hZ�s&�}����t�`h�]���J��bˣB�s����R����fv��"�"堧���a�ހf��|!L�|%$���/���P&� /���M� W�c�	`xyL|���/*�:��z��@�|�a`eI�K��M��U��۟�QP�\㨫��V�?:;ea��^�a�湟 � m��%���J����0�³�s�z�^�C�i�����/eI낭�i��"xw�$1G}�p.���qC����)����w��- �� ,��k�1� ���`��I�$L��������T4��
x#�q�����2��n=��������Y[	���I����w��z�j^!���HC�fۉü�=��#�*�:��7X��BЍŠ	� Lr<0ͤ��c�z�#����:��F^�����A
�z
s��f�ۖ��n!eKj)��i^){���O=�<"��*ݍ�5��ſ�>���eR���
��R�p���)G!/�n���m,�t��J����0������$����C��U��t7�����AD��f$�#6?���M�06���0+C�.�Zےsِ۷��H�۔�x_�����w�Pp^w�g���`zܐ�A��mv�V�K,�
��9��6X&˱��r9�E���C����w�s�<�r\tsUx�dh�
���d~%ױb����v���zb�L�=?�8�`��bn'_���X�f�t�Q]�b�� ~���߁o���]�K\��]Y Z��˕�����ē|��R[}��S/�����8�P:k�"Wў��ðu�@�<�{O�t��Y��8�yj���ل�!:�ݧBA�DՕ�'Y��a��k�H��k ��%8����Sox\��0T.V���W�e��"[l�0�>-8�O+cZ���}��=���<���^{�h��&'a����p<�=6ګm()`�wf_3,��Q��ܱ���UUa9 �z�Ii��H��~�҄S`�X�Tm�p����5 vψ,��4³�}>�|Y+tI1v�l~sʱV�|Jd��a�:����E�܊I��#��j2b�Kn��t��^:��2�c퀻F���)w]ǈ
�@�`Bd��f2��\u���F�WNՔ��n���*b��ƍސ(R�_2�=3�T���⢌p|8-�_A��I"ݧ*6!�n3,Ɉ`�v���޲l�Dn�".��3�q-ǅ�zw�������b��Om^���H�j�`�
5m���-N�Qn��X%�\dm���#�*.[Y��D!I��a
��wi"M-��[��k7�/`�'��%SLZ}`/�%>3��8���i5��c����R�N���]�������[An��Q�/�f�DX��Ѣ��Ա��ad\kD�)g�*X�p��5W�o��e�͵�g� ���F��Ĝ�5�lܔIw��҂��Q"6b/WA�U��*����!xΝ �4��4\,������*^f�~�"2�P.<��F���B��l^G����;���`�5&'��|ߘ�ۘ�A
W�	����z��Tg�ϧ��tY�I����(�K(�����>EXw?;�����{�u��M��K��a��طT���B�i@���[@���(�g�I�xV�'�܅�ӝ}���(5�ogӋ*F83�w�/Nϔ0�j�@��i����� 句���6anʎ���i��.�1�e�N0��p��gdC���.(��Z�lc}���x�"�V��yā�\}^Ց����k�4�݄��H�7Uxf�v��!s���z��	���a��l͑G�n��*���)
�Z��@�Vȑ�L�z���ED��e���]q�-ӾQ�x�J�xƺQ�l�	ת�� qOm�@�� ��!i,�}i���?6&MBO�980�����3_��5���A`͒����ߘ4�4����{�,O���w�*�5�PV�J����?l_)��ܸ=��.N����y��|��$&2JD�CK6�F�8��ѡE�ñL;`�����b����,�^Gv~�!f��O��!����Dʺ�J�\���x�R���p��sN��Dˊ^�X���['S'9B]&��EH*:$�V]���ɟ�/|�bq�Xp���Ny9%����և�nU���+�����}97��7��_a+�2��?�Ep�K���Ϛq+>�YA�������7+чt	^$�⛱7�hB�r�pj�9�ݗ�g��Q��� ���O⵮Tu�Y`�f�,,N�P�A�(���
^J��P	?�-l�c���9�l�u��5����_� �[$a�A�+����C�2�\!��Ty+�Sʈ��}��a��۴f��i�Nb�=5[��zs[�/<�?�Gn��2(�4ʸ2ۃ��`����l����~y�P!<*ԝZ�(k
F�B�?DmҔy:��b�ؙ7�^�2�O���;�C�p/f�I��X�yt��*�q���zS�k�y�>,qe��WEȴ�pAz��7~W��.��޻�{���,a��!�p�� � ��(/=Xt��r�������L?�O��ݗW�Cq$yVE7��s�ɭ߈�+2�O�2h�aZ�:�Fn�;2i a`g��ن0���6�~6��@iѴ}v������?'�椡�"��V ����+f��L�F�^=k�V;b�>c�/���#�MU4�|R���fu���kG*
	�M2�kn�E�I
p��El��M�A������;ye �	�W��;�i��sиб������f&7�иoPe�&��q3����[}jK�x�j~X��8�NX�B^/)[��6ޭ|��[4Ǹa[���2�b�w�ρ�s���Qc�&%���[5嗠����Z�xtUz�O�m� o,�������wNʜwSi[�}q�ڑ��ihK�"X����TP4^�lY�ה���"8�T}J+p�Q%y�6YMBU"6o�YP��ˠ�]�@w���N�٭}u�`���Ɨ��p�l߱E�x:�-�o��n���p{^g���!v�6�;J�Ej8�R�0+��S�lz(��y����תڴ��\�?���
��`���Tk/:q�EiS"*H�E8��vOvZ�_gO�w1w[�����l����#Գ��n�Ǥå����$b2����[��l���-��&��!%,�m�kAjq��͌(�n)%�X�6ɬK�!���A���א�gA����E G��[Y��	���1Mw4��<���jUp3x5��Z�w���K}���ph����O���X?�vA�(5�W������J�hDYk��n�	�Y�����i��J¥0�rK�݌Np�{��禺����ޤ����ųUs�j �����k�GP��nkF�;=�Lrar��B��mc�'���[��M̈aဩ�*�G�Ũ���f�P
�6Q�h�!�T�a��J'q�X��RCZ|t;ᢏ,q~eπ
5}k��u��\e��4�	G�5���if�|"DE6�5��SFv�c�Aa8��*<3�۹�J�����k�M��>�MV�x��2�Ӏ�*�����POm�K%�����yMs)욾�E^�7�ڸINڮa�Њٮ��^r��=�V�F��Õܯ9�!�
א���?��;�D*N�=1�L�+Ȍ�S�2~N~�(���$�y�22������c��8�}_iHd�$)�<���T�9Fq��D�k�Q�j��#��Gz�@(����컖����P��>��h�*���(��M~'�^D�x�K�n�p���R>{2\��M�gp�y�&�z�ٛ(�S��S�5>6��� iq���p�(R��dN�gmH��{���J"B�b4�,��G����gLQA/BY��8s���K\�K7F}��f`(�:�7�5��P��|�_�BU�r�j�W���J�]�E�>�Q�q�0M��Jm7���d�gy��X�A�*.P���� ���Eh��Z9���Z7���my�+w�B��[{Ӯ G�����4m��	�6WT�P��2�FxG,
�9�5P;!�H���9+�o�T(��b �ܾ���Z�����8�t����^O7�d�c=�pUn��P�R��4S�"��#`��k�=���Z��3���_8�hG�Bg���Ni�_���ѡ��SO��ߣ]�@�w�d�e��i�, �/�ac���seCO`hʔ(�j��	�v����O�qx�P�a,��Ѩ8LY����7���-��tZ��!5�':�W,�:��?6�n^��F��|ʥ?a���+۔��v�D�_Z���Z3��\��	�'��#:�!BIB���!л���]J���e�mt�B��/i�~H84����w��G�I�H2��W�_�]��.~��W�8�B�j|�e'���y��eVb<�b ���(e��ul�Æ_�0:[�W�p<�쑫X5)�}�)KJ!�ҵ�k����H�Hٹ��s�=�{M%kG\>�",���ҷ"FAH�ce��E���Xts?��SԴ��g�)��������J��IK�v4���J���o�"+�<�\��0^I�n�)-��V����`����@�����
b&u
M����Ѽ3k��i��S���,B\�=}�/�H%�������l4��=��R��;�w^*Z�� 5���xvi�-�P4n��e º6�:�m��TɊ��p�N3X:�IB��7		i��Gy�N�p��7�X)e�J�q�.1Q9\5�]��n���K�Aޗ��Ef_�5�-�ܡ�Ȁ��;��1}F.z/kb����^�j>PCj����WN�r�����O����Βa2RN!*.:����2�p3�8�<䬿8�}���~DA\ns 'Z���'N�7n4Sd��ԑ$���#��A���3<���@�~����Y���9��Sf��	�˷��DGr �$�����,hJ��%yx�wVy�y�R�� ���fѭuY ������'�4��R'l""4�+^���jE���,m���� [���H?���u�$�EX�M��׆�J����(���xD���̽�.�0�� �t��+�ԓH�hymd`������h2Xn�� �S0ĸ���U�&���Л1x_����F��+	�~��;VXJ4�����gO5��»Wq�9���Ӌ;��ē{���{X���"��y��%u���5���ϙ)6�;���!K��)�Y�����0����[������r�.�AM$�Ձ�x&ȗV��,��dO��#��{_���z�wD&��4�ջA����	����`D��G~���ΚXE�C��:R��"{�ӣ;�4�	} ���b��h�$ott��x��0��J���MQ�����=��{�g�:��I�R�C�7SZ9�߱��tC�P��MH;k��r���������sƮcD	m����sl���"Fј�{�^�4��op7����}=�E�h�8�әV��P����D��DP?�/��=�jՊ�1B�;������ʁ�h��X��#t�����x�t>h�S�\{c)���G�h��|�A&�G^J������n�mĈ)�0j�����k2��*�'��(G���!a-;I���-Q�ٮ�x�q6Z���ݰ������bY�A����a�h��y���v�ui3}���C��\���ǁ/5�����K�s�%�R��Y]J���5Dz$:�rc��]�PY�_��Z��P>#���<�a��c�!��$W���Y*O�����,�KR��Y��O�p��#ěfb�WM���P�y�F�5�ȴS�%e�r�49,V۹���;��_�w�P�%�ɋѠq�<2�bY����.�[�E�]tC��m]V$���g�N%�P��Sv����g��JY����,%D�_�[����g���)�ٻ�2�Gf���]AD~���V;]��Am���Hsʃ�٣��c����-Qf����0:�g����b�- f�$d��>e�:�%�yU+�oc�D�~V�����?M��4�ᦅ=�y�`������3�|����ϊk�AL�M���?�,P�٨�gppt��XcE<~I���M���W�&˖N�L���[0/��iF�Vb��g��j9nJ��
�/.�2��eiaai��8����q���O�x72��cQn#�^s�˝���e�5�b��1�).�;��k`�W�Ymj��U͡�4{��!�'����	��G�1t�Z<'��{J���T^� 9�>Y)�a��)He�X��L��ǧ+����BGG����P�Ms�f#I�3�稍>��R��n�����~��'�u1��5ݻ�+4�k?�XY�"Ӧr%���B� �ET�N�K���y�Y,>�E���
�B84�?�_
𘗨ק��heK0��@�hBd�T�+��&3ַ�m�e).y��F7��D�- �^�%�Y휕��'���@��[�Q��07��swov��;�U�%����6Γ 3���b�A�����m���ׄ��5�$��F�)�x*r�<�`.�h��a�8x��u���Xj��� ��G�~�o��Ś?m�=;�8;O�i�f�GJF!�:*�(�K4"d|�MW �m�v���V�t�q$�h�}uF�g5�U��Z��\y�sv��o����K���[�E�a���<t���Ҋ�
��$��tæ1�˒�h_���m-3O��ow����������<{#�������C��\�hn�_x�O�"�\@�v��O����߆�xi�F���9 ��Y*X�Ne�����ӫ�Z�����hVl�����)������%�1�h�eX��ئ���Co��Q{s��i_���0�4T+5��qUQ6�{���
Hq�}7���e^�XgX��t�.�zy
����be�ED/�"�s�J���n-�)e���a�T�����M�r�΋���RP ��g>S�"�}jpn���0W��I*!e@�ll��4p��2�o�/E��}0�ϭ��7��B <1�T�+��	�0ą$��j�e�@�rN-e)�"A�з��Qux�7��0Ys���Of&����N���*S���4��u[B|�n�C�IN9h���LI ��PN$�0�7�[.|������t�I�[\���D��|�-������h�$4� G5�i��m|cQ0��s_���I�C�G��@�G$�!���b�т���^D�1�E���+=E	��˚G����G�1�x���D#�M��Q��G�����9<�f�b~u"_�-$��	Uȑ���5Za)�z	���Y b���),� �r�6O�Yy-YK5��;��G;�R�����[ʤ�`���v���oO�;`���l����ѭ�=&�=��_�61�P�����b,L�s}�@�%>��rY�C�3�1��ކ��1Bb��)���l.w�*�����K6]�wk����Z�x\Ġb�/�l�Z�+Q��Ѡ�O�P^�?uO�u��3�L𨑴��̼��+�s����s%�o)�6UL�[�t�7"D�%Xn��.�C�8Vf������躛�k�*a��m+��7��Am<�ġ__��ح�,���>�������U쐡�4�'G���� �3j�I�]��jXf�I6�>�n]��vƭ�M7�I��	q���	������+G	]T���o;[ J������!�ފ��m����#{�f���	b��"<����>(��h

k