��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|Cd��D�����������<��ݪ��r�~���6�s�%>��h��aq,��(͏�2�~���ԣ�㮏a�"�f	^��S��E���b�@|r�-��V]3n�d�YR}���2�B*`IF^4�������8ʯb�2�!`J����0�L����7���6�t��V�_<	s��UG�SI8),�؊�FD0��h�d[����d��I�GQG�Q�8��h�z�T�߰�
�d)���8��|��-眴<<��^��w�jjS)տY��X��Z(�Q��[���&�l,"$%��Ď5~�L���&��fh�B�+?K���Hi��0�4_�50S�1������3��p|$�e���Q���G���j�<|�GS���C��i��	n�ڐB���H��ݐA����B�e$wٓI것���>e��$O����&��9e=ѽp�s��Φ�;L�&���gsOO		�U~ �gɮ�l~���o��� �����0u�s��{E�cîؘ1s.���`���i��+�S�s-v�b*�L5�F.�p��@Ǎo��7倭m��o_�/�F6�b�h�N�����Aw�-�q��ֺ����Ӡ=9��et
�}�� �����|N>�=�$�4H����P���nP���5�,�Γ�u�\|�L��5f��xM���@k|��1?5skġ�>�l,e�qu85��=�^�j$�i �.�:���z#/��&�}ڬ��Rŉ��Dy�CT�b+�ă��祑Q��6G�^���@_�ڱ��$�}B��qT3������XT3���9��ap�bg*�f����fYܽ��#��[����g���̒��YF�������,�M*c����J-�d"�	���Q��u$ׂ�鱄��>1�;�J
C����v��͵�;ً1�A{$:�Ŏv�!��H��R�I�Rw��?k��W��r�Z���<@Sqr|+�	x��B:��T���rW=���~��ӡ@tj��T�`�����u�o�O��9xM��	�B'��	�ۨ��>e_���ca�4�3o7��>�o9�'��{�X=�\�Td�)�2� Ǽk9'�AߵXs�W�32*M�0"��i�~�b��<����'�Z7��a����3`�W%#kM<��%'��� �v(�����~��Pg�Ú�����*}��u�D�\���J�O8��L��2�����L��/%��������̙z�D�͛���➁kF���!]���%�En���(��;�l���S�)��%^{I�0J���|��>�Düƙ.���eF,N_��{(�?�B攊�`���'O��[�\�3��3Y�F:�Ě�� i�4����;	ީb���a'ѸѻUo�;�7=�)����c��<�`����v�e�	=4a@�nv�~kӰ��1�{iܱ��d�����w�04�3 u������<ߵ���������6�c;���g�>F�����ky��"MK�J�;[;�d�A�E6Ul8�`>��u^U�S����x�n��q�C\�7�
�����Ʊ���.i���'Q���|�w3��Hg������S�M�h~���t:��J�{X�2M^�A�+Ѱ�d���LIu&� *6,I���G����և���h(�c�G~�B�~���/X��� 3��&*l�X5��1D�j�`E�,e��2tQkEŀX��u)�*>����e��_���v,�f̱�T�������aVH�z�x�{s�o�bN��&a�'H5~W����ю+�'��^H&&S-���dZtb�W�A}��Xډ���/�Ɲ�S�H��'	a$>�/�s���X�\���������x���=�O.�}f��H�B©�����'����kYƬ"�.��k.����P�+�Y�9l��s�,b����w��=�l�%�N<Q��Γ���c���e�����3�2y�vҀz���;�?y����4)��R���`�,�J.(�6%~�C"a���\���������p(*�GO�IћZ���b}'���5˖�)�ؕ"�Ԟ��=�)]��+���E~;�E�B�FN�b�VCƲ'��0��Ǉ
S���.3�|B@�x��ss��dv^�O="����q*�G+�ѫ�aݯ�C�E��^���	�����2���b-޿�KN�z3e��f^�b�=��}8�E�QŮs��9@����i�zYbW7c5���KF�q�Z�W���!0�*�N"�2Lk7ә�,����P̽�֜]���?�US%.�:H����F�9��B�7�t�,�;�+=n�����T/u�H�SY�wŕk��P%����	 ���n�B)J��͔h�ś�
ˏ	�ݞfݡ�%�	p�0M-~�<q%�8+*B�c9l���ەS?z��Љ8G�!����J�ɾѣ�8uy���C���v����hD���:�7�:_0��gGL �(6C1N����5Z�kO����߸�s&�p�*6�Q�@qq��|8�C�������4��KG6"�/�%{T.NFU�����Ic=��#�1m�4	�߅L+u���()���,`�ŀ6P��i�I���_Z�9"Ӄ*Z�fU�Х�;yl�F�ݒ�VӏSD���.П������-�pC�|�Ԍ�u~�O����JYn�QgW ��d�aIT�dV+�b)���c@�����D���5T�lF�y�q�^���ə�(6S��ɦob�N~�^'��5��A��-��.�e��`�|m_Rуz��/쓉�Eu�ػj��N�}(���uC,���?���0%xm�sQ�sY`2|5�eC�s���YK���`�Z��xT�)���f�2`��e4�d��+��3��[���5`U�$Y��ߒ��>v��E�"p���a��/��冃ep��}�gk�d<���B��/Z
���}� ��:ITC�Q�.m� �.��[�Y� ����Y�U���6�<�L� �~�*�R)T\�G�u�7Z�ED���4�I\�L�+s��]���\	�m���;x�3<�7�����)��PͲ)U�ΕN	�?S b�'��}~
��$�XC�J�ٿc�,�[/�f���H6XS�Ӊ!l>`���Ds��8�6�z��^�����NI~��VX3�>�hK�������J�>�