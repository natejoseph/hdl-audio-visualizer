��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CB��na������om�z��3 �$,x&^,�0�[.֊�~�CM�~�����U(�G�M�]��YOl��\�8E]��^d�]D�{����9�O�Ŧ��m��}�qJC�ܖ:�s`2�,Ҥ;��F���,k}����֘ï���̶mY#{�V����n�5�E�fZ+���bkMp�k+�f{�˯ b����9L��{<�A�����������&(yR&bī�2��/��ֲ;g�عs|��!ǭY��pR��F��-*8�8Q8�����-���8��7��^�=��.(-V�.�g}�S�r���y{�<��{�qE��_�z��3v��\"��#���T�W��T��(#��1ۀ��햣^����	޵����R�Ȉ�Ě��a�g@�M�����O�8�d��i9�ڃ��1h�NF�([�|�5i�9�C�d�=:s����癟R��p�1��zl*���$��A+���Z�k��>I'���	�n��aY�2Fo��4e�$,6����
��Q^Mn��0��B�eh4�*�xX=p�¹�X���)s��=Йi?�pi���l�~��L���,��@�bEk+;:����m�M������8�1�������T�]X�9�5�����ƹ��d�u�%a���פ�G�1T�x�L]D�.�����	��� ���Ȋ��S�!���2s�Z4Mʘ�ѻ����SҢ3�_:���"�~jXo{��H�~��Q��� w���g�Nr�5���LRŁ0Aye'4�
�&+��lW񃎡�k��̧
��~�+��-W��VHfe�RL/��������eF�S1'�u��I�b�槃$)x�2jR#_ܗ�Y��0Nh�'YK�;&�׿Y1�=#	p��j�4�(��a���&Cw?óh\r��/o�J���� =/������w�ty��L�E^o �N��E��#C�f�;��Ȫ���Ѿ��u��;7:�Ӂ7�
|]�||�2�9]�C�C�V�>s��=v~t��BR[�D%�Fj�|ǖ�:F<S��6\^n��<�e}Cغ�5B��_n��Z�`�A!�8Z�0�	&���$�68�Z��W+����y\9�p.��?֚\��.%3�ћ%Zs��
T+����?8�CX�i�|�:.�[Y̲�����N�E�	�3FI!s���R_�DAq9�я�4�r�Pz�/3oft)E�Ԑ�q�EZ���ܡ��47و��{�v(y�k�ӗ5)qtO7IkTӵ�t��� �I|j��Er�/[Pwm&l�'�S.������Z�������B�wm�����'�oc�"ex�a	`e�T �^w�`t�1w\�O��%��Bq�h*�֟�i<x��fP��Uߏ�}7��㈒����8�Y]Q˾�!�/5g�7-
�1(J�ގ��2�7�.��x���`�_�u �f�%���BU~P!�e~�B�d�]�H��ɀ���T�%�z'vw柈�	�I���L710�p�Q:��:���9y�����z%a{���0N�3&�5:�2��u#��?� 0�כ6`gC ���h(�d�k|��z ]�����;饍��	̔��\����΂H�(�h�S�3=H�[��i�	��/륦���7�+�c=w�b0���0��f��޴�3:��nm]\n=���3k!��]�u��	mwOf���Ca�������P�P|���67��YFl��ZRC:G
�с�K�����A0أ�Z���ɗUY��%��~���}@+��	�A��y�/
�mA�­�yNI�g��A�#���Y~J%���ָ�%�z�p��1�J�_���JC% ^����H/�A�J&������t�?+�:���>CΟ�r�cۢ���=���e欻���jfG��*�%�.䷥1���a���]��Sn�;i��9hȂ�+�\m�~��nOF��������Vj9˝�?��r�|��
A�X�<?N�~�-��a�sԋ�r��=�����d!1E�*�����E�̭+��QdX�]q3�ϭ����!��̪$�?���+�Pd2��oH_ �f0K�v���H�+�+���j�o�e.t��w�yt�Hݚb�U4Y�Я��CSyq��o�[f}�/��$�J�x��G%>�ا93 �F!%�9A��zo&�,g^I��,�;�z���Y�G4�nH�=ޘ�=P�K24�!ֆ}��"��P�]�����)��J�Ln�J�	D��'Ʋ���-�oȤz��i�j%=��P�:)~V�/E�=P��Y������0X�}�ꉅ3��Y��d��1������vZ�E���I�R����-q>լ�+�	����|�k���Yΐ!�*f��6����:� �I��Jt;+��ɁA��b;��M	��k�H|�P5^Y/82����^�p�7���.��E�G�|�0�Z��y�����: ���h4��D5�ݦ~#,�.�乗��3`/w�C�\����ϛ>�b�hu�1Xk"��O�!w�����V�%�g�0:m�����ͣ�ҰXo���w�^"���Ш���a���fg�G�r������^�A�=�^.R��A�G��έ6����#wǖ�*�pf�搔���|��M��v��S���0���"5���|~�$�f�Y��݁����.�05����*8Í�RZ$#=~W���5X���q�@�/��`���o��=f��#�7whCMj���pb�+*�B��懱��2"9��Z��?�Lu�ժ1LRF���(@���d�soVwhS�.�:�>'L<z�k����csQPe�3�L}5����uEf������ *PO�_���?�p�爅=�$-�x�7��O�H���":�ͩ
�P��r�CWˀ���Eȸ߰����~�5aO���:��Wg�����X9��~�t~H(� ���
�J�Oa+l%��m ���u4H+RB]]�MQB����� B���:|��?�	"sg�m�4M�xK��f=���_G]�a7,ي-71�"@��'�,� u�}�D�z�.�Lo������|-�>�����U�^�.�������g�$�"�� yې�.����Nn�'�hbs�ؿ|�K��&g���3��C�XyV|�EY�[�����#8	Oi�<0��;tבQ��w��	&�t_E�L��@��PdK��ڥF�e�4\���إ���T�۰#��*�P����Ia?�rڹUJ�΁�0�-��?9�v�E��U4zV�0Wv�l7�FV*;��?�j[J��Ek������Jr�:_'���1cSï�oS�C�V�;��:����	i]���[��NTúTź4Zh��o��&��;��UpI�8r[�������0�SP��2�yGą����]��#9�w&�MG!K,�R�LS(��Ӗ��ȳӔe�<�� ���5/�#lR�w^Ŋ��>qD�8fv�*7��Q�T0V�Rr܎��n�ֈ�bNj
.���B-c��`�L�U�� �n�݌�-�8��,����B�y�8<M�ik�0���{X�='F�/�����4Dw���mw�BY���
��R�IJ���r��Z���rhq��u�P<�	H��
N�y��!a���v�|5n��v�*�;V�ߨLL�Y�C;�O�h�ϰ���L�?��!	�n �ܗ]��"�K����(��?2/�2'R�L�	=�b����b!c����S��2���F�ٟ�{\���^���:�8�G���P�q���:��r�ﰳN������,�Zd�ՄJ`Wo��7׋L���֐m���m�k[u�%����?1���Y� =�j@}
�.���WT63'���s��tR ���s�����k��85���A�}�"��hK�����]�%�� 
j勽c�9��T�;qM<	�� ��}�-JR|�.��ޞv�)		�%�;�w�C��Gu�+�8��*�H�8��n�ݔIی9�@Wg�Y�_$PA���J����n/lsKcA|�73g�pg^�ՑV��߫o��W>��}Xެ��s�qC���n)�d�Х��!׃M�Al�X�0@�cD��=����1c���Ab���?ɦh���?����m �-"�qtFah`���TT�RY�|�ʵ�%4�J��?lJ=�L3���ؽ<��ޕ%%�ju�v-D����qc�c��*��F�A����+,*^�]�f�j���H���\��-C�4���?�9���x/���<w3��w�KTs#T�ҕaq/b��8�ĳ+
��,�:�OS�=�k[������|l^����ջk}f�aa� ����@�2�G^���\�h���w�9���8n�43\�?2����nr�3�Ƈ��E߬��<�/����M) M��.\Y7v�/�W���;�uaۡ+)��0>.Qw�P;�dXo���j�C~�S!&���i���1��Ų�7C�^�#�,�L#�WH�����L�o����7��s�[
��˖����pM�,_Eu���Qgw���?�^3�����e�9�r�^�w���;|}��P�mIź�
͞��Iq�1�Cg�B8���e�[�FE�W ��ף���7�*�}�c8�Gsa֔s(>�0[K� rՔ�����nɥ��E�Ӟ��nS4�h�AGe%�������V�N�S�B��b\3jL��q�Y�IX��T�^R��o�j�l�g�!�"/$���%�)k�����V63 ́�=��2��&2��@�6��.�B\#��a=�P�퀋&��v���+����(�A-�k�\�������!�WT�}���xآ��f�ą�g3�=�`������<9F!�ȜoEYL���8�h�-jnS�ѓ:gS����V7�0�?�Qcm��۪'�`9d�?~�B������W��x'�S͈ME��i��q�cd$a�_�H%��� ���W})A�`Ev���)ȋ6}K2�ໞb��5���}[D�ôcO"Q�]�!�K:DqxW���c���>\�������vdGy zL�(Ma�Ư��\y�ay��z�1n�Pß�����gC�T�j�l�j7iHB��f �J�����(ڧvxe�mWE�5K=���u���[�����8�N���n�l�F�g-!�7M��B����Up���cl��׿�5'�`�z�g�V����U���c�y c�m�c��&��]y2q&'�ɿ�B��C��aܢy&?�΋��t��S)�����X#���c+����!��ѭ*��z}rk6 v���
y|Y\Gb�FɪL��f�����zOB��t����}�=,��j��d�ߓ�K�r1bD	]W�z��"_N?#�K�}b�L�)!�y-��yłiӾ��yk	Y� ���hIN�~N�����ޥ�%�>u�b����T��\)	xzu�`����3����tb#�QL��qТ\��e��V �y[��N���u��dI�iT��S`R��#$���D��]*7p�t+��1WXll�"M���=n|]�����{�y�Ύ����F�:���W�M~�̣��%����}�O�pUx=Z/)L��99�+`*��hl��1J�]<�ng}FC�w4���-���Z�����H��9Qm��}L�q����׶a��z�[�Q�U��;��\<���ʬ�'y�w��H/ç���	�y'x�z+� W#ÿ|J(��m�o�8_Jy��᧢��l8=!��D�����ޖ�
���y��s�����Nm�;жp�Þ*���rY]���بᇘ����ʹګ]�H������`��~��\ض�Z�] �^�s}Wox����r�;��05N�oC
��힁		���,���(l�HtӅ�{J|�fUV*)�����F����!K s�Sa�e��k�]�d���#��>�'d�R��ԫ|����'���,>_!�S �/�)[�3֘i!_[1�DPt�sD����%�>���z`���~uv ���f��� �k� ��H+��B�Uͧ��9��۷ή΂��T�$�U��:e�M3����p4��Ϙv˖��=g����6c�rm�KbPk�Pv�*z�Ѕ\�O!|`�;Y�ӽ����`�W�4"�U,Ec��E��{>�1̌��7*�3 ��h{_/e-�uo���-]���H4�1f�#Y���C��o8	ʅ�#i |��8@�+�FX A,��t8 ��5Y��|����w����k�98&�!�k��#�}6<8��i����8�yC����ߨ��2
�0*�X�w_���b:�M��x��\>�-�v
��[#s�X��p�*B!�aJ.
��Vg�h�eВ�G���2Cby Kv���'˂9_�G��ajC�7s��5#C%�����s�y?W"���_X��:!}��W#��2��R�=C��;Y3�{@_���OL�+��?��/�x�td����}�\m�:���OQ���֊��R���pJ��ˇ~���G�PD��Y�*?`K�����q"lb�����;��="����ʷH���]|��چ����;����X
"�5kZ]�7e#�	�ϫ�iQ&�붞��l���z;2&�t��'�nUp �}qG��H5�K%�SH�;�����hT�v\�>r��9D�d��z��7D��Ma�t��훵����Jm*�zg��I�4�p�����	���H��̲�U"G��F�J�
�k��W6����9:����s8��:|����S�|�鴪���Gb�)�����s������ �1Q�-<�k��"�s�#�+&8�@{L+�.�o��(c��[؝/�c��o�Tڣ�a�(�9^�v�%��7���4�%��0gﲳu���ɺʗ�q�1��cb��	*�١�D���:&�� ����8IU� R��	������ ��R�`�~QEE�ak6đ�M�m0�y���Ͱ����^]��%GIGR̘�J3ϪՈ}�TkI�O��f��7��i�)$=�JK�d�=�S]��
]�{7R��s�%·����/�.� �)o�z�&�
πmJ����2j���\@y��>��/�����zb���*=w�#��ýF,k�Y��m�_�0�R��x�b��7�����U����=��&����4��?ݱ���|����s��Y�Z��ʎ[���`J;���05j`�W�4Մ����#�gT�Oے~���	�V�>{�кF��G�?h0I����&�:O����y$�D_M�w�1��ퟖp��u?�jy҆9-8�Q8�ϣ}/�Ф}���8:M��t�Eq��{lI��<_|�j��J�2��dTȂk�cׂ������
�7N2��CKK�9nҥ�1�>��8a�k����Gssz�����K7s�[]�kwu��Nx�������MOΛ ��:&���<���^k}D�,�L�t%CM�n�D�y�}:����ê������g=�G/�
~>>S�
������F���&l��o�HXjgz#��2��b����C6�����H$�N��;�*,Y4V!��E���f�Yr���у����m/2A������CZMת�[ˀ���V58�Zl~w��l#6iNЍ�%�c��UBm5k�=b�V����<T��<j���c�>U�W
0��ח�X�%���y��I-�E�r�8�j7��j���[U_6S��Y�&���)�r�W���Q�ׯ�sPߺej/k��2㟇~'�d�٩�B�Tk`9�{�La4b�l����ܤ�u
��w�g�}.����S��D2"�"wgIj��וY9���P��k���~,qZd��lSS����KU�`�^�/�?u
��}�n�	�DVe���mK�׮r����x��70�=�����׉��ʵS�MJ�?���!�.����/B�-T�w4#6�uXu(*o�U<�����V�6���_�u�?j�\'Qu���{ ���"6[ 1�t!�攕��{�'�G�&�y���}E���5�x<���������t4U�O£�+�SG��NV(�n���CSfD�C(WhJ�EM��\7�����9�->�7��i��z"��l7�k�
2�Ow�;�������$>tX��5�Z�����Q����a��^Gz\m��M���3F�n�r�� �3e�]����tW�����.��ud'�l-��gp�f��7�o�p��0ܱ��c�����=�\,��z�`sFF3���j&m�j$m��
U4�����}(�v�_���D��<��1��Lf�"�n�A���p�c�*]Ex�p��f嚁Ʋ�q}���&��}�$�z~���0�)�ٱ���D+$��
�=�BPfy���%�h�NC���\�0�T�-�bz��3����ϦI��O��L�&S�%o��s��Bq�?��G�w�ح��M�?C�ޙJL�4�}=��D��E"���ѳ��Sc����Yc
H˸:,��gK[���.f�$KF��f�� ��l5Y�6�����O��t�<�O�<���yRB��z��:g5K�I��!�b��!�pG�_�8.d�-0�ܫ|��HJ�@4���X@�Q�ڬBfmmɭ����oL:&o��soL���Dڀ������As$�ז�Ѯ���X�^�oZHbb����(:V����� Ģ�0�v���C��58y�P��x�$<D �� ����M��X=^Q��7��%�Uex�/�)�<��?�&`qa�L~���b�����u��ju�`�L�����L��hX�a����W��V����ף��9��$먪b�eJ��#�aW�	��3l�ɩ�z�#�!<�94uzv|��8��ʱ�x{Hy���2�aAr��SKC��i�������V�/�8����Ra���޲����% ��C�2dn��?G�8��;�ݦ�Ǽ�(av:�'qVO,���å��_M!��NK�<+mZ�7�m�NX&�4#��i���<v��ǂ��w��e��s�����-'QN�m��ꇓ��/~�ᡫ��ǚ*��n����虔�,iU��D6�!�E����1*��o;��D��^ (��X�l΢��؄����9�1c��4��w�� �[c�����a��z� Zqh�;�p�/*ՁO�˦�9�Q��6{	�i�2E4�să��r%����7Vd1����.��:V��꓁�'�f�$�qx@9�4���(�E�Ӊ���?eX��A�M|V.T�q��)��X�n2kQC�����G�6�|z%�W����ø@��b 5��9�j	�W��	+�0�M�:�X0p���~���-��Y����Zի8�1���|����xyj�^�x��^$��AmYI�пnC�C��49���A8h#I:40s�?|��1Z����NU����@�Y+p|����.�o���c�3�.h�t�Ku�.�'����1������a���ji3��>L3�L9jL����!��Ϊ 4�{�q#�ja,䫣�g,��	I�mL[�	��Y)���3����΢�$�Leo������T��`yFFm�J�����BEG탠�Jq.�D��Q���aYO�oYUDa����"�¶�t��Iy��m��T�����q�4y�����`���Ly-.VSP�_(@��n�V�5eF�Zo��pG�+�j�M^���/J�@�����
�_
p���:�쏕A�-��AJ�t����P$O�?Y�%ڲ�%G'�����,Gc#���7��&��M�9��=�:4p,�>"�w豬�1%�L���2���_Į��+�������BvO3v�����n��8�Q�j):��|����0���?��G9U^���m.Œ����z� �͸��cFد4��		0M9q쫩�AT��m1;Qk����j�J�`��>�Ff��ã��kyc�d5���(|a�#�$2@s�O�2"i'�pO�e� `,wq o��/���t�v˿"��J�8�����;yf��H�����:��fAQN�O,�C6e�Q���#3�h���ґl�r�R֧�
]�݇}��5lrynv�غ��IRY�!�p���r<�$�:"4�`Yh�h�p8n�)7���t�Z���9u"�������k#�z�����5�)R��Y��^�yA��iʚuu#;�.�zN^n9�.P��:�$�hk���q��0�q���@��A�#C�j�F�^�ߒs�ʁn����bo�Yp��k�ϳk��=���>��z���m�R�f��x��.5R@,Q�͹|[�.��b��y��噶�N�쀏�2����ú.�:���pc�jA�A�cNHpH���	��'��N���e����Uz�#XU0 ˰��p�P�1�Wi���@��W�+���W�3��/�����b�����Fip+s�*w�r�XQ
,�Lm�cS�yqg��d�:�n�ӹ$��%˓{�iRiKa�l�}�B�>m	���A9Gy��X��2h�_@R!���~�0S�{��E�<0eN6�{UN�c��1lD�,��A�>Z�����)���n��LrU�"�"�ciAX�ؖ	�'4A#���s�=M��Mai������S��O��4�qc�2.�����[���y���-a��F�a87�7�A�Tss��,��E��{�y:r��	��d��ft�}0|��K���_�ky��P�*CK��i������{��AK(U>7+ގք�0�Jj��;_�8�����+
.�I<�<�|^�D��5[���{s�p�b���q�k��XX�T|�q��OָUyq��:is�٣l�	����PS�Vc8���G�B�/-�;���2�(7��a	D��2_̙�iT�P}xW�k�Erj��T_������\m~��Έ�j٘N��Tq�5[.ot��$;İ����_�HJ���C�:�����k����q�X}
�Wkh�����w���}J��#�0��U�f��$�P�����:y��5	��l����v>��0��F�/8�$��"�(�s�1'� 0֋ ��%�2�8h�-�'A���=��=�"<��