��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CB��na���+.x*�?a��h���i26x&�,5�S�~��M�)��C%�~���g��l!�w@a��L�qj���G�_z���v2�2><o�)/L��p�G�
u��5pU [W(,@���:�E�WbK��"+[Ӫ.^z���Ȇ�N���hÁ�2��R0ةT5��-���s�a1)�$y "����4C�p�"��.Kb�G���㝸mJ�W�ٗ(qג���Rߩ��4�f�f=����2��Q�]��	� zc����h�҄ϔw

�+�Ca>�4�W�wnPQ�v-�g,�gG���A@�>G����:����h�l��=��R�J�_��h�}n��͉t��#ҽ'��j�9�q8x� �\a@�o�*�ۇ����?%u�.�ո@dL���?�"o��E8 �� NZ!{Q㪡W�g�쓼E@�����ъŏL^�'5�x��y��l�GZ��>A6�n �ؖ]kA>ӹVy�����ɧ!����1�c����P f�p
��^F]?2\�f�?I��&�a���<�^#"vk39$��r$�iH��X�$�eO���N�m8Ef�n�+��oN���Y�ұ�8H�`�eM��xc�vh�a���	vնV��hͩ�'N=�T&�W&�=��:�'���x���$?J�G���|J��}~O��u�ȶ���������"��pӀߐ���בn�/,O���Ȭ �B�]u��Old��-�N-�*f�H�1�����:ہ��Sd���;F�A�}b�UB�8̐������/���| A�0�a�X�5�ۖ�k�Bp罰ƕ�������k��|��!��%�+����ڜ洹G����Ə'r�G�D�a��ll��y�0�$�/���s�&�9�Ʀ�fj�ܨ��^��d���_�J%w?͆5�i���(iX�6-��^NdU����0OJn��/��cAl5J����DTnW���<.E�{��ʢ�S��k�������\�x�+_��?*4��T���4���N��� �_������9�|�'��PZ��e�l$̸��/�
��E��n�us��zXO����e����.@�ݶ�焕=FE�X���Z�ň�4�˥���kt_��F~G���@��y��`����U5��A���tyK���"K�WL��.������s�L��Ԇǡg#$,����{�����_"��^���<�Mf�����������d�>����~�HY�5�i����w,��G��8=��c̐���Mc�O��W�/�#�s�2�ZG4�	(��TF<�P��ѰX"�:��Mi��t��WP(,v]2;�[��ƭ�WR��VϻP�z~38�ƥHp>h�'x��e���m(t���ix4�;[ �Y���I�ۄ���c�[����z�c�Z�4�.��j�p֕��-�|1?�/B�i�j�5��[�����Y����RS]�@\�q��kj�L�~ǵ�eT�rd�Q֟qQ1�p'�6��O]X��#V��?��� Wi 9��R�f���=�\A��x����v��I"���7y�>'��3���3���@�H�g���?0H�v�e���͖Do�C�\��Ԫ-_b���>j%L��*]ߺ��v�df��S���`XgG�Q�F�4��u�O����_��� a�y��.�kZv��}ˤ�̴�$;L�i�m����}$�����[��%R�����'�Ȝ�3e> :ѼQwO�D����Ӟ/X�A�����y^�cTǑ����pF,�|7ģlsL
x���~q��+I2^�G��}�왲�)?��O��>_�x��Y&"��d��(ZoP:"���O_���5���⻦�q������z����o��ܪ�DV�����Q�]����B2�ʛ�}"��S���V��&Px~��sTg�,[�>�RŵvBs��-'%Ι>j榙Z��s��3l��$E�� ��Q:]U��q�O��լ��R�pniy&�?�D�1������᫱�U@2�u0����' v����D&���ns��SR�:nB�~�$� ��e2������$���0d�bL;g��r������t�ٵ��ou�#x�M�w��g��V��]�K�(��9�P��KG-}δj�#��V���k�>"���cӴ,a(.���YQ������_F����V��$*ʍ�îċ%	���Yh�z��v�dHTc$��b!��7�x
L��M"��@	 jp��y n���E��^� �C9�Rgq�Π�����no����&������<KtM���X�y�$Q����/췦	$#\���
{	��|,���Ν��	f�F,����#vn>���]��N���˂_�
��گ|��"Y���#>��͞Z�.�8�e����Y6dL2�����E��uY�s�+�D�Xdk���H�Cq��'7e9�L^ջ�p�o���qi�bҥeQG�C<$��	���C/�/�L���u�g����d^o=��u\��M`�0g�@�Lw�d��י$�%I.��FpYOw��r�*��RR	�>[W+Jg�y�8��&�*|� �1��xY������T��S��6�葺�L ik�fζ�G	<}�wL�*1��y(!{U�tW�7�4��[�zA�J�7X��^.'�c4b���L�Ӂ���Q�tN΢�O�2qs�2�O�>��=����6ޜ��W#�Lg���wIո'�{z
"�" ��˜�S-٣#)�&�u*}׏8p��rv�J����������$;��#���s���k?ٌtz�2�� S.Ӷj����<.���ق�e�`����#�]s���z����;�����<��V~���qD/��H36
n���X���L��e�]���wyO�����t��ɒ�7
1E�௨:��z�f�`J 0��J�1�?v�p9P�H������P����i�k:-Q���o��]\�Ū�"�E��]8�=��Xx�܃��d��u�:���up�16�A�a�;�-7���xMa3�ܨm:a����d��Y pU���]�ܭ�t��>Vɼ+���0G'��ݖ�(G�c�аgh盖���O3{/q% #Tq*�_���/��%y$?^@~�����m��Ե#���Å����5eZ�PVDj��66bB}EtD�U�1��ǱGH�]�@�
ab��;�a;�h��c��w�2I�u�o�qk����r��޷���Z/��j9bK���>�u�`C����-elv@7E2�@&�W��(����H�F����*-��;�$�K�O�gK���(��B0|D����h�5ß�#�A}�N+��S�Q=�<�~��E����*�
v��#̬?z���l���'�;�]�j���������X0Sh���`���(c�6�qZ��y�My�����Ie��b���U>�5S��:�m�e���ip٪²�|_��z�I�)���#�ؿ�^�e�\7I���C�Vk>2rm;@��<����Y9��7�"h��']V֕��s����Da՝�H*�ý=�p���J�O҉!��̙��3�7x�p���m�j�we��C��g���X��#�S��m� qi�,���%&cV<'�8A����䐠 6�Ì�|h4/�8�0���ϰ�1BNa���$s�xs��l]֣�S�����b5h�aϮM�(n,I��X�~:�=��~�.ђ`9D�*M w�%WW�-b���B���wC?AJ�*�>G�c���}Is��ݘ���j��;�Yl�c7ZI�)wC#�f�Ʉ���/&PO#?x/�Ѣ�ņ��m	�YA>!�?*��H_���o���ua��a��D�����$3��dA�1��P�Z2�-}'"a�h��.tM���Lo���yh����0��n���E�+B���ORCW����N`)^f֡���� ��@�䳑�NnH�^�v?S�~#�#��=1m� �����	�ڨN���c�L���G��3�1�kZ�rMD���D�ˠ]e~�c��g��&h�4,�-��88���>+s]� �^7��%ʷ�ʨ���m/�q >��WGU������4f���U���;���� ��B�ƚ�.��=��h�xvw54���I�
*^�ᬇ���[A,(Hވ]�ѳ1��-����@�6C�|Q��X'��&\��ɱÅ��l�z�-���4�j9+E�V��=\�H~Һ���� tJ�r:7u}L!�M�`\K�6����Kǎ̽2~�_X�r~�Q����f�P0s��K�pc}l�Ri{�M5:�V�\��_���UZ�%�oh�J�M&��˥�^� R���4V � ����k�:M��9�C�%n�7olm8�PC�D!c�� ]�7��?���p��z�G�vE�u�ܙ�t]��(��k=}=��Vn�<��F��pmg|'�B��c���$�Z�ÚRuQ�â��.� �w(	�<C5�E�s���Q?Q틪�P�p#n/�|2J�2���R-ؗ��X��1�l��m���|@���yq)cB���/�
�o��d�fٽOvQ[�%ZI�h��o	Rgm�D������)�4������#�5Ds���n:pbv�t`bp_ۥmiu[��6�2D��?]PQD35:���M/��(�n����>���4�!�e�=m�,��{w9�CK��R��&b>�z�etNL��N�^�D露ק��dc�:�l���(?��::)!����{��A���җ6h1�9��j���2f��<�S���gUa_��C�c�<c<'R���h?=�����w�#uu�	�xlzv��K���돬��Ȏ�y�i����w ��fE�@��λF]1��*uRQ�a�.��/A�l���}�P�����ٰ�5�Z��
��I=u����%+<�4���uCH�%��o$]�s��)&��nh�׵�D��/��[lP�Q�������[b��&�� }�����B��%\����4"�⛿�ķ͔T��ݧ#>�q��3�c*G�?XF)�82ķN�Y]�-Y�M~~Ƃ�euh� ���H2�k#*:G��S1��s���K��{<�ٳ�[����5����ufE�PO�[\H;�:�e�v,*�F�Q��D� ��G|��3�����Ʈ�q�
�L�z6�mX,��VS��o�;�H���3z��iedZ��
$�_�[)�M�`]a�o��)��:����۝Ӫ�����V��/-��߼���"�'�'���ӟe_ݮ/(����\Fi��=!\�ɹ����$\3�j�hl�d��E���վ=�y.	��+�)�hď�q���[vh��s���?�=y�jW�@~���'�E#3&Ы}� ����\@U۵�޽��^�b ��Pt4r&U�aKT���@��ր�r�`x�b�S�h᫘yYR��4�\9R�������۷%�Dm���ն ��.�"��#f�v�������//�F[{H�UC�%�����2(��0����.������	%��7�Y�0T�c�Og�OW�C}wS�Jqĵe�t�2�T�R����¡.��O ϯn�z�E������{���߇E��@����5�h�.���e��u4�j���TJC������y�A�-�<�H`�,jj�����*Dec���ZC����aO�٤1���0
� ٓ���niݹ.�!��,VA %��x��N�J�	l�0|o�_a	�$�ME�	�Z�)t���EJ}��za;���T���lSM���?re��Pd��Ey����<#� 
h�᥺9�� ��7�R���aS�el�RZL"�Z�{����˞�a���Uk�R��l�n���;�?���:�n4S)l�!:��N"�s�b�lzK���YmG4m���Y����)�~9��B~�����d��%*��e}͎_��P_ez�S^�AM��W:c~�?�tL��\rZ���4�l�#��\+^C�
�Ђ0��-͓]G8��^��S��;e8r�mC����o_M����x�� 0<����t�E���rP���cphM���X:pS4�c���VK�f�=�O��,C�S��� q���,���Z?�8�lWyٔL��D�F�#���ͨ'ڔ=�G��|6<��8�\����m�#��6���G�n���ޒ�D�fDZ�V���xk|�U���q�Q,R�W5h���r�_����.��>|~Yv�$�@,Wv�����_!Ť%�G0��q{��q�o�v�B)���N����䏅�!�ޢR�/����|^F6ʟaBڿpAT e��l�FL����5��)�����L�]����jC�bD���Q�S���!V?�Q�Ӵ��=	5:��t������7{�(Ŏm���m�Υ��Q�sǚ�!R�!���%0�������C����k�?�Эf�1dkJSjOG� ߧn I��R�?΂	y-=�3�?{����.�#�"P�b8��&�)2�RZ��:wiI��J\(G�������31���HlUO@�vP���݃����X�� t��Q�@����=� �̞���$Љlޱ��-�+�x+�M�{q���F8]�9�B���������n*�Z��V��xb������U��L�:���l��m֓�|0��RݑS=bG���]'s�r��Q�^�\��9���bN�5��@d��4j"�ƽ)}�f��/!��u��D�'���0-�Fq�cX���z��r�$.��ا�32mݣ��Q�����B(� �-���jgZ!���Pm����A[�n�w�o�,{���t�����iM�D-1�K��p�<�k�=���|St���E�Lw^�n<~����d@�2.R�ݣ�OJ+[�-t�ٍt�s7�R��ܔv��ݣ��տ2�RWvK�C�%����!9H�<Jp�
R��V��+�p5m��5�S���"�*.x�����j9/�5��]��ΆLU�L�F$�&!���R�ӧ�r��e�/&#^�<{�sR@{��
t�.¥Y���� �ZG��a
����))�;Ʀ�g�܄\��	�~"r�\7{���'�eF�k���|cI��.�~.�鶵2MR�49��U��3Rʒ���c'	Z��v'0���ڼ)�����^N�'1ѣ�o�\�US�5��H� ��b"eŐ@�5���S�T����To�vܶ����V��ۚS���@_��W�!|����>�ts'�0��+g�ީg�t[�9Zy�}�gq6���k������(�X�b)';n�D�k��\��w���&:�"]����Gtf
�R��=���؏���[��;fϮ���+�f�"J�k>���v3S`H2�:�d��tbE��S�|��8�x6����6ѕ����,�I��e��~�����M�^a\���W�1!��8��5./V]o�[���G��~�*̄��7� ��h@��\��J
��$O��ed�Ę$0���'D�{��Lk�;�j����K�y�����iu'Tv�ؚ�1��M%ǥ�w��>$0��)��jܚ�XI������=~Ј��hK#��st�?�?��6�"3�I��*=�p����L��tKS�&�C��ʭC��64���R7�E�K�����i�S��cg�>C����-���]�OBz������3����� 1�b}�������cʁ�dq�.�a�^���;��b�t]<J���eךc��ih��S����2������__�4[z���|�j�|���8��D50_��u��g*<P�T���	������3��ې�yⰾ�;s_�;�<k!� n��0Dy!-^R�h,�{S���*�{��bP�ʊ[�݆��P!�&=��?��rd��hBH[y���'���hN$c+�3�1P�i+��������1
%Ó�-+\t�&}�P�>gF���z��Y�Ϯ���\��o�@y���>��ki6ZQG!w���g���g�c�|3�RqP��WZ��}�9��z1t�E`t�E\��X�6��M��w̖w1��^^a��to���Gה�%��%�xƧE��p�xw>�8{q�B_m��
 s���'Ԧ@%=�Ԇ_�{'�4��V2��J��}!����f���7�}tɬ�4\�{��h��|_k����
)h��E.�N^����xn�����^�Ob�����PH��㥺��?�H��|6.�%��CwI>zfh;���]Ml"�|��5GB���G
�F�i2�^���p�bù�I���x���ۆaf���4�D�#�K!�����ު��ϩc�wC�6ԡ�0Ŝ+��?vE�q�	���}2c��+6F�@!�G��m7�ŷ�}�Ϝ���(M"������1bkѽq�:�?2�D�d��<r��\�������n��)�����?��ɪ���#޳��m�r��uQ�[����^}Dy��)����/��^��qeDۄ<Iۦ�(���EMZ��6 ��qi?xMRe'+�M�VC���l��R,��i��_G���]�4W��+K4z�~cm B����A�a�k�Y�/3s��L��pS��A.|�~<Ӗ����wLR!�����\JK�h����V(H�3���V�?��kI۠�d�:5�^cʴcyD�%��v~�쎁@��I_Qib�k��n%e>7��Z�����q��O�3��?,�,�7��k|���:MB& 1�%��dE��A)�����ҕk�6���ͱ�OT ���{���)�uم�o���zǺ�g+��\ޟ�_�	�T6�Ne���=c}Y��+Uq�p#C(�󾎹H��  �z�7,<w;�N|:�7U������^��\r�,���s���ిȭ�q�� .z4�0�8<@���;qZ��U��v��?�&&p ������a�F��k�E*Ջ�w�	ۈ;v�"/�k�AF��#/�y3е��0���|�ǔ��]+�ж��Uy��noP���g��U*�ܗ��2i��rN#F��s�|�0��n����wbv�^��.�����yq�Zy��x[d����0͇�L<��%�uDh��'j\n,M�AZ�X�Hf��T�l�a�S⑹��CBCЫ~:Y�1��woܐ�䆬��g����Zvk9N�>�<%��+e'���X�m��á�*�K}X�sX0(A)�S���^��.f����"�����pm� H̔�$�=���S)Z��V1���lz}a���KKF�@��AGts}I�G�j�x��bJV6ceKGKXF^�P��Y�}���^�@G�����ͪ� ���焾
o����!�7&>����X��eG�ȅΡE[��#�&�L������;�*U':����=�=���	=c��Ə5M���}��vR���	���	L7� �@�UC���n�}�e5=�өxo4�F���Z�����WuLϘ�5��^.ٻ$dY������f��\3��j��1ct5�¾#�s+��ꀳ�/�A�@+�w2�ŗ,'���Ze����`�"$�J��]����b�������{-t	��U�\��vR~�W���:.?��z��#����$�_��8m�q��!���*|�Q��(��T]�+�ە%�8�������V��Y��!�s���.���
��hB ���MO�����hX��K.KO�C�mm��ć��!\���}�	��Z?�B�F�h�a���~[C�%��J�yjhg�^�9;p�[� �ѵX�_��ʹ�?u/T?t��n�'+ˬc�BnU(B&AI�;)��-�:���N��2l-�Zł��f�B���R��­�H�T�(�@�H<NB9;��N%KYt7!�l��J��m,�����Z����m$Wc��$�{-O�B���1פ��R���t��� [�Rꁙ�}�<����⬎�WZ@o��]8-YqG���'���=9�\J+n��Z1* %�Rgʤ�IӇ�עN��a�q�{�BF�_(C+�4:��)�ęB� �r�C��Rk��
�ڛ��AO��Vꨣ0����PՌE;�	j;�x/�F2 %ʍ�7�J
��S��?e%r�<�^b��Ω��9��!�}`�:8]f*(��4��[��1{E�_����$h�d1�����\�2��A��G��n2���G�<K��S�L����LH.�D���!x~��:��8����#-���	'���~��4���jqgЛ�V��?c�ڄ����]��f=L3�,��%v�_��'Mŏ��W�����EMm!(�եhouB�t(�J��U�<Bln_<t��E;��N|���̴:�ڸ�����?׀����ٱ������&����Uw�`�lz
��#�!��}����:/���M�q�
�dRy��a��D�O��$x����`�C:�a�o*����X���6F��5���?-��_W���'�c�h�aP�NTX�Z�Y^]��1��v��X��;�7t{C�5z#V�=A��,.�����2�3��R|�>'�Ⱦu��ag��zv!m!0o�vqv�O?��3���ԝ�ƕV���`��r�">�T��䘴�#��f��E�l���.�q���$�^�!E��0@D�Zi]�6B��|���Q	�`dgD#�M�%�N�%>�l�����Ԃ�,�B���x�'gY�>�d��U�8*E��9$L�7	�Q�7�.qŝu�Y�wMx���^���i��o���C$/M	CJn]g϶�~TH~��:�yΗ#��kx.�F~!��~�����}�ix�@�����/�Cs��q
ue�@�ڄY���MuNI�syG��FquqH�]N��YQI��ip�\1���g�+a�g��.�~Z%ۏfG&�ju��l}����	��f4VYV;C�Α����t�H�B��E\ م��"���t�Lf6�w��2�xu�p�W�pa��~DY��]��lP�l��Q/EH��î�X�E�9����O�;C+_�(���ҫ�ȡj���^����pf�n���b�TN�����>�yu�3��Jʑ/�vߜw@<�C$�����٠/d��i?K�\<W��\��U@W�`����Za���W(42�(J�
��\��[H���-���z	u�!͌��K������W/
��H����?ģ��w���h�{� W�6(Ur��\@�
78��� 곞v�z�n���E���"A�ꕪ�8Z���=p8F��<�O8� ���R�,��}�r	#J� M��j_�ż���X�&�I��+��P-�3�=���|}$>�1�H�wq�fD��+�W�l��~8����*3�	��vK,)h�s�#����{����/Zf�{���-�.��>ص]�ih�[+R��GZKT˗C0��+��_Q��R��.j���+n`$;���$�f�u�ω�S�F�|���j�dD��͋�u�h[{(6�Ct���@j�N")��c?w�ʃ��U��'�a���MP�uܲp�B9_$�I�פk�)�����o��F8:|u���
��~r@!�TS�L%���)�w���q$S��q��XD��q4)H{ � ��DӲ�'�T/��e�M��w-���3�ᶉB/R*�5^�9���}~���G�-�'u%-V��6�}�P!|ۣj&ǒGM�Kd������ � ������ ��oE��\�o6�a"J���W������n��R'<ŔA]3J�ޔ�&���xl�3&�i���t�ϊ1�]6�[���A���rի>i(��G���`x2�M�c@�$ރ>��?��Ɔ��R(��'1Fb��k���{E>C���S�5?�~L�G���Ü��v�s��)v_!�8<tv��p�������u��r\�����CHv��8%v�;	�+�MZ�=W:�HK��� ���&��QT�"pc&�%�r�T�|�k�0@�B�R[~��M�M&?x$�F��.4�9̡/(����o�l�Bʄ㈯��� �bB���d��!�A�n�4���b�cfe,��)�67z�����1���\ȢXi����=���оW|#�8~"�+��B�мA;��N��#��^!��9�x�l7��Q�0�3u���Kf`�`Fcٷ�4�$R]S�@��hAx���͵�����HZ��q�m��/����������Ͼ�CD�����tS7j� �	z��̍�"ΤBlv���)�Ѡ=�.�ҫ��~�)d�lI�i,������u2�;V��h�Z���qxlb����T��?A�6���Gb�.g�`9��ޕG܌6�1V_3��fA�S����i)ⷒT��?L��3�+�RT�c�a�4oIx�LU��7�f��Z�:�2*����9�,��_�8Fw��?`�0��$!=j�:!�2\�x�zg;���C}���놲�R����\�/^�Ör�(�Wg7+n�h$:Ǐ]�/)��X���vU^�2i��|'�aˉNwl�ˊ�g�UHy+�FZu�k�j$,1�_�h�RD�QK���s�$x��l(�>�yx�j���,'�kQ����Mr�$�I�ڠ���ߧ�D����jȫA�M~bg5���?t#�_��v9�(�K�����%c��4;((ʞ��{�?Uε���J�|{m.���}^*��������z�����H���k�|��@��m �v�����88?74jt�KCk�:�ՑH٢�ߨ�z!�Rs����c��C{�D�E@�1&��,HT�ثW=̽��d\'U쌍 K>����>\�u��1���1�P��uKձ��{>�B�s����a>}�k�o�!�I�[�c�1��K�Q���������5�G�B�S����,Q��}�B���-J������Ss��q@X�SQl����������a��y,���qH*N�^�Z�Gi�]B�KQ�d8�p�o4J� q��B��r39�':��#	d|��r V�8��I����L����A=+����F{�Y�)e\4���r}��%{�U{���L�"A}��O[ܫR�R�X��̤�E�M�JW���Л�z�^jmp���6eE��=T�a��A#�nBK#æ{�2��F��0|f�a�W��߯�H�b"T�����`ްC�Iu�{��'O����vR��p�2�i������"��c�$y��>-�ki����kR��e���i����`ʉZ�Ӗ�u���n��l ��?�2��~�y��Mi���|��U��aQ��cJ����j�8�d��F�hMٿeO���pcpb��b�U���L%;
�3z�K0���;X7)����ˑ��P3T�LV��>3�Y���[�ׁza�� =�;�Ԍ}9�(�%����L��Xz�S��rP!$4�t�ذʸøLa���ڔV"�8t�P6��7���&���T�2B��E�q�V��]0�x��2U�D�D������?��#.8=�+�7��9u�PJ�HH&���㴦_/Z�[�8�G���Yڇ�G���J=��#Tp���O�k���������L����x�;3��S�K�4)	�Glt^ t�aŕl��(SZ��2?3�In��������F�.��8�?1�cḷ+5F�R�%Rnn���n�P�~&�ͩ�(�&	#��UQ��Ӹ#�����*�/�9���@r�Fu�f��Q�.��-A�S�L6c��?�fm���(Ky�/��� A-3|d��B<5���S���ro�^r�j�g���BU���n��-/�^z ��R�v+�}��*�W���q&����g�d9	i~��RֆǾ����_�{�w�&��"](C���*�rV��.E|�/�7\F�6����Y�+~�r���`"m��Y�˨N�1����b�w���K�^�hW�"�~�]��)k�/=��x���KL����l6ڶ��L��(휐q��t���+�@_�I�~ۑ�g�٦0!�|��'�Λ]��XH�eFK�3��Pqy���ڏ&˸�*��!�������*y���i��ވ��H$&���(cN���d�-p�ٱΛ-�ܨA>��P��6	?��lܴT������i��b����˱��Eˇ)/�P��]b3�=�A,��E�L�]X����Q⦏Y�O�JϠ����Vq�^UD�ٓy���2\�����[J���OO���S�/~(� =7�ň��xX�=րr	Yk�ܐ	eZ\J�|�M��_e��8�aS�C=�� ǯ{�_%i�v�:��0�i�e�4�ۭ�V�m����P�0j�\%N^���K�����bqK�M�g65%'B�a�k,��U3����$��e1�C3aB�/O�65	.魻}�c�]}�*fY���|wn�E��ͫ���\���y�+*�2���c�R�Yl�λ��o>2����ߠ�nC�Y	
�)L�����^D��Zب1DȆ�+��T,..��ϳ���_����2l���-����ʄK�=�RS�����m�M��9��be�J=������B�%9���>�W0�U=��0M_&��vO>\6�>���L�;[kb^OwI�E��k�T��6,; 	"X��!���מ�!��)�6\����"�뽿��b(�Э� �'�T�
*=�\^��O������l�8���"�UVe�`9kt=�LO�>������j���g��7�|�ڳ��lx��&�JK>���n|q2�!j+��*`�ӻ4��"J�^��_��;!���e�g^[%ǡR��*�\�꯬KG�02���o����+LFL8@%{{�DCf�9��<�AИ��rd��X���$�	=�0����}�l����x�u(�R�訿����9���9�Z�]��Ö�r:��Ź7)I?���j�c�^ُ����S�t�β�x�	�H�"��F;3� $�7#4��yL4�I4����qY&΍/;�	|s�����A?m?[�ɢu=.*���Jj����߻�����h����\�����0�­BZ�C��T-��ɰ9��H�B���bhr���@��ǅ'�A?x�Y��QW~�=��0�~-�úK��9＆���g��Z�!�
=bzk/$b�����z�-ޝ}��w_�?��<�96��
@�C\�:M��ˏ��r>���Q���qm!ugw"n���'�p��G��6�gMQ���#W
^1G�SV!C�^���=їc#���aR�}���WS�(7IBK��P�N]��
ad"�A��:�9v{}��Q �͘�|��{X%�Q����v��LͶ9�S�+ �Y��?�*y�P��w��?�e��X�0Sme��]�(�g��\i�L����T�m�+��!�}�0ǺݪT��K��G�^�P'�7�Qt�!�[��N1��X�JE:���c
.q�VR)R���L4��'��\^���L8�}���ݍ���"�3���`fc`�1A5�*9�'�N��C71��k�6d#�w �ڥ�� ���i*��ũ��0���Q�G���K��?��
,(S%20V[�<�Eo��Z֦��ģ�V&@\K8Cweq�g[;�-�.'��-W:��4��Q�ing�2�����t/v�Qf�J�J�k�Ժ�t_��9��<�"��0�y�2�Q[��O/�iZ�y&�5Mf�l����$�������p9/KK��H�����5�Z� W���U�ZY�	'�4���Q�����-j������	�P�<�(�'�j;�R�� �Ea�/�dW�"�0��	�1��rh�y��E����>�4��w�4Н�8�*s���v��@g+˂oTMs��]D6�-w(t�nR�P�����Z1�����w_k���,�Oڏ�kr����)�Ե|�^�"WX�2'C��n��"�`$�o��@|*~	��C.�|�"�K��8T��<���-�Yy^@x�E�4�eT�~E]��w9�j�"�ԩ15�K����l{�6ս�mF�j���$�������a.�ͭ��j�,V
�Ed���]P$/~'�m)�f'^���
[�a�����f��F���%[�1�D�R��S��y��l�bcߞɵ��yr�@܅ñ��l�k�0	������ǁ/���#,��Ӽ�=X�xΨ;w�������;��`yZ�3!W�D��!���ڌ(p��|�Z�w��D�K��㘥NQ!Ͱ<����ҙ�Ġȟ�&�N�zڶ�\F��o�ۖ�`�u,��v�䱶�*:MJ�>ϢS��D->j�dG��;R	Q[5$ؖ���;s82�{��҄ՉoF�ZB��Gg��2�o��.�$��N��L׮�����#���+�D�96[��#DI 	nìgO����&a�Z��W����������b�yO��X���'�sfНa�;1op�K^+
&��"��MG�Ͷ��B��q����z��/Y=*@
��v�e�fH���m�ţ�qI'�A~���qd<&��O��!��h�I���L�r�Z�w]h=�f�AU�0�\
;	Q��4/d{e��IA�޻T�s#D>��TT�x�C�"�%�H�Vӣ!��@0�s�T߸,Oi ����q�s�f�0\��P%�f����f&v H^�"/���L�c��'+���7��G�F���!��>��*�%��P:�|���P~d���KtS���A��7�S7R�`{QCy2wz����"=ߣ��Ĩy⶧u��R�Ȼ1P�����͂Q ���+�K�5?����p���fKiՆs��-O����]�t��;{��#��&�N�f��_a/��¹n�,��Qd�������䅤:^��΋��7"Zʬ��$�����P��CG�4c��Ɉ^9������V�E�|�R�Bis�T�+ņZS�4!��Y��Tm�ќ6iO3���4#C�<QrG�5���K�&4q��z��F ,�W�EѓJ��8�x�

F���7���m=<�\���pl�8�ֳ����	�4z)��$�Y܊PN���lUf KT���"0��~�b���s��\�S�!���A����~�O�	��}�b���i�A昙�kR����ԙQ���SEx�a����8���=	¸�|k�"�dH}����p{{�T}�|F)[+�|��YCH7aǕ]��_:���ۭc�9�\�#����PKvI�?[��f]���&��-
����F'�\O+T�d�o���I��[JZ}.ID-o'@�gy�ak��̍�N,�(=���<�o��/�:�V�髫s�=�sU4*�iy�/%ӷoU���1��KaƗ�6�_Ϟ������VA�=��'Ύj��Q�=S@�Y�S�w�b(�#^-��Կ�����>��cWo}����ɛ+[�j9ֿc�����{Q�f�j��nC��썧Cqw����^9�g��Jn?���b�+2#�kf�|x��|J%$횞G��2C
њ���3�1*�6}P����{��q�<D1���ؘ��1������|��'ytu;T��V*s���2T��x��A�y�kBT�_9��]���~�
��I4b�>����In��s�*�,�z���pݺPg2Y�2"o~����雬+4�?������Dˎn�h�ku�a��k�B�>��/U7Y��U����o�8��Q�T�?�$/�1� ��9�9`1���i�&V�-�����/uR:_^��0a?@m����D���tD�"YBiv'Q�J�I���Pʅ���%�qm���S(D���Oz�D6-J���Y����NE�x.?�Ca�3�!��2���`ݻ�jz����������]0Ȗ��8���i
~aƭ���[}��( �����v9�~Ct�PRG@�O��R��#�^�3G9#�����m��K��ޙ�� �,���w��t=�`�o:��ېł���5���3�����	��� �UIF %���Au��_s��sBNA��j'�/n��`+���RU���H�e��q�|)ը��f��kK��Vs[-?�K��D�!��~]�~��ɹ&#��Ҫ�T���&�M�⵨P%���Ӛ2E<�ŦQ`*`t䙢�h��b��#)H�ֲX���z�T�߇��%T�ӽs�:������rR�`�3YFE_��?��<ץ��'σ���m�?c�S�a����Ǭ[�D���\�	&�<Pײ�y�uΔ��)#�Ƶ�f�K#� �����v��Vs�gh�]7��"�����f����jN�rqU����'��?������ࠔrֵ��