��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�"��6�t۬���]�U�3j1P
���a�O3:�K�*K�ʑ[j�� ݎ��d�(Z�D�� 5C�U�]~����"���F2W�=s����ip"I#�����سVYCp�}QZ0�W��r��)��T	L��4�,g?�F�1Y1e����.����PW��$�39K��/}���%�-���Bƻ��3!���|\9�)/)��P��W�X����b���@��ͻEh7�!�1��٣���,�z+�IX]���b�^d�R�Ң�Xp<�4�?๺������ހ���<* U\�>��N=��n��3��5�����'����G�n�<�<f�T�8� �q)
�>U67�wA.�rߜ
ն�t���Ӗ���+����L��K?�j}f�[�	^�ث37�J�j��C��%��a�`�����7��!��n��G���zR�ZA�?'��:�����%�:u����N�b�x�L0fk���"�i�(p�c�`� �	mZ�y� ���$���Fq�Y�Jo�w��2w�r��jv�^EM�D2 ��l?����\��xk���Y�������jQ��;C��ki�Ƃ�h�y#�FAD�~���U�(�f�s�eF?���$>� ^UO�C�S5��b᜶>>�ޛe���F���<o�'{TQ�iTk�#lX������J����Uji��^�l��*'@�/���$�w�����C�*>��p\����;���pX�䤉(���>\t6��[���W��F�!�����A��ٷ�ݥ�z�!�}���S���5��i
�Z �n �fD%i��)��e�"g���{�<Z�]�Ԫ4�o7"���i;���$T�{����e_�Ft}��gö���ݽe;Fs���BL��� �� �Y�$X���+׌�_ud5����St�m�B�ܒ���ZId�!�W!�h��y������Ŗ��ּ\�Nr8/��rد�9k�#^�ǐ����K�}/��I�Az���?��C=�:���=މ�&y���#�j�q͐t�I�u��#e�XwT�CH��-z�S�R������������M,aw;B�p�OT�*���e_��,�,��.����Oq2���P4��`!$�|�Ơ*G"aM6����\r�޵��S��4"f��_�n��"1��;��QZS�阧�x���	��t�]�<��k[���it&���y�/ݪ�4Z��<ӹf-�(#����M��go��u�@�0�����ݓ��Ҏ�Mj���Is��WV�^�
�V��Vt��%i�8O<��b'�h?���܀�{���E�P;�I�E�nXn���0�%���OR�@|Ҿ?c���ف'�����x�PJNj_r��;(�?��W�5����L�oxW�y���\�UE�H�e�-W(���h!�O��������FЭ��]L��6���(��fd����\t��T3s�'+�mP�(���Ŭ�/�$~N���De6��;�'�m��%�@�0����t��*q%Z��vVD�r���H6�h�N��^�����#������ͤg���M�I��� ��y�h��C5�R�/=�jv�����}�����e-�,Dxb
��	��p|��7�=sXi�n�"*?�3�����2��J��ъ"f��&���/{�i�'<��q�Dj?���r���r~�ƣ���.������� �<^ӥ��+<|��U�/Jt�<��*����̤~�`4�5�z�+��{�չ.�&�W�E��Pf��^=�>웊d���������0��Kن[� o��qy�L�K�霵
c�Ѧ2Y`9<��y���J; �Ӛ��|��L��K4���V7����+ �V�/b��+P�-�aN~���@��I�=�Tg�OJ2~�r�@1�<���Q\�I�G5�����b\���Ỻt`���b��/£0Zl�8��1}fʱ�)��|;�ؒb��s�%0LE�p�9�cg�0=�"4+Vbc�5x|8z.aHY�t\����_�S.��j�)C��8��1,�5֖�~�(m6��w;P����
K�Az��H��|�i��<8O�#1`@7;����Z��堠F��D�u�������-�H⤔�Z4���V$�\�����$($<��7������\�jQd�l!Xg�'c��D�&���2��2`�F������n���W����("L�c��n��Ѿ���+�Q�,�gE3�Yf0��z�s̮=�ˋۆ����l׍K����b��A�����F�*����*}+!>5#?�k�N��%MpJ��P3{{8"klҭ�D�dd�*��`���~���A��"}�/��6L9��cMh�}3&[�P�a']�
��D�4$?�+Vylq�2���a,*���{��ܛ���J��EN���a�<�F�L�����_>J��_�<u �<��ςxk�X]���
���҈U%BO�[=���}�M*s�}�<�$�3��ks,����y�W�n��T;G�\��vD.�P*
��7�kƫ �����	+a�+a�������� Y@@�&`�I������Il�MGY�T�K�B�ϼy��T"��̓;�vҭ�GJ �����q T�`ȓ�PE5���:j���n�37�ԭD�9Ob��;��*H�[$6�o��mEK� �0DG�"�צFE��X�����(�\E���	.Y�Ӻ�w�US�a���u��x�Qغ�C�z��o�-j��Ւ�0�T��l���v��q�\�i*rS�Z�|�R��Dd�S���o~͔ �˅Z,�� �������{,�$\A���0�3���_Y��I|'�md��a#�wY�4I�?��ް�|�&�}b�3	O�/c�=a������v����3y�&�� �y�'��P2�8��ޖ�x�46��B"5�Ҧ+~�x���bo�6F����P&�7!�����(� �Ƃ)M��'���_%�,�5��J�A0kA��f*�Pj�}`����A���3�5�u�[L���� ��~v��BӧtJT���!"���X��|J��aH�<��d�����1E�؇Rq�$��F����s���B�pՉv�D���S�<��2���|k���{�ҝ���� �f�d��� %d��1��\A��8��H���+��S�]�;[2G������1؋}	 ���P7역K	��S�FNd�H�+Pk��T�8�?^NaëY�hH�`u�
��#�{�y�֧�C��u�1f�Y�J�gK`OK���l�F���T���k�è!]Ϝ&�����FU �hi��M���iD��b�ixu;�C��;�~�K�r��#�i�Y����w-34Fw+3,��Q%�z�ƌA�ݜa�ϋwCa���[)7�yK>C�tEJG`����B��>�m�D�Iu�1~:�C�gNON��GUΉKXQJ�#`rVc+GE:۷�N�w`F�8�K�#����Gx�/���O	bN<�z/Ǫv3=���2s�<m*�u�6�~Unpx$HV�OMRԖ����{�>wV�_;�<n���#�L>�#C�}���Y���DjP'�u��h�tʛ(� �:�]�76*~�1�Gk9�n2g&_d��[h����?u/�5p�o��
o_k��4�*}���������@B�TNd\cH���e�����K�/)����"r���b�T̔�G��sLP�I�nf����L;,�d/فB����\�h�)�&���N]�3�G0ݧa�����<�J�Ԥ��,xp��G�bu�bhp�c�D����H�3�h=�x�t���?�e�?V��P�|���s	�����e	DHT5��4�q�H4=��t~]��|�� J}��+��K*֒qeђ�$~D&� �M���U(z��dY+WJ��eR$ȃ��A���N[�b����ˢ�¦��|ШH�]�I@@w����߂�\�$�4�! }
n�8��=ڙ� ��2X,`ͱ�#�l�;�E����������Q1aO��b��~xwW���	K��y��������{߫����2FE�o�"�#�r�%�I�~$���M�s���G�z�ͼL��d$\�k���L ��D�WU�e*qg��3��!Z`+�i�����Uh5>���[��z\^3lx���Ze!�]�y�&����N���������i�IO�F�f���T��-a����a̕��>��֛f�2v�Q��·�&���A����uA�ğK��Ԏ�ZM�Z��n���y�_���pX��"��t���jǬ1}�d�1k�μqS1��G��@ьu�+�{î�YzϣAT��+���ʲMZ��;���!�ALg[��B�v�奄�^u�M�̆x㋂��)�vI|�y Q��BwC��DxI:�r�S�RJGhA�����	Wv}a��{A�5̥�3� ��>��)��)���|��^:�t���<�������I�-��E��8ܧD���mS��A`��׸Ä���Mo�H3�I�)���Zf�t�(}]�0��㑻_A��ͪH��j�[f&���^��w��T��.�˴�u�9�UD]��N�:�ҡ�$N���P4)��!� &����3Bp_��΁İ/>i��O�l������Mj	7;[�&Hej�%��n��/IM�0���ʹ�%� �1{`�P1��Lp�Z8ςzG��܅{Ϩ3zj�2
M.���Kė�<�}-^v�^�ܺ�B�;��}�We����[�4��4R��Т����㩏��J����9����NԻ�/�@@�Qo�&�i����}s���_t���]��� _ʞZ��_9B"}n���V���xg�Qk�i�&NV�4���g�

P!`��v�fi+ߑ�_y�9k�$�S��=��ߟ�{��X�]$�,�1[6d�p���	���R�BH��� �O�)�WE����e�O�"\�}���{���4H.<w���2�o���+@�~-N떼=wP6r1�C�ҏoC��7|t�-vD�Y ��yG5��9�d��ﲶTQ�~r`꣜�
[�<�3�_L�|Z)��a#���8.p��uX�{qqU�20D�ue�Bcs���b�T�I��{�q���B� n@��z/�_����n9�������1_G�LU�E���o52��U�	��TkHDy;��Hw܆�����G[p���׊XR�7��t��;JGz�t{����7&�~��L6j�p��8H��tOԡ��:�@{�1����Q���IDxw?s��G�#�SSe���U�a� 2��.;�SsWG���f��F$�	�BQ�g[ʩ@�����`�μ��D�+�I~`�6�Vv�TظE�w�9�s�UPw�k�ᅄ��Tvd���C6��*,�-�a��_mF�|�MiQ�	�~&:�"3 E�o^������ԇ����	��%wh0�v��U���δ���;����\��[���.���ڀ�w��-�z�� �����fF�Y�U����ʛ:J"�<[7��K|��5S�5ԛ�nCh��s !)ڵw���d��k{ٮv�C�2�k�����Vb�҂^�f�*��K�*Ji���!��9��%��������2��*�{��#q�"F܁����g�jն"��*[�#�M��^�����z�R�a) k�t�пX����ǎ��-����<���O�y���Gd�_v��D���:�ԥ����*����m��1�QmeuJe��0��4�w��y�U�	��6��k\��*/C�۞��NX�,2y����o�mP��F˘~vE�6{�B�S���"ƫ\v�X��{G�� �?Q�N]���U�z�4��m�xtF�,`L7 L��z�A����m��}�+�B=V0�z���4�������y0lI���n��dHT1�ey�]wS�}���E�Z��L�ɹB9E�~� ��»"��E7��x,����
�ܝ����U��Zu��1�p.5���R1�1,�6?��{M��2�|�=%��,O|��?k	o�/ET�Eld��q���@VRXv_{�\������q�Ԯ�� ��\����t�̔��.ۦ�LNDp:Z���+��*4�A����y��E�☑��ӟ�
�߮�]����F1���ZN�W���wh��sFuP���	+�#ª�Zd��s_{�����@��M
��mO��\�as��:��j�(TSR6j�߫��~�V�#���Ec���B6ޢ�2J[ ��>��7�e�0�6O@�!�d��0nX!�ʨ��Ng����1�4>;8�����84Z�gb��
�|�H�B�˨�b8� ��μR��G�	LN����_��n�.�[����+��Y�J��m����]��eg�ҧ.9=E5�����i�ȗޢku�3Y��;i���;�v�@2b<�������0�)�~�%G��0�Y����hר��Y_*���C@W�ѩ��c	u�SFr�wYb����o�o\��k�?�1�R���g�U��`Ղ��S���XBdF+d�O��VV{x"w�7��H��Fy@�x j�a�ʌ��AO"Gqr�郪����w-J3�%�Х�!E���������}��-�����s4;e>7RaE�B���qN`B�
�*}{>� a�<Ĳ�eW}��'��M�,�J=���2�-��M��}ʐK;J(.�`�*/8H[?I4{�	���ݥ���W;PUp�0C�3|s�}��c�D�;�%�Z�����D�+.h??�ATe��� �Y~�a��@���-���O�a��'
�aP�bd*��wcbN4�?� ���������
�\��6��N6���v��7�ʸ9��#� "�: n���1m�	4 G��c����'m�|7s���3�CT���r�ί��Ž�w��;�����}`�Q
��߁��>j �:�A]��W'f�c�J����/Q%�Mj��������tc�r��F.� �����Iǭqr�&��&�ܝ�W,�#zL9]������_�����S)��D�x�I��)�x$
[`w*N�� oG�wH_��\Q��b�Oi�ł�G��wi�v��`c{<q&��	
t�d�aM<��?p�n]�]�M���(�@A`zeЈC�p{4��0�(���k4��"�h��15u��>�i�x�����UTK�]3TO��Hr���}6p- \rxer ����G��I�8��+w���6wf����c/CTM}�}Y����9����f:d%�vA���%-���?,��b��Xy���(*������]�>%��M�C��9(X����Қ��6���_-S*��h!"0���^�&����4P��a=&&F<�R��������1v+ZA�� ��:i����Z���A����*0Al|:h@b�\YL$�F��2~�4��r��x�P�fi����@�*�8�$��'�U)F��Y�|9���MF�:��Q�������`a��e����[�1�����]�$�N2��P�?��M��-���&%]7QQ&Y_Zn��u�\��Ad�.���P)x�{U��L��B�,P,`�R�#���\q�E�n�M��'�eI|��e�Y.�h̠<�P{���ޘܕa���\��̈́W_�56�M��8��Pa(��eD�+ZP�H�E$�h�@wI�%�M���bc��f'�%�wT�����^h6}�:7��Q�8��(4���Y�Ԇ��J�Mgבy����o�E��c�_0����Ԃ���YU^Ֆvl�z�[���g|�"��s��C���R��_�Y|�5x�1+r�H�����x?<栴bW-��lf��G*�m�$��M>ٲ��EL����Ȼ̣�C���D&�3�S�^@��vHQ�_���$�{���7��2|Y�r�:R,꼬���>b�u3�r��X���"�u[�5�t �� 5�����2�}�2�E�ֽ�
��'�����!�?2��X������|��r�g�-+=��T���V���#ƅ)
ޑ]����	f�����۽#�(�͜�7iV�B��P�M:�x�a_�����$>�2�fJDz�~�6#�=E�y9vܧzZj���"'��V�v���� ��D
-���4�@&����*Y��v����3ꁅr�q/�Oy(N�Ͱ��I��t�握�Ih+������)��X^�G��|#4�la���n��ET�����g�D�`�D/!���)�z4jcƭ3�������{L��W&zVs�á]��Y^ָ��g-|1CD�w�SB+(O@�����4�ݶ֕MĿf5"�qm�{ㄸ�/�{RW�m"���Kf:���
�D��hO�y)@�tSM�]/�b9�8��]�Eg���X}��?���t����`R~(/�.���r
q���$��( ���j͆1gW��'g�>�r�E��2��A�ܶ�;��	���B�؆�+zR�����-�$wrtC�O�B�˲�n5(���"��p�dn�쁃x�<�z���b��Ǹ`Ò�����w&�/��v�+���ٶ����L`����<`�k��$#B�Ed��O|~�y�A�I��E/��65ɰ��8=x�J��([���15�v�a9Mk��0�P�~I���|�
���R��C �7߹�w���$j���Y0�>�W V2�bC��/P_x;4�G���bC�&hɢ�Xt�K��|��~K]K���XP����f('ڤ �D��w4�گQ���0��Ԅ����[j�J
ȵٷ!ā��'L�&��,8�p����):�F4�����e�sa�Z\�6���
9�78��'j��t��h\S�E�N��g�ٖ��12h>�Z���W��Uj)�)e�r�}�Wzx)�N�x<y��D��٤P pC�{�9�z_��+Ɔ򜢠t<ʴF��u=>cl�ysC�xV(����c�Z�z�3�f����4��j~8<�5>9���!�ِ~�&spWؓ/iS�����"!���
h�?�I(����� ��@�����_@T�C{����g�J��=��f�63M6�7F��#�N���8Q�4�0�
_��Q��םRg�g��X9Q��
�$Sdn�Y�#��op^G��;w��k齯  �6G\�����\��>H'�Q����C�jX��堣�b�4�������[]��/e�z���4aW�v���h2��B�>���"k���d��pgd)����ݪ�,�	"�rȩ5{ɴ�'���hMG�h�h��R�)a�8	vj)_t�R���t����p��#U��Dk���D�`�DX�� _%>����_/h&7f���d+�[Yԣ��(��������`�����o׊O�Y�)�߮^�E�M�����G .S��ZNV�|~��X&X�����@�e4��EIl��@���q��h����ah��k�:�^���|�q���EB� ������V��/Wy���$��\��jH�ܮ;�z~i�^���\_�c��n0��l%����̲ݠ�U��)����^t{+e$)�;�Vxq�j7��oDI� ��k�}�2&��A�7�9xh:��qmTV�c�T*�BV�)����)MM:���R���Rv�wsy�RΪ�n�6��<xy,;(�]����n��ɷRg��08�����ֱ�*������[j��@�����H8&8.�(/_�~����[9$X�'ꀵ^'e��C�R�w��2s�t���=�"�"��)lw=#A] �j֤��Y�z����xd����:��~9.�t
��Y�v��C�S��. ���ѻ�9�siW&q�>�.��X��#�(�Jh���-������6y�F�k[�����
��C5o�$��؋��"�4Z�>�:�$(]�p�����ȪN/O���K���;�o�7���XOj��9���ID��®�H��^�ن�Wa�t�%K�晨�=�2���8���	��VW�����J��Bֳ�R����1���hzS�u#�Ս;O� s�H����#"{�7�l}
�8��M�vP~V��ϧ�v@��P3�D�H
�\�Y�=`.x즢nX����>	��r��g���c�3�Rb��Ye$�U�-����	ܘ� �s3gT���$��!��B��7�o��b��ǆt&�mR���ޕ���~Z��W�c��2$䓎�F�o1�@�A�VS�=k�L1���HT��hA�ҥ�e��Ha��)'|�q˔�Z�?�j��V��v�>@�.`z�S�S��;R�g^=%�h#;F�#�M6{�N���6�����w7Zb��z4B������΅Քn-��$z"M��b�U� ���K���7�wʸ�ɒ���wG�|��-����@a��	N{��O� ��F�}?�Y�*Y�Itjy����dJ�[�.�%v�U�WϠ���/���%�	��W�ll��&�6�O�}j�1�h�)]��Fb�'ev�-�d�&�K���ΫN���w�f<�s�{�2,@k�@2E޴u�uNۿK΋��4*�MÜ�?Z�Y#�.�:�.��e��y�n�;u��C
�/��\� U�jFi��O?�ƃg�49H8���𮵐���#
ھI'�����e��R	���T�����X��y�Ӹ��7C�.]��f��S��>�Q��nv��Q(�Ew���9!����(%0Rm���Ӻ&#�D�-r����İ9������yVC�?O�4�m���ϔQ}Xɍ�\��BU��R\nf~�lf'�.9q� /�	���.������9/���فf�*�mz^w
{��s�ZV(�8"��f��W]*7x$��q1(���KH M���ԛ�N�6G\��"V����YZ@���ɘz.k���������'����\��&��Vϛ�0�%��92]�� ����aGGr|6��u����J4��#�bT��CZV�6c�/�5�a;D�����Ͱ�D�2�m���V��o�d� �zw1�J�GD����ia,�軯��0�˯��tHU�2�æ�2���8��KD��1� ���Q�\FƉo��Q j[xE}\��(�m�tV���R�'7�b;�!�?�x/�bk`$��6�w�����U��>l�t�LFHY8�!U%ζ�^���;g�z�iJ���t��1޾���yV=��!��k��p9�'�lG0�3 s��ʹ�-�,:�Zh�v���W�U�ai�#x`����	�L�=��bS�P;NC0/�)�!	">��Y�c�Z,�.Ğ��r��o�;�.�"�GU�>^N������	yU��3XL3�S��6
��mˤ���µ]LGe��0p�X��~�c�:'��A�{zͫ�9�D�0�~Q]TϫYņ`&�L��m�}�:��9�cJ�A%���	j*��]�},�d�����;�1����d5�����@.dלK/�nU%v��	�=�f9Uݶ �w/9g�����Cʝ/i!���Kgr&:@�LW�!R6�� 5t��nX�T�����˟��hiDfvZ�ԗ�*�>
��C���%5޽HI��QZ�RC�$��oe���g����T������y���r��%������5'tp�/��~���v����jv;*`�P��#�y�
/����_�.V���ȑ��_'SI�e���Ց�ѕy~�-�B���sȲ!��R�)<%u��!�HQK����t�b#Qe籣�A 쥽"���-$C���*ة����S��ϊo�΀9b���BfX>?��v4����ݴ�&"�>3�ǯ$��P��2,��	`�"��{���5G*����P)���Z�D�b0�e��(�a�,��J����T"Ϫ0��֥T@YU����xW�!G�>����{f8�U�����n"H�UR�{�� z=�u���Dm-1����e'?r��)z*yJ���g^!�%Ͷ�^Zd���i/���B��<�td$�W�\"��P��v3^�3k�ĵ��Tΐ�,0��EV7�U����Nإ7`):8�X��7Ө��HmA\bbX��Q�܆��}%v�X�䆄�ȇG�OWW&�}����mD�?�-Ĕ��*�~1)��X�0r�����^��~���*�RD�C�������1��l����d�\?YE>�F*�#]������X�j.'HLZώk���%�!�g��9t3>d��w��O��,oWI��?Sg��r�^}�[_DG1c:�/]��^��x�aMe�Or�QG0Ƽ��m��Χ[��k�R��n�h�N�r
P`�V&h�S�ܱs[��K�Q¸��%��E)!��,�i�<�խu��9�0��}����lp�n� �$�~��*'��N5e�m�1z�������t�>����`7	��!��>*VJV6P앸����9@XQ����Ts�� S���1t��#��1�	w��pf/�C�>�G&'��q����������NѾ��ځ�G�ۼ��C?�$y]�I�9`�4��(�\Bh��u4c>�A�/���cy���L���h��s�r��7����z��K�8�Y��<Ѝ����m4�ChEHȪ��kA�N2E3U%���nY{E��(�w��,'�ƫ[	ʙN×5��Pyk�8�]Tx�גQ��"���������MF�ZƴUλ�i��r��ǜ��'�z��%����jo��-��WvCr(�/O���$�TN�S3�.pG��nԚ�[���nwA�����HJ��^&���^�On&G�s�K̜
e�e#c����:T�4�/�-{�� ����T	
��o�2��������a��ߛ����!�Z����eR�>W:3^�����ɞ�U���������Zԧ�1\IP��J�8)t�#v' �M�;����G*�M4O�Y]U��D��@Y�/��~�;�q�$<c�B�yb�.���E��Ļ���ID�M �u�X������<��Q�q�ފ[]V����Z��J&�F�����%E��]'����7���{��<$r"�w|M�#}<��רZl���}�*W
�՗���T+����+,G��}���X�� /E|U���ƴ+��(:�	�﬷GF>N�b�O����[G�"fu���P�/�:4�}pέ������t�����5Ŀ��R��9��R�q��"رGIv��'�����Y�T,��V��mL �/��F��)�'�Zg�?�I������&x�h�>�M�m��E��<���I#�{zX���/�S�Ā(w t=���m�M�!�ڰ5��?�zRn*D�b S.\M������\��6�߁�U%^Տ�J�|B�� �Q�x�m���O��*��6Lf�k���V��ge�0���ܴR�u�0��c�2F�jo���H�f�����/�	�V�Ƹ`,�i}K������KA����pv��Qo�MzaP��zZ�}�"AJ�F�Mv	`}ĥ߃���Q�.PnX54v�NĘ�lW����ye��/����������"���d���$)�֥��d�N���?I�s�\d~ϖ8�(�{O��/�{�Ř�G[1t�w�y��z�[��8P��܍��B��h���K�<j+ ������P䬧����5Z�!��l���U꺵���M�|��5$��lیZ�~�`��k�X�>�$T⢗ĩ��̞��EC�R�xW˪B��o�SE(Ь�� ͤk�h]�TYLV�fY��ո`^�<iX�<����fYm���C (�b�zz�ԣ�����4�:-n.nL^e�m��WOT�zT1H�*v��n��L�W`"��]T_��3]C���3���Bʻ���+��9����p�I������:xg�&�Ĳ䈅\uZ#Vb� {6i�	8���"����*�=b�pMdVPK�G���Py8���Z/����8Ǧ`å��ׇ���`;�� 0�
XaJ���o�ͮ��?fl_є蝃6M>��\*qUyO^�@nL)�e&��b��i��R����{�P�x]'m� ݫ�_Ua�D��7 MB�Es!!�9��i� G)T#�	�?vf�8;i2ţ쩟@�S*l�ܳQ�䌪}z��)S~3Cn1���O���wxC�T,�!r��j�od}�r4g�~)[�%�`�J��1ܟp�Ut��~�Ɋ��;70����5Ww|w���g�?�Y)j�ȿ\A���$��`���_�!\�����d��N]��-��Z�<���׊R�KC��3��n����1DB���;ON=�����iv���!��׸塛�~���9j�k�-7&���Bѕnܹ��������2B-�2�og�=X�b�p��+�4I�'�,f+Vϵ!�	h�[�rְ#n���#�Y�Q8%������h�:��J�g He �}�˪#�L"��u'��o�>�ZW�\�P@1�U��{��nd���A�/�~��	W%Ϸd��l�dk	=��wC�!"�$�%�l/�f��
��<g�p(LWlz?��b�cmL�h��]k�\���|��+�̰]UQ5���8^���νJq�������̻��`n.��k���lr��˷>ą5�t��pPܨ�-����,أE���/��ݻ݇���5���0�,>���:\5��ծ!ĵ�E�7{�O��f(0�w���/��HV_Z �5Ͳ��@��ߞ�.yڥػ�Ѝ;��`�}���V�� ��(bffT�Q;�%w�C�y�V^�t_LC���G�{���j��3����T��a���	��Y�dH��g����NgC���5��R}Z5<�~\�ٮ�Ã��| �~�{�n�#q�"F�<!�� �^M�}�n4{�i}=[�8�϶����"�{'�U��<���%
�Q����(�|{s�Yx�A�Շy�ig�N�ɍ�)/�eSn	C����E��)��`���#�4�.F��g���K�l��Le5��ቂĶ�"���[8o�߷9~퍪��^XϩI�5S�~��_U�A{�E}΍C?��j�+��|CXJ�p=m�I9�;\�n�$Pg�%U1�C�:��c�fO��}��׍�<�ɴ��ҕ��0h8�����ċ�Ø�2���=9�.�[_�v���X_~8F�u�
xeq�UX:���g^���1���U�E�Mf�Bc}57��yo-�#4�]��7�[���A�TY�k��u�TW��1��G����6\�
�%e��o�4`�c����h#":D��t�۰T2���sSc���Q�8?[���%rd��
6NV��$��8�Zq)1:4A_�N0��a0�,B��o�N9��Ѿ��kA�<(�"ދM�
�_�\�bw�EtS:NHw�F�q��>?�+����{�L��]�[��N��i�eB��`PX:��t�⹫�m�S-�J���#�.ȣ�㝙�K|�(h2-�ח�l����w���*9G�P)ʔ�:Շ�G1�u���K�r�룢k�9:��|��������`�~�Q:D�O�j�;�� �!=�q���s�?�j�|��O��A-0�M	c&���QB��M�"�?E#�@m�S}5�SOŋ� �����c��ͷq�D�����$�_P8|	��NF���R�Nc�\��vo<'��7�u�OdI�ëwg>�����W<�1_���4��8��"l�z��g"I�ǲ�V�n�s�$�Ly��]��s��/�w���(�"� �`������p7
j.�x�6��p)��Z9�A��﯌�ԫ֗eM{�-�RLC$�Tax����s:�M��؈� �6��j���o<=2f�Vc����k}}��^H��s���Iz�H��e]w�ӑ���ſ��	H�>�U����1H3�����f�������%�J�.�{���=^�3�R��h���;mi�ͦB���:��v)�Gd�18®&8�|������G��~X��k��"�"_�n�6D����BZ�㜜�|��SJ��>мd^��b��2�;Ȑ'�t�s���h��;K�w��;�o z�ϲ��h��0wwD��Aw�1s�:�pS���`d��o����w�B!�'�hލEW[IZy���\�`���ݝ
E��x'2m.�/W��X���z�/sN,M�Tv��KC�@���p/�}��`_���Ϗ�}�R�-����,���
�޾< \I����*�Ə��p6sx�E�wz�· ֈ�A�X�EPfT�#��q�Cȿ�i=2/���v�d�$Z|�H%�6\�p�gY�,�WG�h��:�\�8�ud:���q���H���ߕ�K��tiZ�k$bַ+`�]¼�'~nhv�G�O���MU��Zݵ����=��9>Ni�\��p\/�x�u����L{x�TA���ִdU&�1�.��L�(�vN�'�ű�pr-�҆�OO��A�0/}L��Yg�1Њ߽�y��j���83�� x?@��C��̀SQYX���"���қ&q5��Nٶh���b��n#�K��Nԥ��+�=V�[;�I_�<�⏂e���$����w#s�@�����&��L��7�JL���&��v�*���F��| �>�Ҥ�E%7����7������-�����69�d7VT�/x�[�!n`����Q����2���,�``M1������c$�u���Z��c7'�wFi���AG�v�ko�ݙ#9����c�]�3=PQ短�e�̆���?F�7��sڤ��
:z�^����m=���V��}oD%9�S�xA͗�<�d�ԅ:7�ZK�{��eiZ���ct��DFHi�Ͻ�Wm�[���9�y�"H�WH<`Od6�M��7�¥vC�{���^�^J6@Ps���b�w'���U�ivj+����{V�Y@�Ɩ�Se�<�8a��ׄ\2Ji����ƣr[�Z�]��ЦLkĂ��@�x�3q㒛�+p�|	��||��92����J�鰵I�d,�>#�)�(M��
�V�tGY�;-\�:���+�'��8G%���2���$=ec����k$}��7�"��ƫ�,}��Q�3,c�>B��2�i7�U�K�ؔZ�o����p�ul��ExR�bŖ�ۊ��OJ7��gl�:�����$Rܞ*h�ވe;�GN��E����g%��|�`�"Xk
B��?������������"π�]?�z��O�km���ҝ1��P��%MU�+�mE�s¸қqv�7�8�u�;|4f�8y�,]�8�mx8����*B���eX���v1*�L|濨�f�#��x|�\U*��]O��Ь���[MX&ۂ7_�eS���a�?Z�G�_�Pi�\�����X�G��� ��s��X�o�6�Mz��������6f�����J;0BU�)���b[�@/�O-ǡ:�ꪚ46P�b���U;��#)�b�����XF��̭�m�y.���s�w��;�uj��V�Yh�뾴W\���)<�̢�u�ei�����茇��*8b�y�+Z�@2����&J�������|����ei<��u@�ålM��o��w��ݱ�#u|����Eϝ�G�1y�B�uC��j-�E;Pr���7��R;7��ڽ����ci1�!.��bg���q|����(�e�X�	q0<�{/��t��%��Uv۔�,���fA�N������RJ�@|��?�$<U��W�)�X0c� �h���J\��,[�$����Y�[�c�PT�b@���D=��z@����
'ߋR�1_����1J/�t���%�}&���m�b�Uđ�����Y�_n������kg\R��J�3����m�%�d�h���=J��������V��2��f��/�/�^�.G�O��/[���pM�	�6�=(�r�9�4�l�D%���Q����[uO�/�ϼ�mA�=�N����]Dw7!3ap罬a�wp�Rl����d�U���^j�0���Mpk��D��1%U��٠h�y�����I��]�%�ޟr��C_��μ8��Pj~|���x���7�t'���VFzpξH�H���f'g�?���$Ȍ�y)h@����JS�Q_�j喓B�����հM|l�	�V��O:h?������f%� :����"m���+{J���D��`�i�sIe]!2�+��;��(���z����H�U��cJU��m�'2VCWjƫx�-�
�L���Snp����!"8p�N��\�2ɻ\�)D�l�����А���d.�h�J~�l��ȮUm����/��g6C�M�iȩ;�É���oĩ;y3��eM�U�;��"o��½��Fh�ޕ3ug wڶ���T��+f� �q��c��[�ON����=F}-Vs��lp���x��U�ܩ�~|�x�G�š����~�<S�
	�/�阓�6����.D� ���=<V�u�p?�� �؞�����}d}O��J�jҒqK�����}a�`ͣS�.bϳ�>3F�gT�)�߸x�d�ȿ@��6��d�0�Y�����T ~�U��0��cK[�����Mu������.v[[H��~;.�/��4~�S��d<��9�(�O�Nw{ �-� 9��'>b�F�,���0���S�Mc6�3w!�mZ��us㥒��@�EO{ �H�K~�6���rg-������}�A��X���_�}�J$�!� �z���cl�Z�Ef�����E�+�V����N��Ђ��;��9�ֿ��r.����`��$P�g���y���?��E��eY�g�@�wSJH����G�0�^N;;�Fj����k0��/��}�8e�RrS+��A���G$k�� �פ4��l�]F�r��5�c���,�C�c�6�'"#s*Β��h2m���>����r��Y&������ie��[1 ��0���Ȭ���DW���ź(}t� ��
�P'�M�qa��WU^9��XĄ��G��>���QJBwD%�n��QM0���+:����bv	�����À�> '�������8��fJ�q{�t,���@��f���Is����$�@�>�G�~38�q05��y+k������
�m�T��se�gx6��9�oJ��+Tg�oH��Ϥ��/^G�)UX%�'����iR�Q6f���.�5-�q+��y ��c�����"-P?@h�~�;'��cI�wQ�g��Q⏵K$��3���Ck��GL�����	x9��n�QNE��׃m�i�I0V]�z���@�P17R��?���8`Z��~�8�2M��dF��H�K�@�K6�j�1�DM�`�yuC\Fn{�wfZ�|�!�f�c��v�7F�X�Ϻ�?�n�Ċ�=a`��	�c��FB�V�4�%�j�]ȝ�hT;���I���?v�ώ�^�6�V��R��� �%ix�>�|�m��Rj=�B�����|�(XB�ά���?��'-�%>�����Ǧ��L;(l���\�Jf+��G����/��V��vw������Cx��kX=^^��<ƞ-8�}�Q}�]i�22���2eU�;�M��;�4�[�CJ�:�[j�.��>���~�������vq�d}�Y���j�W.���u�Xt��-j��+��ݔ]Ñ�V��)=ĭ�K�B�C���Ie�ڟ��u��f�`u�k�<���RV�xgɄ��%J~�G8��c���i�v�!<�_׆��`�d���
,�5>�Y��}��_)���犽�,ndB�dͼ0:幂�x��%�W����d�ۏ/?ٲ��%��j;v~9q��`;�����S�:@C��b)*��NL[K���T��0�9Ld���۳�}Œ�]V�UѠ��s�-@6�P��2$��4NŜ���ߤ.sߍ��C��Q�؊�C#Ρ���{P����||������Ս��H+�"D|���ͽ^:f�K���e`�7�
_	rW 㜽����m�5اw��C\V���ԱyU�D�w�}���K;������(.k��(K�Q/�5(Q��_V_�աg_d��.�[�FI������J�h�6o�}i�zx�xf��Z7�nL�@q��ɷ�K�!�l��H���RL�`v�V��P���za��*�R:f���ēQw�&~�P�mcf��!J9�ax�d2���t
(L
=T��]h�*X#�
�IZrI����8+ǒx�X�nƜ3�`EZ�K�6Ξ�¸ĽGA�̩�Ť5���t���m�EK�؀`�Z6H6�G�
zg0kނj�;yO[�[`����^�������:I��_��,����/B?�76ȇ	���u.��Xe��9�8���ڠ��^I��09�݉!]L��5Ũ���Z i����H<y��)[�9�x��smR�>s�+D	����A��R�s��+攊Xv��ua��ZQ�yɠ�/�=�ؓ=�c������^�ހV�-z�>���������������d�b���So&�p��F�J%.��˝��g� *�q�P�r�*/{�����N��XTK���e;0�<���Pv�g���R�Y�U.�>ޡ���0�6}LiW�)P��Hɺp��0��˶��y���o⸟���B�#�oL�=��2������C5 ��ڶ�+��� ��nrB���4QB�'a�����d���;y}��g��(t�r[��3��^ʿD�(D]W�r��,x^�Y����&��䍐�ϳX�|z��~�l-��R��\�MDN����@�X]cJ�eC�����brܷ��[���m�\�������J�2�v��WK再�*O<�?� �J]��rX��)�#�3i�����ϱз$ע�P9�Ғ[}��(�nr�p~�^Z�6QU�^�;	T�����rM,�aU�aZ7W�F���M���h������yM�
܎�����FJ�+rFD���D�Mi�c�@I�~3��З|�BU�[N��y ���9�#�\��&���S�$��,0��e?ACX�C;� �T̥-�	�w���q��T7�K����<��'�]Fu\ۯ��FM!�Dy��M����ee9%fCʋ�fl��ى�N�����![G-ht@�	�Fʞ�Ȣ�pAD��y� 7*̮MP���O�s.����X241�Y;��0p\ux�1�u��~8<Ȧy��r!d&��Dv�.	�O��T7�L��B,�RS�{���a�T�|�B�år���q_l�6HA��d?o���;fX�bs�[�	j�Q�v+f�Y�׋c����+� �;<�c��R��VI	�]Y�%� 0��P�Oo;��]f�B
NZ�{��9b��W�hI�c�xL�}+[��޵�C��T��>=�#�s���8��pϓ�1�F���Ą�D4����5H�0b�5�S� ,P)xn8��g�׭t����̜�3�A�p�e�J�THS�b��~�`���L��^�1��I���@تw���m����f���������T
L����?T{_�`˅8s{J�A��eO#]�J�c�0F����;k!�g+Z{̈́h8&A9'���Q�Cf�E�]C��j�!����������Se8�:��1�y�lf��9����/�za�ۑ���:���` �7��$��y��R�qF?kҸ��c���>+y� �h~�L�ni'r�wϸ0�Cfd�x�:�%yܕuq��Ԧu��Cҩ�Ħ��> ��s� ���KB�X	`顑s�a�Ң��j��Q¿oq�����%��UnT�8�E�/*3x]�^b�v�m�o��㧥g%�b�\�Uߞy�ɾ�]���Ǫ�gط��;����-���N�νCL:1蔘�=�@#+��ɑ�(2e�og��q�-���ñg�U�
��>}&�W�>Ǽ-�<m�������.G��hA��u0��Ǆ</A�5�`�o�mhl}sY�O"Z��U��F��A�r>fm���b���ɁB� '!/�2N�e��W����Ki��L��$w��'�%���0vL�L,�(�Y��;�"5?T�(��/���0l�����ID����I�9��Y�?�e僋�f�@���U�eo�U�u(/�DvV^[�)��_#ز�m/�#n���S�HK��4�fN<��w�ͩ�t<�E#��4W��A�(*�9n����ϸ�֐��9�i�J�K�	$;%�����i��F�"��E 3�c��"'O�ɿ�H�Sv�xws� ��!5.�c�u˸0��p���"P�f"<VQ��55�SD��j�v�3�ﶛ)�����lA.��9�J��}z���'����Qda��8�3���@�h�����f,1�~�Rd!�:�a����0�W���/���dF���V
.]O|Bi���;���@Ƥ�� ĥK�n�T��	��#P�'��G�.�g��3��n�)]c���Mf��/t��N3Bo��Uir��
e��dL(Tg�RrG nٶ����@��i��E��1X|M��H�:�z��/�f2��Xj�~����%ej�A�4�	��+"ܗ�Q:M\�;��L�S��q]�G�2�F�0�;LA̗��~dr�6�ݫ�\D�/�9����iAUŦ�ƨ�[�j�C����^�7�y�9�^b�t�#�q7�n��R�8�<ɺ�0��+��߹��r�Ω� 8������F33?���E�JR�@Tf�⯧�%�k	�X3M�aHͲ<n�6k�a@�����0Ǔ����v&���2�{UZj.3v���ԝ����G�J��J�	�Ɩ.�L�c��tUʵN�k�;��)�vk�5��9�Ѡ���~���8�Y�!�o�t��~�=t�D_-T�$]^@���B	��j�"��k�g�/���M+�h"��"f u~���.�*E�z��!���2T�jmۈ����ZS��Q_E!A|C}L�v��o2ue��.�`���-A�A~��ħ3�����l�o$�XU � D���h��MHY�č�H�PyB?xDD�G2�ݻ򆑧dy�C��*@i��3�9�,po����57��o�FR<�v�촋�c�\�m�v�mV���-��
�i鿟U��њ~���o�@<bN�l5Y�@�\�$�������3���CY1��}���u�J`�<��oH{ė.��D�۽J��%T�	��Ka5�{��{h6�>0T#8�-H_��{Y���k�-#��qƭ�#� �/�J��{���e�/f� ��`�:��z��u(Q�$�HU��8w�$q�<[��(y��wd+��һ*uw$�E���Y�1P����ڠ�� �E$J[Aw�D=��/�b~�Q��C�i�����ˏ��?��)r@dx�'��u/X�����I��ѰP��c.E�o	m��܀D��t��,uqx��tó�P|���U/�Z�4�q��d��I�f�z��VO�:��,���V�96Q�4�ѧ�|_H۬�<W�ːtæv+��أe��?���e�뫦�����H�+!X�N�F{=Xu|5`�����D#}�Y��ђAJ/�`b�ѧؙ�l�Ѕ����]����Π�I�l��?��v1�/����g�l(ia�S����OS#Z��Q��z�۳4���y�6�7W���E�Z�E�8��|6{�xT��p�/@?j��������S�Ի�	�U ��iT��ʼ��I}�������>40�O�e�&,��Z١�1Vcy��a�昪G��Q�HL%�֑h��@ͧ$�{��{O��eq$�A/��U3FW����r	��M���M��l5b��T�h=;�줡ʑ;�|���0m�����t:���a,@d��4P���鷊G��k�`����qs&i�Z�q�x�h�a��u�^bt�FW�x�	+U'��P������[!_/&;�r�<�3��ݎ"=<�������D��|XFlD��4��SmR>�y��mm�t�<N��tnXb�1���Ba�Utm�@�WG�B�90Z���,�V�ЗJ�g��^�l�f_�!�~,Ѽ�q+~��jAU�*�y��W,�i��Y=n >
��x+����#��۵�,n��jra��!N��e�u��WL��:�*�? D06c�hI>�!�5�m:y�����a�σ�Ba���vP��� Tլf�͎(��N��^46����_�{i�I]����M;�G·{�vɘ��V���z���÷��X����s�cG�	���	].���ڵ��	�w�a r�F�;���mL��:5/�kF�����XeQv��r7����%��[�rr�N�萍�Ᶎ1���������I��Ե+L��#ok��&����s�zǴ�|ёRQ>X�Kr=�r�����My����*���B{�ZjӢ�;k\Kݐp�k�tC}�p��%�K
��Z�,�S�U�{8���4*�d�܂�ڮ�}�������,T Z�������eAŢ�������YK���A0�tH���g%�ɦ��.R��}�b,��8���ЬF���fϣ�6ΨN��EϠ��U��������TL�x�e��m�/=Qbr���	Jlz.,�X��#��U
_���S�st��?��/U��C� '$ug�`���8A��裆���χ��I�5�R6:�`��aHE��[���P�@q?u����&Sv�~H�$��
�sC���BE�)g�B��:��J캺�����>d��)e�:V�J�Tm�R�9 x������Ȇ�7���A�k�3n���)g0r!��� O��|f��@���I9w�Ѡ��r��?�� ��o����}����������3�)�	�\ô�Ue���j�)W���L��ONlѱ�N	�E�E�
��Uo��I;�͒���s�d�><�����˯��NN��Ѝ��YZ p�� �Ga�+�0�>J���q�3����x�����rS���Q#}!��k�[֓LēL樫}^�$���P�P�e����d,[��Ѵ��c���҄��E3��iq�jϳ����hWr ��ͥ\T�ѩ}�[O�NƲ�Z��Q�����!� '�Hϧ֜����_�u�E�mb�K���dy}�e?.O�~%[��Pau�{�?�E*�4�ǈ����"��]�Ki��Mq(P�DXPC#{�Ay�8'����f�ю�rNLS\/Yk��r1hC�9��1[����M��+q�,���3H��H�:#�Cm�.���N�Ý�"E;ԤWꚉ�^[�rI*H*��v0g�u���[g�Jo��������_�5b$2�>�T~��˥�^���[,��[�-��q���ӯʹA�ISZ��4N� �ZR�%gZL���?'�dI�e�~�` D��`N�AP��o)�H9�q��'��?�L�v��b6�f�ݬq%����j�6"CՁ��r��7)�)qa��x1e8���@]�ո*���<�φ���:� ��*2(�^.�.a����*���s[��qE���V�_�_cr��]���x�>�l�L�����������'�x �K"̥��������薦�4��1E�`���8bA\�z��y���!��vי��rR���;��`2nP��,c�u9/m���0H��zJ�Y�h�'PGj�BY�'`���,ZW���fTeϵ%+^'tM_��E9�GG����
��2Z4}$�j��FN=K��wz�7C
�1a��]!̀��d`��*�w����z�L�|<�<ޜV�$���8�3rb���c�t|�����^M�?}�ܱQگ��Ok���܄����*�k	�]�N	D��}7	p�܆9Ax���Y�����X?��ǲ�y���6�} 7U�\ �=����cL�d[e
\P���3����dc�8���p�8�4`Y9�-���C�{�_�w�'����Z4��g�n�������Ȳ��a4����b���ι���4 �߅a�����U<��h�߯H'?��;-�.n|M�`�.���glm�>"/]5!�CV�O�X������c��!a��=MZ�V���T���a_#r�̩&�Ԣd��P�oE��U��c\
Xv��;3��_U��S�r�v�T��	"oV����gWO���VD��3�{��װ��ܻE�������CS�[���w_�.���w5���НSb&���к×��r!���z(���@�]���[�a%&��,`!�#�e��sd��t������f����RS����y!<�!��۶J�hAx�;y�B�5���i8<"���i��U����[H�,�Q�g�݈KKn������"��+$���0��隭�@}}Ns���Պ�T�T;�c��@a�� �B0�����Y���X�c(���9j�cVd��"���.�y��l�I��ZY���u�{ؿ� S0������O�2k~��fdW�ݿԞp�C'X��-�u@�Ȑr�/y/��>�I���w��$YaI4���$�ݐSc@��v��;N3�d�\�hN�[�5V�g�����"k�J����8ީߪ���n|�L�)����-�����IZ�O'�?�P�w��(Ӕ{�P�y]ye���H?�g���v����E�\��~۰l���@� ���|��Seȋu�-t�j�Юv�qd��jxQ��Ȟx��"]O���4�yAҺ���8%�7�{�5�7�}�ܖ%�����`5v����,[��
��&�ƋC�5��T���	͖�hx�|�*	̠�TrY�pi���.�wଥ�k]��O��m�(���x?����"�գ,��]T�^ii�/�!2�Tw�Ыŭ� �)F!�J�{1�4��C�w���u�C!�;\N8��Cx��Ú� v�8���А�9츿���W�o��%��M�#C�m�#&�K��]P,Bc��}ӽfg;!N݈�qI��a<������Fb��:8ͣgdm�S�]:���^w�RE[���T��$vi�G�.�βO�q�m�h���a���҆\�ry�?�r	nC;��J����E�#��V��<Z���o�!Ꝿ�`\i_v7������qwջe������'���?�׃�|�-�E�p�)�t	7yҫ�L��j`�,$��e�WY_(���g�)�X*�ׂ�^�r[p�'d>Y��������qi�R�˕z�1�y�/����mYAuN��G 5���ۆi
8J���z���C��e(�{��߸N��.Ll�����P�wd��c��n7$��$DnN�j�B�Ξ}�vAm��pD���5�R5~ƈ|V4��7�cM�Z��Y���@ߤ|<�
Ѽy���p�]t(����z�g�IĦi0��MFZ8��&���E}%B8�V'�j9e%Iϑ��'4'o�Yf�R>Uѷ,�P��ql��Z�j �]��Eեg���i��tE��H�J�%��:ʨ�@����M
�cTX�I+���Aj����"$��4�������d.G��]7�x�ѣ��q>�3���d39Z�(F&�a�}��'���&����/3���9p.ά8��	j��)�H�؟�m1M��_R��tjEj��c
#+@Aۑs���B�;�a9qT�)����-?����$�lz��aw"�95���C�6�d�<%��!A�4aB]����gʞ���A��ҳ���γq��f�%oL����F�s��$༢E�Z�[��b:�Bn����>��՜"ڊ���4����ЍZ���d�s�3���Q��RUip�jz�{x[6'�����&�����3�B��ŋƬ.�.��%��M��GsZ�o�^������W
�[2NKi��cso%��C�`�7Eiԭo�5�����^����Dx!w]�� ��apgu?��� EĬZ�M,���QI�HY7x0,��a�(=JC�SA�l?ռ޶NS���ɩ����t�ʼ��y�,��},U�{5�j��"/� ��j��7ON�4�I#O�dpR��v�3���d'@�W�I����֠��}�� ,2ڣ�BO�o�}��Պ��:�ɞ�7ǭxXI��F�y1`��I�����#�ύr��4e��*�&u��x?��Ϩ��N�V_��ۤ䬐^/"/̾чk���t��j��p(
2*���e�q3x��$��	3	��Z��$����Ě-�P��ܬ5@Ӵ���؈V���� 5��~�d��2������k���'���-�eEk��0�s�g��	~6���nm3��X�R��F\a�}�+��$&KWVf�`N((�����j�����L{/�b���wQU�љ �x��V)�_�L�n6jn��d/�Ľ�2(��3�u?'1�f���V�@�oI�!<o&��
� ;��h�N�(=;18�m�j��C��!K2Æ�-��K���7��%\\��CH-���U'8�)�
�ʤ?m�����v�(��v&tw����|��/%ù]@k������&��tl��qd{;Fv6�Gxg����y\�	c�G+�j!�c���u��P擈䨜����k�F�jO�!������KR5�zA>g���0�*j]sϒ��t��?6e��Q�ɦ%�N���s�z��#\�P���r��Z����k���'��	Y��a�D"�i �=1�^\�լs���nVR�O��h �a�ڕd�â8ڟ0xZ#B�]�D���T�>f��%�	4��},O�dџY�Y"�?�GV]�3J  PQ��Z�dղ�0M����4�i���s�2��ՠN�j�ݛ��ynC~֞�!^E����p�"��T���n�3"�dR�}�VB��ΘL�$s:(�Ф��>M?�G �%yXi=�g��򟗭��W;�ik�;e���k��s>����pH;�&��%9�D �Yj�<���y`�!q�j����n�r��;��'!�5�	�oQ@)�8Q�bi�>�:W敵tF�x_��-�D��3pfG��0��zol��?X}2�:����Ws�'�=�X�����B��:�O�ϵ=�rӯ-M)�d�I5a�|�ѩ_��_WP�[wH�|���g�U	8W�hdp@�����ji8S�З.�b��5��Bl�M:\|$0�/g�y>���b���L�5F�n���v�뒬�*���p:ǈ��/����CjqgL� �_fI����:��f��ec5J�����,o}����?US,�b[�ї��q��S���D�	mM��3�O��}y�X� ��m��_"Ꮜ]w�<	��-�@�,�0���w�)�dh�) 7�Y�z��0>��WM��	����'1�[�Y���ֲD��N�ޡ��*���\ -���Z�y���Yh�A�kM}zf��M�LO�8��ѝ�ٰk��Md6�Û��j�X}rI�=	f^��4�	<��yg��z�F���`���$�mZW���Y�/����M9����!�LJ��/�H+�*�i�̽�B$��u���s�m�XY�7�x��*]c����;��ʮ���=K�H5����B�����Ͷf�`��wf#�
����H�0��>��I1{騰�ӝ¸�;P����Yz��8kp1o�~Q�����+T���*5�K�c��koj���!��f�nn�!�|֝��Hj����?I��zz�ʱI���[H�c�\IVl{V�|4�%��UIGB,$� ��fx��%�����E�[du�Ù���w��
��t�1M��	� h�ф��q`�� d�T'/��迷Y�?�cE��+�ֳy����C�?j���W���w%aS��	�6J�҂�Α�t)1E�qT��Dޟ��'*6PYG�Ǵ��W {
��A.��߃�>@��`�cx�裢���q��[8��oZ��_2�L��	l 6]ǊS��:��f���<𻙿-��"e�<O9���0� j��d$���ၽ�����i��Ʌ?���&����]!P�Q��<QJ�'"����;�.���I/�L�tߐ���"xY�5v�6��@�N�>@`��B��U^
^ on��+ dWx�~�����;��ab�i���xc��ߙ=�i�6�� |a���#yC��G+�]:Vl���mF��^�ֆ��/[��m��I�L61�E��z:� ��hr�ٶB�37��-ID�?�B4��Q�wHx���o9��@$���#G�����aՀ�G�%/
�]�_ �}�Z�G�i��qh��X��E$�:˦s�f�1J���6��>y�&Y��6W���~͗i\{{"~�kiSb?�9�P"6�g-I����<��h��Ʒ�
����i
���>M�Ҍ����85�_F��Q���9��i�}G��(�#��~����&!B*��<��<�q1���;'?�Ԑ���*KS�	ɧp���]u��v�dL�~狌�Z�)ځ�����$�Ƌ�^6/�3�9�*� �x1��IYD��y�o�U�C�+��lS�e���9�3WU�L
L�j�S���d�Oj�r�&�K��֚߳2!����٪9�蛊	�w�	�tJ�$_�c��+�R&��*�n�Q9��E�C0lSn8��哌 -�
"R����P�d/�ʭ0������\�J0hx���� :O���G�T�\D�Bk�2����=^lX������@r5=�D���L�[��͙]jz�	����y�^/���rm-�* �����N�P4�|���舄�~
 �D���|6�����m����}�$F�J��:����(l#c����ɝ�^�9���ǬA�� ��l,�0
�;� `I4�z�"�1��K�e��D�mLO�NRh�����h���'K	�W�d�VYWuz�^h�g9}��1~Il��f^�/o��U�������p�Tg5����8�����v�l*/���a�Y!Y�j�<�R/�'B1�G���ך�X{)���J)�3���$Y]��^ڙb���(2�K?T�}�"�ok��
���5g����|���l8A���Ģd�B5A\��}�� Ww�BԷ�����j4X_�*�a�<"��6���N��}q�s�.,���DT��8kI��� ǚ[��ʆ�x���1v�0�\�ѯ��P��z��"��N�vz4�n�[�������'X�X�b�֞����N��ˣ�T�'z�w�p�6�#LE��,O�P�K�
0b�G2ږ���Z�0O��x�yu���g$X8�!z�F�$��w�� ��%=����=��nv���+Q����[�S�H1��ִ�� 8���FO6���w�M�*�'�2Pkdщ�B����rT��N�&[�m�����v	��*�� ���X�ű+�� Б'A��d�8�������@f���b��7�
V	g#��#��s����}٤TC݇Rȟ?�rb�7��pnQ\H���pzS�/@H$N*�C�?Pa8
[�6����$�L
:������G��~|V�4�����V2� 9v��3Z�	<��2Z������������3y93�TIh|�m(�&�V�8�3�w�?��-������ʬV+Mv�y�c�����{��$ԆN�'�Y�U���s�ĸy\�e3���� e�]�x�d{��&q9��~��\��E �
���b|S��L[�g��O/N�X��s8��Z睑���a|�\�j�)�U͉x=��.e�b����Ņk��9�����(/���,<M��E4�7{'���}���ӟ�?%&��m��ÁN�!�Fl]���=����C�!D��	.*$��(��p����vU�ڰ�{�yxt�}�����3�[<�/��Z������jҥM����4�%�ǌy]W������1m��7��s����Q����ANk4s-�E+�Ѱ����_9�(Տ%�;��X���C�(�q�A5�S�5l��NLe��"MKҴ�nc�'"��9�[F�sG3hs�1�u݋�LZM��n4�li��pu�E����V	�N0���H;�H�,�UC�pR��lj�� Ҙ�1o	oK����� �|�R�����>Y���}mcm�J�gy��D��:]�Rt�Y\���Px���c}��4ɉ�~LVXb%�-1v·I}]r-I�o��Yq-_����t+��tN�֟��W|�INv��I�wZ��\k�rħ�}��(�sO*�>Z0�>[N��GCs�S�5����#^�D��zn����_�����&���Ҧ};� Ŏ���W�1����$�.Fk��O�����t�!���̆[�<��b~GJ��K"sӕ���M���w���߭�P��\����x�k@��X>�/��*;2��ji6r8�?(6R����P�){�ʡ���!�-Y�O�z�Q�m�|����q�Xi��l�no7�5�=�r�\�ƕǦ)����ƣ޿�1����8�F�a��U˔D��x^�ɩ��?��E���$�*�ٛ�vM��י0y��A>V-����젭��Z�q�Săw|)6>�U�Ohx��L`�5b�%�!q���'چH�M�;픟B�J�AMY�H�X��gsK�`�/��K搥�=/)r���`�N�K���GYZ�Aw�� i���=��Xd�M䮸��T/����EQ