��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�۞����h��wdIv��t�o���G�QM������VrJ���
Vt�%[
2���w�c�W���p���NB4�q��7��f�`�{�#��Tg���'�?w����E�?_A,��6v�t�:q��)���[nI�D^��ɵ�.��r!��(���Ym�? �{��'�U�*�>ԙ��(�*�0�Q�M��V���H���^��_��.��tv�c�އ��.����F�D��P��լ�MI�0�~$���'p2�Q$Ǯw��C��Hj
Qzm���f�=���
h��ث3�5�A4�[Zi��9&=�%��\N�<>���4|yǮ׳-�t���Sh����
^<������6�>޳�Qb�2�b;�����O{X����ͥc���h������d1x|^�2����e��b�]O�ڼ�Q"-[U��ްUެ-�[l�	.��@��8Vm��XJ⨍y���`�*!��k'�o;�ۖp����׀,Cm���Z˟)�~֯��-�\�iFk���w�r�׼�x%��Y�Z�s1/n�YXm�_���#���Q$�������3�ח�vd����ݔ)rБ�cv��se=����̏�G��z��1_�>n�Ho�k���3��]�����h/Dex��s^ر�1�ԑ���ݐZe�`u�����jVjjD�\1)N�&�ˍ�$�;ZN4PY���޾��r���J�Q�^%�V:��2��,�l��H��1ٕ�l! ��At�B�vd�5�U$n���+ʆ2�����	Vb��s�h�v� ���kT�37V��57���U΀�􎤥���r�[�XHd�~8c2��8��b�}�es��~Ǻ�$\����!T���� ����p�iO	�	����F��-�2�k����O`��[ݘ��]�2X6���L�X�,	�� �`��	�y{7?©]�L�3���(Sg�{�K�A�ilxф�|K��,.}�G�*���6��by��3!n7�*L �Xkw��g����� ��VE
f�c �$q\�^W=$o�28a������e�y�1���(���Y�{O��ҳj��x�3	��'wR�%�	^�&޴ߠ�aͪ��*,�����rY��y
{�.p$�(�B��oW��أxH��Vֺg6h�X]�={|q�W���9U?=�����hXk{i��;��/)�S) �q�I��c�1�i�|]�O����b~
��%h�iۚ/�vWY�0D�p��#�G��J�h��*���8 ���Ń����������>i`���E=�����k=�0������Ε�dMg��,C",�	X�&�M���@�Q�L}1��&�e�}���ȅ��.��D(m���� /������1��V yL��)'�w�Y\�`"~;؄DD�~��p�_� a1�ib�Z[�s�_�y��[���*��=�yp�m�@f]1jJ���:���,�̝D�\z�9�r��t?�,q��O�}wW�Uo�V�A��@���1�kM)�$5Bܖ�׺�]Bw�����~`��(̬חjM/�-���
��e�2oRȳy	�NHzަ��B�=&2:~��� �<�o�UOnbV��YN3l�mt�~� ��0w�~����J� VJͫv1�O#$��+��4K���X<��(B1�q����ح��j�-�|:၁���RO4�<�`e��Jtmq����7ؚ��b�u�cMI�f*Er���3�}-�t�ճ�+|����A�ɢ�nO}��)����D��;a6�u�!O~Q���~,�Pmq�}�>��G���\h���0�� ���[����/0=�f.�Bp�p�Yg�No)�+���̻��V6_�X��:�,*��)<C�޸�p 'L�Ϊ�L7���ײ�ťغ�2a`O��W�K	����pĥ��d�[]�ϸ�\�-��>��2��6�,���X�(��%}�҃>iu�L��Oz4�9`X��\�%<=S�DL�>IUԧ{��\��_�5����V&8�?{5:�g�o#��	Ju"��Y�4�|��RIL�[�M�	"��Ɨm�sVj�i���5�z��wb����ǁ~َ���w�4Ć�^hi�x�s��{���y�gAA,�K�S�*[��R�