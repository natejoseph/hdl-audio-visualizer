��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��Td��dxC��!k�h,�_�p �]�¤���M��<���BJR~	��FdcB�t�J_�7R�x���F��a��ƪ�~��C9 D���˕VF�H��f��n��(f�Ek���o��"� �&"3=��*��B
y\��3�vC̟>uF��X?JR�����ҍ?	s=E���"k��"L=����U)ݪM ��>��z��m1a�T+���6�4��zƼY!*��W�3->���!�՛�r�,���@�'���\��У)iC�cTjϔf���oֶ�.��+O[��=N�B��O;�|���`W�;eq�)O�38�/T�vޥ�[J]K�S{ �S%2�'{�`9�g��=嵵�za��K"W�<�_R�|i9��W�o��u����4�����(�GZ!�|#l�"�ۣ�q�㣤;��)WWT7��(�a�{gp���1�[�î�g�}$�`uL!��#�y�dm,̠6����)٥w��M4����=�ź� �i�-"��nF��-������@zr��.&t���Wz>�%S��R��AN�c,j,��ei��"�����C�e6�~o�%��=.S�M;��7N?\�Z���\�H���"Wv������>�s�"��ҿ�6	��5�_n�}H�W� l4�8W�B��:�]'�c`G��F^�g�a��j��t�}l��5ҍF��ƜD� ��sܘ���c=w�z�x��2�_�*�����{����"����Uh\��#{��%Q�
G'?ךptt}��Fmg�i�r�᠔�o��9�Ąo������2H�q���ᵜ�f֨��F�;�g���5�5(Z�1֗���j���KO����9"�k<��b �V��adU[���j	�m�-�ח��s5||��*��L��	�+�]�*0��������
M�'،�����K�^?<^���UP�� �zR�.�ե���/��]�*�Q��ɐ��:�6lu|�Ơ�>;d�+M�����ĥ>r�?+���$B\���m���-�W^f�j_�=�<A�ȱqD?�����8�]��������_��ݦ�;5��v��/��*����4��ˇˮB]��*F�&�]EZ��U|D�8vV�̫�x��@j���&�����bwu�_u"��@�����3�P�����iX���	�#c�m����.ja�%�Y;ܹp�j5M�.���;L�ox��ǔw^ǲN��W�8iE�B���2�]SK��^/J
���PE��|�$I�*��1���W��.� �I��T��լ���P������(�3=�ax��/*I3Q��ԔA�x�i������bS>��+�hh�N��t51w{�X˾΍mB������KQ�lگ.�fC��0@WJ���w�(��3�Rj�Z턀� e�Q�dH!�H�bRO�r�����Z�l��I���`���L��f/���ތ�,>6�n?�g8�X*7�T	�V<�T�2�k0%�\m�S���q��Q7��("d��{�ڒ>�\#4h��kC9��n����uJ�=fh+
s
A~�O��}�֏�31��V�������<���g�Z�G�n��8����oO�P�%k�J���,�p+�Io��@����΅���_ŀ�e蔂Ҧ���'eį&&���H�d�ߘ��w�X��a8<����x!h��8�M
�:S��5<�S��_��f¤*�����\�*T�`}�d�:�̷���@�^bZ��q*r�!�e�#R�Y�ᔙ~���fX��x����۠ﬧ`�Еn ���W��V�tۅ������<;qCV/d�z���~�
i�y������ iQ�l��#K��g��C ���+���X>����U�N�2�:"헳�
1g�H�g���Nج�f�N��$��!th����<�i���=�m����%V��po���wL�jm��'�4�!�}��ݞ5�����aNĈ�.�1x���q�L�s�+�䟂,	e�*3�U@S��Eh�Z >�x_�!�#�$VL§��ŉ�/J�܈�%�| ��O�6vڎ�ب^��NfZ�`쿝DΙ���O �6���GL��r���a#qg];����.X��bY�ZoPZ�A�_�k}��Cm�I�?�x_l��~��0��4ǳ��w��:<�[�a�Wvk���{*m$�ysB�?+��l!�8y�m�󫑼�Nb@;1R���u���{�Lvq�K)3΍�q���0D��~T~#�G,u����?�s!�є�|B�u��Y�B%^�%9֨�q{}��ch�©O;�����o���+�f���Z�=�ƅE��ls�@����	l���,A�sF	��w ���S�0�zB���)�����3��Rc|�a�%j������"ݞ�o=(vSOH��T����+ȫ��N�vv.�W�Ԛ�M.K����nhi�`c"�>��H�d_�������#M3Q��.�S&��8{��cxM�d��L�#�֏����8�H�hyo��,{�M��:��;��}�}kp{G��98bu�\~ �Bs��&>�vr)p��%s�1cQ�AV�1��Wa�/1	�J���a�m?��� ���]=�gf[s¾4�n;E��E�$�8ۨP/�ͦ3�7�싗�R�����J 5ߋ�v�WAч@Sce�y�u���
����p�+���4D�.D�g��z�M-|da���0.��'f�.Z/�'�Ɏ,�[�)�����FI��v��p5�Q�T�?��f��P���9��C�D�dc%ވ��(����s�M���`=?�H�=�  s�24<�ia�[ �q5ˢkdZ�v�ǎ�Ĥ٭�7_V��+���u�]?,����9�.��.��k5{cQ�X2.!Ǒ�(�\v��z���rÈ��a�_`�CEj�Sd�����B�h������b�Y�ԻÀ�ӳ1��H�v�<6E����<~��I0��4�Ѝ�,�Eq�5���W�Ti`D���j�F��Z��D:�34��,&c>�t4.�����G�8�����it(Vt��D�66�.���-�?y^͡1�<po[;�`E�{.��0;�$�`�Ġ�x�mزQ�TF��SK½�.t��'i9�i�(�C鸯�\g���a��X����@(2pT�(��h灦��2G��F�(��1%�0����3���ؗajIu���J��D
��c��j�y�J�'�z$�y �=�f�����!��[�Iɇ�`ˎ!U�j	��;tl.҅(tW�/ҟ8ߖ��%7.	"�p]}7��%C��K
�b�۾���Hܦ��Ȅi�p��T��
��4v܏=���ev��T<+p�)8p
��.8��Q�L�v'�$B͇��