��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CyӉ�$�Z`YZPE��;�Yh?NF��n�? �Œ�>���;Y��A�p^��*����j�Cl��b�ds��+_3�����Lf1dv�E�:�v�&m�gUP����F��X�!����3Xɛ�
��
˦���*����!���W�e�Y�	V�L��m�kR0?�̲��p���]r��m>�Z���Μ"���n.�\��e#��].��v��'�l������j圎��Y��x[�9��@�)"~�6{��� �j�.����ّ����`���=����M
?���5��x�X5����J�?�}J��\=�^X>��bd�fw`�~���Q��w�	��c�Ԝ��x����v�Ar�`�D�@A�~]������i8c��)���1�����T"����=TT� x�aŘ�[�_�u���魖��YzÅ2��Q���4T$*:���]�/���}���`9Up� |�v���:�Mg���e��
}>nn��^ILP���T��1�T�s�a�}�j.���rR����C�l�h�%ҝ�ta��ٺ������UK��(3�u1a���l���U�*�5B��g}��9���x��:�tt~��U/�d�t�g�p�:!�V�UV�Yq�ւ�ܵM�wt����G � v_�O ��a�fm���k�'G��Y$��7��wv}� ��
���;�K/q�p\�ҍ����o���gX]e.%~�aLK���A���X@�e$j�A�M:D��-��=�&�:����Z�h��Eŗy��`�iN����w[��>,�`k��N���IqM��;[��s�W&L�ޝ~�ܧV��0���x��N�����.��V��0�ij�H~�J�!�=>���a~jV���x�b)w'7ŵ�v�&LVo3�!d!^��W��'t��FR�b�FW})��^��57��1CU=w#�D":;�FOWۺn��OD��dؼ��U�$�*��,��!ڮ�z��cVϘ��`{�����AK�G�����<�,Z{#�a�.=n�V��%��S��Ez�����U��.���H����_�,x(��]�a{�&�I�N�`��4�WU��O2�x�	x\y ?c���ο�:\���݇�E_��6�=�բ��dCW�Bc��*��>��m�m-�c�\�uMNHy[kBr��W���R���	dT��F��]�E�]��54���dY�	"Iޢ�i�۾��Z����]EE�X�����L����pA#Ns*oI��B�S2e����GtWMB��3czc�ITyw����7�a1�H;ޭ3ʯ�|�����K��/)�R��f}Z��&�¾��R���)�}bv�h�<�FD�{�>��j������p/qŚ�7���S��J��Q��{��S�bOX	�%�:4q!���}"HW*�c�$�I�	8�&ɦ;a�ʅ4_	�rw����.CXѸ����}q�olT��
ڏ�
��	��"�=��ZκQ�b��J����y���Q�jC�)���^˭�#nj���|�y�pHj�[wN"�tp'D���K�i��J���)e+Cϫ48tk<�6�/�����p�����[lGCp��KL<�N[���ψ��̏p_Å[p:lŔ�_N� rdg�l��3)���κro�~����,�����F���&Z�:�X;��j��Oi�	/��M�5�t�|P���[5�c��7G[�Ly�)���$��IL���)+��*k�e�>[�W�0��/����tZ�<`���;�y�`��K�]<��J�T�4ސ� x��]WaU�:�N�E7�}��f�����5���1���>���گ{t�L2y׾��贆�F��ke/�?�-��,��)Gŀb�p`��<��UFL��"=bJ��% 	����}���� ��Q{շ��Ǵ&,!����P���`:)�%�؏�s:cБ���۶>\7�ta<�ĵ�!����>�L�ȹ��%�*�{�k�%8D���#���gs�Ƀ��D��yn��а�b�0y&���DN"x�?�7!���{T����p%�N�ڕ?�f�ͥ�ڗ�.^_mٖ��Z6��'@z���"��E0:[ҝ��Vp�/���صO��DKy20#I�uu����TS1�c�X`ư(8��?�X����j����,o�:2������Ļ[+*sX!M�ȳ�Zkq�����9)1ߗ,r�������GJ�S��\���z����j��N��3��s��� �OQw^��$���w�0 �吻R����I�r��ƺ�����-{���U�P� ;'uujW8��$w�q�`v�{R�~����A�^�p�3��J�C1�N;ċ�Ϲ��(߸������-�/��M�؏�G�Vx4��I�O��}�:ff���W�=�����I�
�1���&�)���"}ʽ�w�(�z6��)�$9�o��K�l�)b�tN��r=��,�P�ф��~�8�]�	�`%��g ����R���o�XPL�d]�Xc��?�5.g0�qZ7g��3\;�x�+}�ܳ�dÙ8�"Բ���Ͽ-�k�Z_*��g8
�}�HR(�kpz������,�����84�jB�OW�	T"��*���N��1'�?�Ǥ�������w�V��1����O��Z�VN��rH_�B#B��dj�0`� ���0����O�+>�[�������A�Ip���7��������Qhj�4YE��*ơ<���/X۴��v�M�'|�-`�m1WW�͇7���۔4k%}��j�ͧ �)�
e�;\�İ�����|-��+>w�f��!fʂ�.+8N�9?���b��j5�1��,葎�~��Y��Ɵ巶ɉ�d�(��K EB�ΐ���u�}[)�����#,w����n�G�<R~��!��#� ,{\�8�u�'(K� �Fq��
���a��󓜊o��(�1��{x��t2l$g-���]�<��02��T�����s������Ƽ*���:��p 7���j��X�]e������&�^�F(tJ�m���1[�����]��vD�E�����`;0�����x�W0&�Bʺ��N��_�yB�U�E7�oAX�V�$��:n�
�9H��7u��{1c�F$�s��C�C5�y�o��o�Up8�V�ؒ����QX��v�kk3������o�'�� a�i]�6%â�?� "��p�e)\s9��ִ�s8���1�$�����\��� �v�Dj�c~��aѵ��8�� �1%��v�]9���A4�G�4f	6
'�mAZ8���f���6��&���H���D��Π�r3�u�lEN88Fu֎CĈ�"=�M诲�Kݶ+&M�ږ�؊,��$�|�TDdHT���!"��[�+�M�0J|�X�*�L��r��h�b�_��s���������grʥْ���	g�� #j��#�u��,1�;,G���ڴB3Em�d_��R��^N�(&�3�6�g�1�۽��_dN�D-̖�0�`ܥ��.:�r�\9:S��m� n	�Le��1���Y���S?4�@&�_�I�`X����i����-��DYIW���dͮ�b,M,�1�+���{�b�(~�gHG U�q�r?qΣ�iQ󃲮s
T��kV�A�_% T�u:�W|Z��'��Q�	�]�Vbᢄr/���>�o�/��E+��9�W�*S���+�0�U%4��"��>�Z!�&Z�p��_)n/�5e��D :5DX�QO�Y��1��-���4��p'9�_�j@�Q. �_�'L������fJ�ܘEI�Q�)��й_������(�SF��Pu�����S�zm�X��� W
z	�e���W�u���E�#I6©Sƹz�l�r�����3��BO&�b!���`?y�~��e�v"�ᬯ�"���J��>{��OS���CX�YȊs��GH�����I/��ھ3��$��'g���ڠ����IPt�;r���H���Iz�����ԑ��O@�f�Yߍ�_������P�p�)�Y�s�e� +�L��Y�(�ݑ�$�P���y �Ė�v���Iy�Z��CzQVO1��f�V��+Hv�@/Yb?⍄�Ϻ��)֣/�n����{X���7��z'�G,2yb�z�E����sr��*{�:J�Q����;W݅8�j�z�����x�rg__#*�An�%4m�4�@ڄ� Z�*ٲ7P�����פ�;�YI�����d�?���gC�G�H��/D�Oc�H�{�=B�%3y���D��`^2*��LEM|�g�yA���՘�v�]�m&��G��Y����ozoT����q��,eC
�1�>�_ ��
�p��BK�
�K�DK����3��GΌ�����R��*syr�6(K�@Yb�!w�"�:�R�OY�o���*y�q�R��H��AQ��������� .��@����+4�E�Wz.��v�K?Ҡ�����)sĴTf���>zVX�q*�J�#�VV�W_����D����O����F��k��g�*�r�嶑��h&>��8�u:|�L�R#��1_���2����K�Fȕ����(�#���}ܮ��y@�*uY���lY��t������I4t46}D�?�]X��zo �UQ� -pa3��;��<rb�����)���0�N;��0vЯa��t��\���!?y*�D��L��ģ$��pI�IK��0��0]��7╍rU\ź�O��!�g�Q�W�����Ϋ�aP�aS�-Kv��5
6�H���?���w9P�;�����u�2D<ox�,I��&R���]��IKx��{l����U��t/)�P�zXWF;�+������S��/[�F����"���I��T�8�گ,���d�Eq�C��h�F�l�ʘG֫�0��)%G�c��!K���6�M��o}�]P��S��I���i�4'��9�ki�z.ds��U���r�5�mO�����Md���x�߃�:�����B�ů�Ʀr��o�`�񲽹�����]~���jcZp.�����5�ZE���3��^ ����Y�%�k�/�,zQ���
U'��c���q+`s����C�1�=6����u���Ҹ-X�fFb�1@u�ćE���Rhïk�ެ��6�HL��`��;p��.�;t��_�>�~�1.�4�$D~t����lb�D�jZ�iOM�ה���X�\0ndpo���_��F[2�bb���or��e��E��#n]��(P҆��� �[K�e)�V��(.��b�8|�ӧ�4{�X;x5h�GF*���@Tv���Ծ��2��?��0��B�����4C����GNw(�?�J&�Z�pr�kq�e�:ϊ�*��6�)�N�^1�Lm_x�������*K����d �}v�o���G]�'�p���.�*�����/�l��]����s�_��V,����Y�D��]1�&�nNLA�U�µ5�T�!��Y@Y�@�v�����u�&����,�U¥��5�nI�&�|�C�������fs�į2u/��s�Mަ�#N�MK_��3h���
$&��������Y���4R�c�;�� ��̬ܤ�jt�_RB�QNGD��(���������RE���ո�ە�	�ߓK�Ұ�,V�7�d�SS�3�U�S��M�yk���K�A��8��Y���f�1��~4����҅��8R/��3?�S�iV��/��>1���6���%ˢ	�D��phɫ�֤���)zo7=g(o�À������6^W�7�iDK~�w"�`J?~k{!��F 6DqEn�l�'%5���]B}�����y���K�O�Ց��	Cb����,~�-*�]���
З��}9�FQ N<T�#��bG�E)\��y���b�z�y��!V�|~6����@�82<z$0Y`������ٝ��;V�@�Tۘ���z?҄!0����N��u�ӕ�Q`�\�rC5�H�E�x�nG�7�Q���FҔtE6�;��	Z��������';b�������ǈ\�YALc���Dnw���w��9v��o;6��{��8����q��^�׉���9�<��l���k�В�={MIdW�����}�isA���t��|]r�޳,�	VFJ��b
���ɿ�>n��|���nb���F��9�gLE�ń��ʬ��}�L�<��q��!��]���Ѧ���ڼ*!D4�Bp��;���l(��6�eAd���ϔ�f7a�p���(��3\̅���OO�-��UlW]��`U?w�q�XQO���ώ��[�*6ʏ�uX�}����M���
��1x��OI"6�F�V���o����+lhv����ģ	~��G��j'`f�O��JW���i mG�F7�ut��|=;O9��M]�:�Ҥ��5@DO�&��B=J��"�_z	Ʒ��i����q�����(%9Ϭu��={��x �q����/���I�����<��
�Ú���#��}̨����	I����+ ک3�b��h���#�6ϒ,� rES���w���t��lJ섫�є��s3��Y���H�U$��q��C"����->�k����{*�rȕ����-�ΆnT����|BPd�Oz��m�hq`+U ��B���a��Rp�R
��j����5�s�&?A��:=֪9/��B��P;C�X�-l��{z] �m�y*2Wd���������1L�MrQ�d�@�I�0�?�갤ލ>���E</R�?��b�F6�z\��|��o��ֲ`7X����T��v(�.X-���J"f@��4̾ �A��IA[��u��{���U2�0��#;���q75�, �](g�S�+�1a߁C5b�Q��J+�����SfZ�W�tHK�V����t�y,�-��m��:L�ݥ4퍏����RgX�Y��Xʤ�ixq���u���q�D�4��6�ڡ�]��8qO����8 (���'�!�"�=N��~w���k�_}�ц�j	��'(EV�D�G��h�-����f�9Q�ؾ˾�2���%?{�6�	�ĲN���~�7��>B�-yC�tW�_��E�ya}�n�sp���7Bc��x�A}��f�]���9c�	pvu��va��A�:!�& �O��\��������ب�m��61� ܋f�4���Tz����
�������<]]H�ahH{�0��_��X͊���^��7l;P����'��6�m��� q�l���/WM�!�%��A�-�z����s�V}n�ޫX3!�����>ّ��lG�a�y?�)�p=�F��ǎ�7�(�T'���=�C�z��U%�d��U,�R��F�)��m�#�}ǔt��{���Տ*"ͅ[��*O��3Z�g�}�r����x�3p����'q��'3���Y��́mU).�k��i�3%����]�Sm.�T��jQ׌���u� �Q��~����?g��
>�h�¦���M�
�J��1�|q�3{��]3�y�`:���HK�j�U�&�XT꫺�wa끪G�Ť0�o^�"H%���cP�b�u��?)ba�;�B����!�ML����Hv.�L/k�GEQd��Vqۥ�~Z8T��C�.>�MO��2���rɰb ��g�B:G�� #��������_�Ǵۙ� ��0,f]s��_:�&��!�����ͱ��M2���=��r��2s�0�c��	=Ǳ��S�}ۚ�w��������4����Pװ%^󖰑*�f`,{�G�+��C$�\%���n��H�t�p�!(�O>����(��"s��h�m�Zst��t�;�㎱y25���r�"q�i�o���B�,�3-u��引��:=y�/�z�\�٤v�?TqX��/��z|��.�}�#�77��l����
!���"��Ѿ΍��$�>�D���z���1���1��$plw�7&�:�+��%�2g�:��/��nn5�������c�M	3�1�7����=�H'��V���>��xE��"W��'RDܐwPX�-��"�~�Ք���D�xu�Y������K�!�QG,z���Hz���ae�� �\�ٔ!ˮ��m�Y~�1p�a`���6Q�`4P�R�mtlO�jw�Si��KWi-�O�$4>v�6S�ï
�e�����$����{�C.R���/qs\v�jrD�[��T�b�z�y�f����c�<'�y�p�A�u��L�(f�(\���@+��e孌��!�C���H�":�ۼ�j�r����t��P���P�485ܒ�ד���Bɘ��%f/}�����i��#Y�R�h�i���P;߯����j�8X���-��= H�u[<���	�����ޞ�Z<�~p|�x�k���� &l�R�v�U�:y�dJ��~���PK���6n���#~.���`��J��j}Zʜ�!�T �J�9�cܗy-u�酵�Ja'�3/�ѐF.�X9����1���btj>�����<�@���ZWYB�s���!���Y�{����,\��n�R	R�����*8��Vc��J0I�����>�'�k1#9F��v��[;�Q���g(zxHT�E4���U,�Y7�0�ΥV��{VC����Z>8�Ͻ�fyĤ��N�SQ,�	�"�T�X�����򓮕z�h��y,+bN�2^ncj��,X�t��#�GG�##����hƞ���nod�*��5�3�RͰ� &�ʸ�Ye�育�$�����0��ɫT	�(����\TR�	� �����"i( V���+�6�H��ɭ5o:o< ǅy����ͦ)��]ʍ��+=휏XU�2�۪r�͂����;Ct<���B�G��̀�{]��:�2�:����U�"���W�2�BM�c��yY�c���_��?y�R��x��6��0�z�P�zO8��c�oTm�:�	