��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O����Q��VT���NQ�h>�d%�V9Vn�|�r0N"I��P�p���'�O��q@4��F��*��<"� �`g4�s���F�/+n��_�E�@���6�� ?�hf�v��}x�i��1o�bl��H����8���-��N�+;�l��H�ˁ7��kk51�w�W���������@���P���r��\Ġ(�P���c��;���*�$��)��?�m���h���.#�N��=�8��#��swG��s�c��d��g)����y�xw�X�.�NN5��V��sп�a��D̫����8�T�q�b��Dr��@�u^�E1e�3F��喺�1���y��H��k���cs��A�K�%Dm]��[$"J��s�td�~ջ�H'������%h-��\L�T�w����2�&�����Q\��M/����%u#M����،��;������s�\�>����D��9��	����謘Y�C��ñn��R%��xO}�����3r��$�$ _<��[�~V�P��O(^�R��9ȣ��Ռ������n��v��t��k�<���x�c�r�<C���A������u�˖����o��r�륩���%��XI�3�"����B���a�#��'�W`	q�SU
X�OY����3=S�|%�,�M?���Z}��n�I�7�B:)�����AT�_������ WL)��ًʚw���
yL���(�[,�!G:T�,�J,�r��]��XY5oS�):� ���1�Tz���br|$H�f�"��F�ZD���Xu'y�󻬦�@�γZ�"$�e�(W3�GdЉ�Թ�Wm�j�e7D�SWDE��_�"�~�	�w��`?��'���2S���H�P�/qt$!�F�(O���y�VM����#z��RU�8B�pb�O@�R
p�H=��������}Z���M���`Kō�m�mQp�KL��'�E��X����-��F�_�_��^���C���������fi��C��ke�)�������G����$\���^�w%f&8��ZL����Z�� �����D��Q9�}
-g�ʯ�������E����7���;%�׾'�\�������^0)�1w�z�ٚ�T����Ȟ�O�f�	��9G#�l"F$ر�]՗����@wi�kf��~)	�=O�ůؔl�lvB4�0{�VemH"�n�r��x$��lj�$���]��a��2�1�gā�ֻQ���;w��W I��lj�1}���pe\�֛�f�YM%#7"�G��UxW�|n�@Y9��ZD�h����S�2Q�(	ܱ�=�>;"G-�2k�`%�8l�Z� �L�n1��5��U�B�d�߿�3pb���O��y�`�J���/wz
i�N� �)�>�PE6:��='@�<���i�2B�<���'V�_V���CC�l�B��sa�yߗ����>��@�oT��
�"֊E���W�9eoM�ݹ��vn1��Ў@��eU�k�a��ŕ�������/��q��c��ހ��s;!�-'�nT]��G�8�LԌ��yޭ=brV@��#�^Y�kq��
�A�pP}�e{W��(�5w�_�>|_TaHZ���~�T���V��ɥ*zh�M��+~�n�� ����{8�@DU�u�V�|0�e�A �\]��T{S�=�6i�T���r���	&�iu=�B��lD��7������2Ҡl��Ԥ�MNq���8���OAA�۱}� ���M\T1���]z�*�����!f��%�6-� ��Wzo�Ki��[/�g��[쀆�7Ơ�l��$���:���o�:��U��Cce��T���d�H�,��x�TFf��I�O��de8�{@4���Y�	��E�]G����9�����)���"�F��E��iqf��2�P��^g��b�8!7P�;z(�Yֲz���7��pI)K�I+�W�RF�(\�R7�$�G\@T^;���~u/.���y�6^7l�s�I%5ŏ��5��i�͢S|f�JMcm2Od����E�S�<��~�@��M��|�'�a� V�����'p-!��+q����^0g�B��(��}N��Ibd�8^(���&�͘�����F�ӂ����)ѷ�- 7:/�Y?ݙ:��BXwԭ��w�Y��M<xVo5�"���<g�JS����ɐ���b!��|؆�)KJ%	$�u��	PQz�U$�<��F��cWf���
��)�&��N2(U-��U�x���g_�$�>����A��1�R}��[Ϯ8a�	���9��/���|x=`x�+�l�+�^ɃOlKX��$]Yk� �[��]�g6�V��  �o�����N��b�p,�������9(����i��V*W�/��/ǼI�9}HY�e�/��Pl=�r�$��yyD/�QG�E�*�������х���C*.�t��A-�� �U�V��-��&�Oi�tJĒ(����dK�����=	�)�Ļ31AEr�{����ܨ/:P+�h���O6�8L�:[X��?� $Q�ѸW���T{_*���"z�{��M��}��eˋBbj���E>���Q&[��"��8���m�8]����͚����k��Z<�;���279��h �J/�#pO��z4Ci~Y!ǋ�Y��C�X�O��ۃ�x��j\����Qz�0�͠V��7���+9����KC��[��h��nab��J����p~�z6v���3���Cq�d���	�[ՏVnF�Ҙx��b���(��:.�2���$
��Qc=�9�~+݁§�7��;�z��wJ`i�4?��Q�9�]C�}D>�h��=�1gU>����{.����j���"Q6E��J������X��N%�Bg��%'R�v�2��=o��?�G$Ʀ��ʉ'џ����^�p��vLW3b&�ֈGH����U��z���wR3%�(� )y�9�70��5�y���ՔX"nE�,
�h�Y���C�#ؙ<�˝���L �u� )���h��Z�;S��,Q�X#	��BA[~�$�|\y�0�V��7o��MU�	.�B;����h_©6%�gpPuO�d��14j%]����W��
L����veuX|}ËQ�r!,ݻ��%4Ə;����c�+u��� mJ��B�h�؇.�{=@���ǜ����lj��{��ц�/�	�n@`�+�~7�X��8��T�2�L��bW���^ m:�4�;.�/�� �c_<�4��z������E��P��nL��Q��� FD�?zq+��meFlHx:�\R5G˻lt��_�3�=0^&v�������O���]?�c�4��[�R&�xy"c�3�$y�"�dI����^\XÉ0xJt�l�).s��ell��
��,�ڀ_*��@�.��a�a^:.���
�"r
�w�9�񯦡�#A��iݟ�V�F_9n9��N��3r!m+�2�����t[��>��3����>��u��Q��2�{2�S�Ѧ��ɒ�Bw���8Y�&�G�eI��җ,sZ�L�>�� z��Q���f��^���u�7�9���:�}^:
-�8�"�e��;:[gM���x�����ȯGr�~A���d��\���p3|'SF9Ӆ7�щ�υ�@g!Q�	��`��E�2�v��0[���^D!ͅ�m]TW�#*����$��/�ĝF�����f챶�Ҽ%;��A��9g���? ����땎[������y_j��`����ү2��Q�ЭGB(>��QV���'-�^���)���\�m-W>�;�t�v>Ѵ0g`��׏��Y��Yëa_,)O?�?�F�z�QFu��ȴKG����XE�����Gk�:�*��{H�7Yh<��pLU���H&�u(�=�2�S�aw�P��!d�	��)��k%�?�aj浀��DR�L�
2+�Sp�z7�u{��)^�����D'p-���.$(A���8˝�-/�b_�,��ʢ\\��:9�zP�����ﷂ�V��8�|���4�f��t��5�_`� �?�w����+��-���-�����R�t��JS���	��Q얼fr�&|�jlT��rx~^��I�W��Zpkl9��"�Gw�=ߓ�r�;��V4S�'����O�E��,V=N�2,(��X��ĵ��W�k�g�J*��M�jj�	����`��f��u5!mHۛ5z��F����Y�N�pnH�|i~∆<�~�ڠ>�)�Ŵ�25Hh�A���� �^���9��[Şŗ} T�{��U;0b����t4���i�Yp-�䍱&"9�1$��Y��My|h�;���~��$]蘂��V��lV�i�}X������4�A�@y.��!���AeV)�gs��	������5���`7vAH�q֔�?\�Ɇ-����4�x��UQ�\��E��� �>�5�<�z�)���3$�Q\��V�*���ӻ9��}�	 ���VN�yL��,���9ל�=��\{y�S>��F�= �8��?���[�cWK���j	�C�(��fV�}�+��)��(Om�V`J.��p#�k8��:� o<,���"K�<e���5>�S׵��\~�Bz0r�It0[!L����~�%��w�����d�9�P�)/ X��ǩ�uM��2:ҡ�ߟX��q��ev���(�B6u���Q��hYv��9P��[�U�����ů�ၰR[���s�8힡����!	���f�Et��Bz�o�:ϰ�#$YGv��ȇ�4�@�4��%vap�[PU�0�q���^"��#\�8u��}�h2_\�0؎��Q{$�}ǟ�c`ѿ�C3�'m�������������z�~�+�r���F��YcV��mɤw��q�=/[��R�S�f+\�]��ްP�=i��U��%|�ݿ���$��4� ��������
�-y���s��'�
�}�K������G|�BXV��N	�ӦC/;�)�V� i�$�z?~�f� @��c�O{1���lDiT�0�]t��2�*�
|n�i���>��B]�P��C�zoR��"�N�[;�dd�B#z�@R�z��>�6������B�{l��CRy{w�XIW���`3K���;��TASo�hM���E��e
��n���,��z��1P.��M�SC�8l�ܯ5ΓE�u3ғ������<����5��I[_���3zllM6|z\)�i��&����ΘU�m0��H��6�f?�o����r,@�"┫{��"+1�:o�6�T"maD���ݡ|u����P+L��N���ȁ�������yyR���(S�爏;��jxs�`�3G��)�}��LP�!��Q�������6a~D�9	��=lUES�eUH�FM4i����,���]�����9��ۜ����Ql+}�C����lk��d��@��f����5t��/�[����r]D*˦�*ɹ�{E�<��3�z7�/G��%�y����ܮ&Մ0��\E��G��IH���P�RK~| �����>Oѩ`aa�sg�>�hǈkYn3Q޶�`�"ȐW�U;���H���?��<��m�n#���aX�.���:HW�P[��	Z*,�v�5������=����P��h�I���x�L�AdE����=�o�l[��1)7� �+e��o��0;o6���(�;=�׸��ઐ�௬����+>� ����7���傟�ˡY|1�/��V9�$��R�<?u�$��#�]S��~<ƴ�s_336`��k������ج]�~�>RR*R=��1����ٻ%�ňm'[�k�3�!,������äye�/y8�տ+v��D.��y`�wl�m��9�ˣɌ�M���w�����ːq����`U֦��%^:�`�B2w��W�v���w7X�`��)��%U��
eZ��g�$��[�9I�|��~���;'L���ê�u�����f��RQ��oˮ����iUS�ޕ�G�<g,�'��β+x�^�L?C��̿nN�Y\�-��0%҂�H�����?���@�yK�۱+��u(�G&�
���o�F/%!6�WN���~>��Y�CV�o5g�}�<qA��`T��WI���,Ԏ校q�Y��6����q�%
;d]ߚ����Z%$�L���04`!��[8u7$a�i�,~m�����0s�f*�ݹ��qy�d�@���D��0ō*'�&�^�3~A ��U�4�s691��F�;̬C�8�v ��G̋�w��VK+���d�;���?R�rV7v�	����Pא��tw�ogݍ��L�@B׆{Z,m4G�a��o����9=���%�!:l-�r��;D^v�m�$���ޕ1I�E>�?@�	�Ӿ�f��r��Z�Ø��tŠe��Am!fZL]x4��0�j	^���+��-�t�D�&�蹲�S&�6��E�!r*�u���/��β��%�Hv�u�E0ظ4�lVt�"�Ta��/� ��+���w�%AW
�Z�#l���S��W���%���裍6q�@� �>rB1��s�d"�B�]���*�����wwl?��R�B�q}��;-�ڕT�����~��:��V�S��=�T�W5G�M�ފ�[_��+��۬@�{+6�� `�7����&~�O~[,1c�dm���#��Ok�/Or�ú��20�zU�ݛ����.L�wJ��N]�J��G�.���V���粒�������?��d�})R�n`Y�TA��T�! ������="�t�h�2��q�DX��~��cP��xm+_pU�扼�7�L� �M٭:^�	�V]1�$R�����/��Z{ؗ9bD���5��������3�L��e�X��C�ЮPK�
�(K3�j�
wӟ����;K�Rn��]�m�*[����3�Ő�7��T�c�g��u�h��%^c�� ϽV����QA���]�lR��\1IR�Gڥ���典	��]b��x.���D6���Y-2rĢ<�I(Qh0�[�_��{�t�j��425��-sڜ�	���q�[n����N���s.�`
�^�Umq��Ϟǝ�p<��a $Z�߼Sv]�&Ԥ5��Dl|[p.���:���7u�� �a��RH�zk-]��r�����m,1��j���<�Mf�UNM�G9��:�1��8R�E�8��5q_�ׁ���~JE�~T8$xZ)w�TQ�X��
��' ��oWp��<�p�Q����~]��a$h~��z�y_eɜtq�tzu��#��9��L΅�Qf�w�[3V�v4	%`���J]E���Jf����Pt��2�EG��_z&ͅ;x�ɿ,uG|Q�A�7�'ߕ'�n}�>�7X���g���B(���'�ܾx��� �r!�`�z�C�9�"�Xca!C��_L�\�Yj{|FOE(<��S",���>�^=��T~���/�Ӕa���Ø<|Z1�OÙ�a{<qiE"P̧��� pƺ6`C�wo�J �f�o/з��[��(	[�c3GYQ���$��4&�ed�Z@i&�A�H�<eӗ��ίsrS�ץ�Z�wL����G�b����-�'���l���-��Җ;;�'�����!��D�	�U&�������F��5p K��*�`�ak�0`baw�G�ZFR�����	rߟp�������3�ND���v��]�"����&6�۔��ܨ�O���]�_]��^���i��v,2�)��m|U�#9�#&>%Z�~�i~1A&5Fuk3��c1ҍ�V����z����?~�I����ڈ����C��])���X�x���v����Lkn�逢GD�E��-����c���y:��R�F_��X�Y!#�w.?6M�\�P �wR����9L:k���+�<�V�^ ��Ct����p���rF�]}�A�n��]�@h��?g�8r��(7���I�f�
^rָ���.��3�t(h��8ia�T���c?N���v�
��D�h��*�I[�#��y�+3�u5�]b����7�JP��ЇΦk����.�o,/P�ؽ��Q_� ���9�͕l�B�z��_�F�yb;8s�yhٛ/a@�y�o%o aJ�~
��b�� �Yj��VZ�e���I� fEw��jT��Q��yG�t�MHs�`��.�
1��1��ڊ�n�B���QK�>��Bau?�34�V�x�dKuFd��4��}�������p�oѻЇ��!���C����n��]D��cZ��z<�$W<*���� "�磬y&䑯�]3#���]Rp���ED��(��z�z��$�д;A|�h;+�z_��}91(A
�LK'0\5��� Y��UMq Hm"��gE���;5H ��rG��X���O.��OGQ��5�\E�3����(���c��e��{��#;�y�6���S�@CYC����D\Э�^jk)�Aq�qzy�
_kv:lmln�nf��o�$3X���$�;�s�Ô�K�Ր��!�6N��v�G��cX;Vh�A�=�i���R��g�y�Z����0$������͹��Y��P��H�u[e��T�l0��%���x?�'x�H��]`�=aA�M��P�Ӧ7錒]�9��Sa1�뱿�m3�4އ=��iS��1D�:�(��f����K���.͟`uC54:r��j��9�9&�-�Ε���i�2�A\Iq(�'o�@���H��lg� X}Q�����D)�u�8<�fB��u|`��dE�}�8[�"�RKH��������g�b,٦���ʩ4����p�
n�ea�m�/�TuP��å�_Z�_�g�#�7K(rP�eg<ru�k�