��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����lĝRFĹf����;���cc��`*���k����������$���ǗV��}�1D�.ꎔ��z����
���i�(�\�a=V�Ѯ�k_�|%#Ǜ������m[��[W`͟��Z)֖�%��k�B^��2����hOo�{�Z`XIs��d�1k��PC��ǽ�����	�EU���K��ō<c�D��[�<�Pk[��ף�^�9 ����D����c;Z`2԰�TDg�&��;E�g���:z\����J��9�)S���>'(^���G`�Ζpɍ��d1q�
*����_8��?�U�� �DBRҦ4}3�:�
7ņ�&�"�:�x�p���Ҥ�l��y�rG�Py����8�Fn"�BBK�$H�����N]�9~��ѰkϨz��]C/\K����!��ie��@�Z�lOZd^n�^M?��s�O�Ƒ�j3����4�	�Y��c{_g1,�;��L��ߝ�k���]b��>�����="�f�A�w(�	��Y�p*�#~��
v��9}7_0��L(mZ-�SW�Ȗt�gj5W�lv�[�7���w�� ��'焌����:��<F��ؐ��I��!>-=X����L%�dħ�!�+:�k��v;�ܧ�xG�7
=]fxzC�Zk8�?�.����k�n�{4e�T7��'�����d�~������^H=�H�;k����
{�KU�vo%&�L�&̎���V��>C���a4����5��x���V���?��.�ج�~ͷ�_�-��;�VH���=`+F�����T �|�Z?ଧ�0��2��f��7%;
J1?ҍ/i��s��=�����!wjk�j�@���z�[�8�\�T�p����Y�O�Ϸ{���U�ޘ��dx�g�^a��l����R<e�]_h?�x8ҷ��ꀴ�-��n`�`�s���j��H��&.�/�k�+�QD+��쁻�F<��x�4�5���^Db74>_�I-��� ������&��x:�@�"ZA׀�Y&��b�������a�5Q��0��G����XPH��Z|C9�2&X���=��qsðQw���c��1.���n�{x�)[��*yR���wJ��_�$;Ce7��`����v�)����ޓ(�㗰K��Dު���Y[�x���y���T�n~�hRT%���1=?\=�r|��-�y���-�
�$�p�qB� ���+uw%�<_��~��km�Q4��*��ہ�����!!g���*+Wx�O�zjК��c�UX�lY+Y�x�%ǽ�p�� C�'I��3�3	��B�X-�y���!�NA�Y����S���m䟩�QO�/ޞjZ��\K,է��f�q4Wg�P���g�T����Ǣ����g/���s�[��j��u�g��8�O�v���O�����FvV��ȦӪ�G%������r��k��
ꜵ>͠b�ak�H��u�����^`C[o��lMZ�sCG��7(a�U�	k�G>�] c𕊪��u�7a�����P�-_`_t^lCvrF���٤D�5���ۨ����	TB�כ�J^��X}���q<�f��R$�ꤛ��A0�.l/7�S�G��C����M2Y=�o�(�A�0D􏃲�܃n��H�[J�w��&��>0���nوIL�����Mp`��7�i��:�-�
ס�_�� {�yj�ȉ	��퀛 ��/���H=�<�p�!�"�eM�ҕHaT������rr�a���m|��%M\�l�P��h3?G��2y+D��AH(덭G�n�p��(�l�5V˗��/H��!�^3�9�^��mR~9"�ѭf� 1��%ZVM��a,6Ŵ%OI���@��?vH�Wq��; .�Cx��VT�rZ+r�~�`���q��6=���s�@�6�Ɂ�Fu�u���!8��DlJ
��$�@ʾTH[do&f�V�#j$R�J�M0�6�r������CA(���l�iP�		��ٹ5ߥ�jɫ�0��p��(��b�p����/F��=J~�ݡ�&�Lv�,���}k��\~��.n�*�)�ǞP��u���q_���臜N����c�ֲj}�+W����e1`�<��g{A��ܫ<Z�Uau`=_�$Fm�����	`V�����y�v�꜎����ݩh�`uPy���@�'��+����H��İ�o|���O�{�
�� ks�ǅ�<U�O4B�B�z\���Sz��֍���q�	����W��{��R_Ts�s�::�R-7U��Qd��N&bؑ>��5l3�G����������J���*����0#��?Q�̪�y� ��Z`�lB_�J?o1�Fw'?�8p�dǰ��_ϰ>���U�*4z�[x�m�;��DU�{��⻭��6qlTEV~�?Vu��Lt�&�E���O~b���*g+n� u1��<<�_tAV�"�g+
�[���b\�q�"���}*J[����>2���R�M��5����ŨR�n� �_��^�V���r���T���	0r�5�=B�� V0�=	���A�pϿz��_��?5d K�H�J�%Osύyѡ�L�Bj/��������w�w()�::��J�JF�%2�8�|���/�����G���@�2/�c;�f��6DѰw�Ml�> =t�\���XM?9�^�0�ZkY5C����M`�1�(��%�h7��8F��YU~���!���T&D��wi5��lQQMcs��!<[��u'�e�Y�R�/$����ZN{��Ӌid~������ǆv?�3Z`���A����=����3��TcF�y��� ��|Z������{��n.\���r�)9�8�*zQ�Z��!���D��?�e�9\��3Ί{L�^c:}��8]S�K���Wg�t�_�R�Aex���F8)��A(�M/��\�x�U�Í3)[_�p�[���HށC��v�-���­6����+�>��ڛ�zj��=p�1�Aa;P��.����#�T<\4�3TMm<G| Y}o� K�=�!/��'~\�f�`�0O����@��g]��[}��DGQlk���%��> C�:n�{�D���)�C���	(N�C��@��ē~D��X: 1�)ٳ@C�Yu9�����1���?�)�D���u�x��<���>���(��v.��ƿ�K�R~Ȃ�x�dXg��Q@�"�Q�p��y��W��b|��C�AK�}@�ό3�7��o�"���b3y�j_A�O���2 ,s��߮�>���=ڤ��\>��ֱ�����*�D@U�H	���#7ݱA�T���ipw�أ|�YB2�5�m���>�ͅd3�ݟ=����?VA:GԌt7��1裷�i1�����u��sb�Kk�Q�|�jh���<�]9`�l�O�ԮX�n{L��;)>���g�Ɗ�I:�}@?w�`�j)��ƫ������"i�	����bD�"� '�R[ͤH�bڹ������Rth�B�%��:c�X.�O�G]�eʗWՈD�0eg���J�u�@���Ҩ�~����&Q�I�Z��Dj�+��>ZL^��Z���nw4+d\�Ѡ��aS*Q� �i�f�?��&�{]A%zy*����s����\�[Q ��[�2so�p��f
)�����=�u��5�n��G��9`�n?��V���c�$V�4s?j�2Śz9�m#�k��~ZDl4����<�*ؽ��~T%�E�~k ���:�����{<(��$�'��#� ]����OD�;���i�$��]�r�W���ix����>�@bQ�^�?�h��S0C�!}l�)Zmk`2K�}����W�Ge��T����IKݲ��fGk�o���@6�:+�� ��9�B@��`O�_;%n>a�CL�u^����Yf*x��ӡ�v�D˖}F�p^A�*��=Eݍ� ��ҡ4��]��V��:�nG.f4�_��9Y]��Az�/��ty�����Sɪ�̽�:�%�'�6v�R��&�n2�95��Q�!dv����F��h��)��x�`�#`�EI��<��es��`�B�N��Ʀ��C�*��PJ�S�C���)��y`�,�t��ǆ�
���Z��ؘ���4|Y3�����&��W�!�n#*��i���n�t�w(���Wߏ�G��Y�W��\�],6-A9���w7?��� y\<3>����@���4�c�����8/_���1�=�\5L�	�z�*���">ҙ��]Qq+B3x��A��۵qщ�ˆ>�$mD����x�N�\���	���[b0�(����Lz�%�'J�abJ��R�0Ml8$����o���v5&��e<���Yj����'�1�N�7Y�����ؘ��#���Lp�����g�e6T p&_��8�^��=rg�%��2*mr��]f��Ȱ(ވ�wpVf�U��=���=��ƭ���0D`j"����� y��NɎJ��:�ş�r��9U����z�e&ߑ�K}){Uʁq��%j#�E����Q�@���d|+�a�M�~SQ�f��{h}�/.�s.0�ޗ�`ɜm�O�إ��H�r?�ʙhNZ(QC<�b4�<�_{�,\���>����X�����_e6'�t��}	
�)k}@���(2�,l_؁�t��9�$?�ݮ���B��T�A��E:_3��+��H�>l�vշjA�D���r�K���I�����!��<��x�B��[so`id�#�0��K��83U���W^	�3��Q�~�sLP�TT���G��^����A�Qz��6n!Cz&̔^It�x8�q�u�G)�T��7�{O4ݔ�kt�{���Y	⠦������g���H��&�ц Thxc�����t0�ς�~,Mɲ����U���|I��O��&&L��b���ou�"�)k��&����1��b�ڡ��T��&�	��Ʊ@��`��!��%�t[�,��.x�X������|�1v��v�6/�2c�~0=.�r*�鲍�"b���c?��C�_���0;x�Zu�
�ۇ�<#��6P �W�jڡ���$�Z��S��`��<����q��&)�ݒT)^<��� ��λ^����P���Rf��q�+g7v�l6���ECp�+C�A\����/�6�ӷ��;�]�P��pϑŊ���e�✀�P��H]�gX�X�uy�\"#�n���Κq�<
�5��T=�CƐ&$+�tX�b����L�D�l���m�
C���ĶrE_ᲶO.�����ڗdM6`#E��+�F��Uݏ�4���;sN~z�&x��oVplD�|:S8_פ��w�ytU�ԕ,pe�������]A��rL�m�A$!e�t��|�#[p�&zu�����Nϱ�ܕ�f��w�&�U~�LkBJQ���=�'�����N��h�A���v�d1�_�	
C��	�Mw����~���Oz*!� q(����ʤ��e1�Vm�D�q/�ߞ������>�m_&ʄ*#����K?��ٲr�TQ9���7�>�~`W��M��Hy&�>`�I=�#�B�/'�&? �/�0i�ą3��� .����? �aײ�D�d$|"'p#Y����5D1;7��ɸ�ږ���C�����%Ku�`9��3�"Vo���b��P[�{��\d�W2L�r����8�x!�����M8�
��)�3פW��xow;��i0MM��8�}f����h��6f��'ʢt���k��M����~��k����M0N�X�v>���~F�jw��� B4Yn�u��B[���ь�@Vܲ���� �=6� ��p/Οiv�1�:��r��h�P={�)���<H�N�FG��&��N���+`!��+�͖wv�5�3#p}��=�L��3<C��i���J��K�b̦�j��FC�v��9��ڛ��%��и9z�hD�E�zF��9��5��ϟi7��1�h4^���dqz`�Po�1�iF�k{�)8 ~���U�T��z�D�{���?f�PeD�-�?��3͑�Ѵ�r)c��o�OfM�g(+�d\r?U.�톉8 �P]r6���"��2&�.��צ�z��{�	D�Ӣ�>T;3���h½l�Lɧ�(``���	���G��|���Xg�P-t�+��<��I�Y%�B� m�b8�9�݌~Zkr�ݨ�+_��;]�L��te�~��~�]�����)�{TR���!�Ӏ�֫3��_Y��*w�a�t1E����@|��Ѷ欠IA����^+���Ո����^����ZY;S��*��RCj���h�&��Q;qz�1%�#�81<��5=���\1�>�}^��>Ũ�sy,j4P��U��D6&aq��7��6#��K��2���X�D��+�+�3S*�0�֌����������{��u|@��1&]Q5`J������$�/��\��4U'���GO{i���Q?���aW�F��yI�� �9H�>+}	�Þz����5\��,X��|��B��h&d���<d8������q0�ۑ-[f��!��_#�vk��U�8�����°���~+K[�ِ^�B
���%�����<@Rv'i_�3ږ���,\�z=|�妋�_O�L㵴�Е �Β�h�=\��˰c	�߲y���&���6r�ls�+-��FV���Lw���<��h
�]��& �����-��Pۆ� �������E�4PG�y4_�V,_֥�/ܧ�i6�t�(s�K6���XY��Px������(͢���ѐ���
]x���J�$͟�yǴ��~r����/��]H����ل�Β�MH@Y���w���%Tל�u�{����x�в"����ͭ��H�����13���\�\��MG$��p�\�;{���Y�y���
�I?Ǧ���F��b��	75�'��ig~NnVrOv����L�f�$s��qߙe�	+��>�V��Db/�"n+N�f�Idw|^�$�/r��"�mk>2��B�P��`=�d,8$�@�mP��p��?"l}�BT�Ӹ]�.�W�ӏ���9aU^<�F= ���2{�i��@���a���O#�/e(�{�!x9rZ^&����h�2�/��~C��A�_Z�$�[�v�$�~�s����l��j>Ƕ���O1��l��Q �t4�D�q1�D�wLE^�`ȝ�n�y�@y�0K͞u&t�w	N�^���Y�Maj�P�~Z����1�h�W�f[Ie�	@�M`�����K�5�2�g�)�>�����Zw���E�8�h���{�i����[��e��������\���xu�EJ6���5x�@�T���x����K|r+=�kId�9*��&8^!��|	a$�ͫ&C���<Wr�2|���M.V5Ln�[�T3�]e��Y G��6_Үn����'Ưj���X-Y�ye̶�y�R%�q �Bǹ�:4�$%Y&F`�j�G�eur�'W�\_%Ftp��8OX�le��I@��\��eV����[|֊��L��aO��Ғ�#�B�PL�jҎb��:�L����ܵ��W�ærwS��y�g%�R����@��W�8��Wb���CA�>�`���(��2��Pܘ~`Q��&�-��=�J&��j=z�$��_�����si}�s��.�gO_:�0M�;�F*WoX��s�G�ë���`q���ѐ��{���v����:f�?���y�ܚll��g��c?8�n���7;A6�)��cT���jL�xh��ls�ie�LN����S;���]/�?�C?G�mh��<{z�X.�?L��x�E�5�ְ�ދ��r [��E�@���~ʺ��9�0�S�*�<)>��0
`�p�"BЋ�P92�b�d5N�:E���S��,��<��&:�1\�ĭ�6rx!T�y)�����c�ǤD6I_��2D;�
�'A��n�w��98a����_��e������&_e�6��o���@�[����/���Tqۧ��L�l��@zPe@*��+}�X���Z�89�����֟�2��l��nl�df����R�lu.�6h&������?�����&/ɜ��)^;�.;��C�Ak��M@�O�st�\U�$��کz�冗���n	��4��ς�����PP��G^/�N�l/��'4�/�T����sF���~�%Ym�8w��jT<�3xL}q�5���\���6-��ԋ)�h���]��a�59�mu�Aq޳�3�Ӳ���m�o�>�BeGxl���|�����N����uG)����BF�g:{/�
5-�F�?�5����44MdL&�T��O���u�����}�Fn*^���e���k�J���9����
GpЄ9���vR��:���<�k�ΚF�^�,�n�P�E�u��(�5��0�c��$�{V�B����p�!6�k~�^��PR��*��Aɾ\Y]nvE��q����E�����v���&4R���.,��H7� ����NM�"�9^LJТm��J�o���Og��8|�crt�2���T.��e���x����ug�p<3�e���KR#pX:�*��8	�[��m�N�<�_􊃌��GW���ȫx��c�|X�ސ*��|�am����u�"[7.�3N8>?�7$��y�1��*pG�Ԛ�_���$ �x���O�БuK�Mu�� RV[!��;�V����W��
ׁ�6�o��.2D隚�=6�
���zdܲ�s�Z���� "c
\.����*�셣�U�P���U���֝�5�}�����ʉf\gu�p���2���x��K����嵑�gr�e��;e��	ӥ?���#�/R��=�ߜ���|h�h�C4�wݔHN�9�z�sX ����Ė觚{�S�A���LNy��s�t�{:Da���<��Rün���58�iͲ���#��4�bx�7�<~Fb �ɬ���g��X(�����f�9�E#+\ś��*0o� G
�����Fؼ}45n~�)�IZ?��|<߄�ϻ]4�B$S�Ku�3�(W>F�!�"YkO�������m�|_�p��jp��d� �h�k' _���>�כX]�8���/������R?�޳����;��|��WL��:���=j)$R�'�!�1<��g	f$�.��0:ր�Gm�M!�2L�BH�,���-,� �y5���Nsp|�0�82(�o��zV���i+T��:3UJ�M�s�`؅JY�sˌ3�8O@U�J��q�3�{��3�ϯe��51��E>'Q{���ZE'�V�;q8��"`����Q�֬i1�Dv�h��ܨ��Zx�,H���f���	�W�NƤ;C����D�	����*��Jy�C-��-�g�9�;[���a�>=�x	9�x�*UB�].GO��. ��(�?���W���W����*���ʱ��sH�h=�悱(g4����B�?��2Iy��{��<�.�(�J0������H=��RE#Q�cO�9�����w�;�^n��f��O�����2����	n���iI��z��i<�~�Սp=@���ޜ`aD������:��e�_,����H��'�/0�{�3�!�xr7����cE]Ֆ��CD�<�$��1ƝfFj��𳁱s��G �jD3���.y���|����iG	8������$+��hq�l�^�d��в��j��<YD��{����.�l�TG�m�� ���5?�����.��zDj�rК�_�T��.�t�[�I:��DA�JYsEw����X�n19��<ƯF}���|�`]r'�0��E8�hŪ��6.�?>D�%�Z�(r���,��P+�i�q���ۚ�#a?�z�/H}�(��(�Wm`�s������@3>�h0bfP�A���rK��d
LW��Z�<�L�[���/%A�+���*Tٯ1y(��9�T��j��i]�[/�`�JT�i��Y���R6B㙰��4D���i͊M\IY���֞���i��i�Ь�Cy�.���9�
�%��
1�1��.'"�/�ui�s���W�D'~��w�g���I
j-�ص M�+��)fɍ�[ʯ��l����xZЁ�����a���S����n�?��������*~6��-��?��Acn�6	R���Vĥ�#o<>kP�������`�fH��2�ɻ�6}n����y�G��*��Ct��gX�C�߈��I�&�,�\d��Vx����M�k��@3c��햧�&��<UhѮ�����h���P!��<3���,@��3��u�U�ޔ��⦟χWޮ`���Ȏ׎1�튔��� \v��k�x�X��|+!S:�*�����!�׶�G��5���)�˻��6$_^q\��YK��D0�~ʊX� ]�>�ʷE5f�;!'�s�}�0��o������T��=�y�i�������e_��N�I2A�-ID�r���EWӧ��"�fiG�֚X���Y0A��������9�{S=δ�1	�Pǈ-\��m��'�����8d��1�k�>1��{�hØ7m�E�~=�(XZ) �iɂ^�=⸡���/�u7u :\C^۾��Ћ��W�Ӄ���`j��u��Tp~J,X=;(��G�ZaZr�	���?)�8�[��k� �`��o��'�QYH�	d��<BTb[�#鷃�
M�7(����­��ì��:J�W|Z�vR��P�;='r�˗+>A�®�g�Jq�Qs�ƭ���H�"�{��k�(��l)o�z
.�Mke�a�g�������\^?�,&n����PX)2��B^�1눻���R)ڃ<U<y�r�����p�%m�́KtNN I�2[\t�	�})�Fd�䌭�$8e"� x՚(��f�� 9��:ތ�5���Rw�P���h��L�B���൰��9!��2�E9���͍Cq��8�쉄�����HD(l)�NP�ʖÚ<i�}�7�B�ɒ�iab��	���G��\'�n1Ф��.߱�.;������I���n��?�/�z��RBd�������$XB&q�ڱ��Ⱦ�vw9��� 3�u��G��y�<��~7��2�PȱY�N_�߼&��F{H5���~L:)V��+����fw���^�%�f�l|��PZ�b��&�]��`8���{8'i{���i|��i���@���&��!��S�|�;�9�Z�����4S�g ��غ�.���=�8�Z�JB+>��*�ŷ�KW�Q�sO�Z+�L��dը�HVT� �FT��L��Q��pV�a���B�!kq�����8�E���ԅ�p��4��l�i�d��&�	�ޠ(�祊��Ѱ�N�\L)�Xz��67C�Ȏhy�=Op�7�N6W_9 �#z��K�-��RM���V.Ա#��Ȼ�|����f�+HEݺ4��L��F��m N�)4
7q Ȯ�w2U�,�!J��8#���<0�D�4������\��)+��<�=B� ��9L�?��¸��V��`�X6�����]6�-ߣ)�!�hP���n��k1�e�b�b$��'ZZa�{���ڝ6��u����Ȩ���X�XnL�K��3��X��И�#�K�-G���O�2�����$��b�m��կ�����q��	�58q��8�L��%�c�B{���Lh���F�����TKĜH
՛�Aّs7e"9�c�M��s�[*?(%ٶ�ǫ�ޢ@1�������ԃ'@Y3�1����u:�|?�W�jl+���Ͼ~ڀ
I�v3����6�L}̔@~n���L!h�<J"n�bV�#��kHjJ���)�R|�Dg�+U�M#�\gt������j8'���?��J�>@j���q_DE$e��
 ��|5���!��G���V�|�|��p(��jӥ8{�~�d� H�������!壄�^�x���Ő�����Q���ɡ����y�7�r��tA%C��E�i��c9K��Z���둔�磀����SC�*A�
�/�S.Ht�)>=v9�)����
�*ɋϐ`��A�<�$�H�;�U�{'��n�1���)"���7qݳ��m裚�u�M�Ѐ>��&fՊMƖ|6���3�j���~%���ҁ@�k�'�X7�R0�O�C�t�1x��P­�X��
����7���[�V��s�
k#�r�Opב�WAM���=4]���{�m���@&n%�s��}Z�O�c|O,;��`����-2��Z	�a:�O�;	��&6
�/9��C�X{� }����w����z�d�|w��	�됧����1~��LC�`�SE:JN�g�����E���B~`ףիY�	!�L�"O�K)_��%rU���*�܀B߉����;�/�5��U�˧
�?OI�e>�76�YT��fՏЉ�22���}�wmo���Vm#�ɠ�����Mx��I�BTo"B�ɵ2���kQ�G��(�Mvf�]oַ-_Ծߊ�xۤ9��(���g.�J�*C�a��|ӠJ�/*���W-$foE����f16�R�Z~;�k2��UR qKM1a#�=��m0>/\	�����Nլ�h(���Y[	�f�'�69&N�ń�\���
Wq�G�*Y �����(�C.�U~
5�oǢ�UQJ3�x(�+���@�1bqo�.�{3L�?�2a���N��8��V�~E����H"�.�e�.UΝ0ݫPpއ�;;c�����Ӱ$��Lf�f�I�vu�C�Tj��Q4��IܘױWő�� h�`8�5�3V��+g�?J�|� �A�	.Wζ�,�O�"<�5��{ˠ���ͯWQ^Y;�l}���ǘ����O�zn�a�6+�������f	Ca�"��[^ѣ<��oxi�.'�KCAVw��S�9m=9�^�ÜSz��H���g5̮��X��I�=�� �P��g�`⡐�Il� UۖR~r�;����p5��� e��<�K�����.j-���aHSW�`o����sU��S����#q����l�����\�y����+� x�j�x18v$� ���p*ɱ�%U�N�F���1:U�+kUd/sA`��Q8��`��=6<�A5ț-V5���-��9�n�ʃ��X*p��C�A��{�H��%Swb�ӥЀk^���?Y�����wV�๺F;q/uO�%`N���;��}�It;MC��&G��7q�x�{cTe!۲���:�U����!D��X�8`A���k$����f�+~I(ok��Ѳ��0���_&��rD6�|��l2�MO��{��6������{���Z��3��>_�A�XCK	�9~K�i�0n�3f=�!�9q����5��I�j��נ�C����f�k>�B ~��(�P��ꔩ�F/�������V�Q����8%�u������T���^(A�g���g�O�t��xC�4��x��䘐�ܩ��].�7 4�ۆ���+!�'ЃP|���Ϳ��%@�v���P.�����S��D��~?��w-U���\���I��������B�
�/��@��|�C��,f)��W��x2�O�
>���3��
�lI��#�,rk�ИZO���e�ϳ<W$�!�<c怗.6�A6��q�[�6B���L�Eu_:�D��5v�$_t�H���:Yts��>�"�>�W�T6����>��:�	)��MT������* 0��g�V`��-��݈-I��~Դc�ءW(��mBL�H�d�Eyʣk�`�|���s��"��ۗr���O̔E�ݠ3x�;��1"7v;��Õ��ǧ��9/�H�CgI	YTh2����!(�����,p�{�N\9���T�Kc4Mz(��I�z �DH��B�pz���,�ww�x�ɏ���e�J�9#�����
.��߷���}!Γ�o���C��
S������ey�����.n�*١F»��-��IJ/B�U�]�NWc�����]��t}'�n�uJ����-z��K0��0;���yF��c����g��_�HLtҭ�mL���+�\�ʙpV���� �� �Y ���:��'�����@N�o����Ͱ����1�QŌ�9�T��{�)�;U��޹>(]�:�،k80�K�F���&Z��ß��.pK4�D}�I���O�0���O^���/��m�yVG��s�v������������ٹ�y��]�]	ū�=�I5��&<�ʔ$�����+���mWA�cj���`� �G�=,�(p��d��+ϕ/b�)���_��6��;Di?��C��P�0�ݦU`mu--ܢ��gY���n��S��e� a�G�J�)�e�F�>�[b��P�-��^!G�������r��^�}s��4Y*FI��qD���b�`gr&jzL]Q��4���zͮ�Py�!�b�	��I)�w���w����+q�|!7gDE`~㱭$;WxlX<�T�a޽��� ��"��/g���?�釢a������_��q��&����Z/3O���A���B�+%���W �+�`�o���g�,� 
|(�S^W�ɸS�S�0'T��wkT�.U��*�ޱ�[@�;�(E��`�
�T�ᱵ�b8؞��;��џ)��ɸ1�:��m�*�s�-�Φ)�P�m@!�[H ��n����{��Z=��O�r`)��9hN2�o���
���6ٵ�;�0�E���Bscid�18�\O�F�ݥ�-�������L]�C�w�:�m��3>T0Ei��},m���۠�00s0�(igz��n�^(7�Ŷ�)2�:��y��Q�OǎL�!NIuC6w�����*�������ಙ<�Q�9�l��Z �w�S�Z�K�a��d�*�7P���sY�#�e�ۤ�d�y��Wbr!M�#���"�4��+"(�l��o&�����ɡYs�E����ߠ����lv$č�w{/�U��(�C�\jq0T��= b7{�CX7C���Z�����`���&���Z��
�El�4�z(�	�,h�|k�X�� \^�����S�Q1LD���9C�&�/,�E`�Flq��i��#��ۿߖ_f�=�hyƖ�+wnK :�？}��z����Nӑ}�:M@�0���1�)OC!��X�&�8iH�k��J"S�P�&�j _\���<ny���k��A_%�Ё��[�o_�YҊ-�N@qy���\��Ew߇��r�B�}�ɾ�����1/�L֊�F�!C�wrz_�RzM<�o)e;��M���L�Ć��1�]��e���n�~�<�x)�j+�O?i�)���ۙm��6���o���I�4�`�`�xI�$��]n����b�r����H�q�:�qL�i�J ���4^�'���f���c;�������c��"�y!��0�1�ŲP7	�Q0��\�*$	��s����d2:�A]�%�d���qʦ;m�Ey�~%��":��yǀ�����+�g��F
�����������\��[Aހ6������E�1Q	( ����RR�/�?�dC,{+7\?�S޿���C����OX��!v�h/rgշ_P�Bjxh�@�j��k>�F�O�ՑD-��Dx'�Y��4�]@�ہ^Ⲁ'���0nأ�6O���_�NkN��&6e�tR���x2�&פ垃o�����?v
1�;�۝2� l7?6Q��x�r6���݀:"bɜX���	�f�18�v7/?��ї&�m�\?�� 1�?Ղ�I�m����ă�_�-��sP��,J��>���&ʜa\%Y��=zFT{'hJy����FR����H��P�H��.�?�j���OI��������Ȗ��W�B�:s���w
�f�ݣ�D��X����.�����=�qFN�� �ĺ�oR���g�Hx����ـ�S����fڔ���Q�?3�IÍ6��eEl5����ٿ�!�F��vk}�Z��_	j�Q���|��t�a7���0�6�E�o;%��'�>S�h�%�S��-q�NB0L*���'��4ک}�{�. ��N=ּ�^��չ�þ��f�Ħ�}/LŖD��j�X9��]�(~�C����p`=Q̫
^Bn�ɽ�A�`I|c��ÏK�����[���')\CH"#[���%�'4��U(cw����ݳ�5���G�Z�X�'�'G>���誙(m�UL�R��{��u�\����bu;�Q�J���V���*���ٳJb�E_B��"��}�1�ud�Cp���Ώ��cA}�p��c��C�yD(;6)�|~%�'n촼�� S���
�J�8�{��[OvN�����Ъ#S��Ƒ{`[?��^J��ɯ#�I��ǌSL�F��&���xrK�=1 Ez����2����(��фt״:K�ZYl���9d�M����w��h`*�t��&|�Ug
ߋ��ynL�{���ڣ.���[6s��D/�ۛ���2^9�zQI��.%�d�)�+��� ���R�+�w,g$��Fj�v~!�4/Ú�-BD���*/����<g�G����Ʒ
�	�F=4+�v�Ϊ���v��,D��޼��h3)�x�Ǿ������ؠK�!��!w���x�k��7�{=�17���7����˂̽�k���U��������bir&j~Ɩf��;�ve��Xy5���*�h�#�#,u�Y��{o�c�d���RÐ(o;���,���8jK�9�(+��sI��1���N_4�߹1�L�hRg���Kd։��J�@h=Sg���m����Nof=P����}k,��~��Qit�:���K���=-
� �((}�#6����& @u�u'�Gl�f�,�H�f�~��%���~<�^�s�	�'�s�9�J9������F"(��N�� �pWn0�� MC�젶�+���Eה��I8a{�3���Bލ�6��ஓ�T��LA�`\k'��ѝ�������3|]$O�9v�r��/�j�����Rĝ�w?+X^�>����kѐZn�z���׻�؋N @�{G����{o���(�]�f�PۛJ\��Ϲ���*f|�/�Qb��X���zx~���EI�Yc_�K��(1����<SG4��92�����c���c�A�Zk�~��}�!L�=Wp?�@9�A�����7oVTg6�Lt֒�m;]Bh��RWd�E��햾�o�}S�@i�'�-�9��e�/j���5��>����Ѕ���jCO�Є)H�{6{:y�x�Gi����f��2D��{~���zB���k�Tdg9"[�>���c�m'�J����}v�[s�#ڧ���c��F��wR�����	�Y��z���WQ9�?�Q6���61ʓ�vDV���zߕ{_��qJ�;����^��;TC[O�
OrHH���O��U��hyX�`lr�n(v��!���X2ǜ�~k��U��,���l����.b�cu�n�E���BZ����m����J�D�I���~�ٕ���ϧg"5oBw#�OܑS��j8]�X �cG�eB����Q�V[<�;��M��$Lm{�X�����fK��k��Ħ� ���7�ZV�
a(���n{{B�Qͣ��u�õ ^1��Q�wֈse�(*e!�|���wYщE�X�l��ij�Ox�C�uEf$%�-�0�b2 g;Se����a�d� sH��j��474hI�H0?�x��S�g!t h�ġ(�?�o��S�����S�#��;����x(>���D�!�EN֦�*�&�y5/Y쨛�r+]\�=��넜U���V�W��誸��O�x0��wZ�0 ��N�4�3��^-�w�LJh�I�̺I���u��C�	u^l1�?���Qn#g�8���6(�]�@&0�<X��9|���O[j��m:n����YsVb �9ހ��2	���Ng%Z��1Wq��w��b����\�=���8�]�����VD֥�]���~���}uQ�3Z*�����ŵYIBN�Z�c�F���Aj����ڡtx%o�]uhSҼ�+��B�w�B dc�����|�c/s��ZQX}����fV�E�0ژdr�׬p�ۓh[~&/.�4�d]�
?�CwۭO�;M�cr��	�k�����K����sF��L�!ta�)��ȎkUT�'}������ c��5�����FfB��D}��m'�|���E@��������b���Wd΢�`}�md��,�X>W�@��y��U�D�2n�:�{*޾&�����8ٵ�{���p}�Z�yY����ivr��P6��L��]�1����]չ�-$9�_+��>'8�z�~�!�u��f�c�*J�^ފR��"s�3�����0���[���L�X8��k����n{�깇cL2e][�M��ļ���c���\8�wG�rZ������ �r!ަ�����Ć�אs{�x�U�n,`]�Hݤ��&��a�~
�#8��)DQ��"mh8b����Z�KN�S��-Z=Q�f/��\_��n�����w��{���+y���_����ZԬ���XX$ީd�I�7� �)��6h�0�)D,�j��b��{�Q+�ԭD���q���������E�9�<�u��e��ņ�,T������]�ͬ��vN&#"�q"!��Q6W[��î�]��fL���))