��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CG�ʜ�S��m����un�%o׎3ke����)�ˡ(c	��&}I��>�!�-��@bRH���$ݍ��tVǆ���2��:^�T��}��S��g�2Y�ܞW�L�kB����Y��B,(L"=�񛨿${f��
��.��C��ÿ�q55�ǎ���N��6n�-���i�E�BES���	-�	BX��O,>_O��ńD4�p���pǱv��]��C�;�sܴ�,}NL�����G���+���Ọ�_cq�煜�����R=�y�{��A顃9b���RPʲ�;W�F7���6Np^�A��˛��"��5�HǚX?�#�ʍ�]��$�ק^L�`�ó�XWv��|�aV�F������`��E%�RT#]SG���sǞ#i�E�T�ͬ^`B1��Z�=�3ﰠ�|��i�\��<+����0��j��U�Nd��o�E�����Y�
/;P��zsҢ��{��i\��\A�ھ�u��^ik;_ޕ��}��eo��H�K��������`_a01�6��YI	�ǹ 	������Z
9�kR�������lOK�$��=��Qԋ�r'e�}�"�,�}k��Pz U%���'�)>�����扙(	���ޑ�U"~����WܗL6�9��##����P�3�8��)�'�#���T\�m�O9M��K�ؓp�.��G�.�߄Ce��Q���{67�����Ї�^	�3J��F�J@�8�����xǽeB��	�uq�J��E���զ��ʛ�N���Np:~"`䘾���������ۖ
��%�,�I��J���S�%1A���t \p8�\]��T\h
�]��t@�݉)E<X�n���띰�J���]geI#x%{���"�Sk�Ơ3��x0c[��kt^����O�YrΡ��\_;�Z��N�p��0�b���	'K�]}�G(��	�H�C�J�+����"�:��n� |�)�9P����f���|{o�o@�5XoB�!g�y������6M���������P7�Q�{{\�5wVW�P��mдx
��8l/� ��:˲�s�~�|ы�[��T��S�x�P����G䭭�g1�v��y+H��N������T'�'�>�oH������j�N�-L	��:��|{�L�?O��$�D9���vy�ք]���Zd��/hc<�����g���c��P�ؘK�
r�b�2�خO8 ;���5��zx:ʉau�aW��}kc�>y���pY�VH�W�
gv^Ѓ�_��#��p�*D��s�&S�:�.F�\��᧽|��ICud���փ�(i�>d�LߟM�]��@�ݲ$U���V�%��D(\U~�>���<��\!C��0b�Ϡ-6A?}G&�q���Zn�:N��>f�J>��;# b���_ٌѷ��r�>/�^F���L_��F�� lN�K/C��(�[����h���q �i��*���@�}h��gX�MA�>���A;�3A^�>7��1��_J*(w��˂�������	�1�O� ��f�l���#��B�&U�<��;O�y <���w��;np�� ��[�~�\D�l�Q)�뤊TB��р�_��Z���͡��Y�Д�q�3������q;����0NuR'�Π�Τ��Z%���̂&҇"��B�&?H����yh����{0��A��Shvv\��A1�-�z1oƩ%eM=,�O���=��m-1�zY���]���w�[m�L���h���/��������!���8�6C�����؜��%��,d���2�KEB������I}��י�i^����0��P�����2Ш��3>20�]��uL�� ��n[�y�+�A�I~���Y�v�&��c�4�����=E��D�6>�΍��x��E5����p�n������ �P-�X'h������Q�j#��g�$/�&j����Q�� �1]E&)�!�t������*���!8�L�$2C��[v���UIw�C���3�2����ڤ@�X���cp��q�3��f��<d�x!T����CH�ynH�Rh�2Y���T���?rǽG�:���<���S]�28��,L  ɒz��F��w��mƻ3�V����Bb;:}8zi��O� (�`3L�Y1.�!��h�e�o�-��>�S�R�c.k����iG�t��F��~e���W�:٬�]�P� �o�v��yv�ۭ�3X�D��[ne�&Ƹ�4�\����TBZ�
[��j�/��/ddh�BOP���������ًn6����I^-��k���'�9���W���ʎ���Q�uFG��a�0��chĭ��ںi`�,$�eH�N�&�/+����_W��!Y�B��Vm�tly��f���f����U'ML;��<��L�I�k %�*���9�cA�Q����+8=cgb��'����l;]��e?��4ET�z!���J��A8�:m��L�6O�@�uמ�a��Ě�(秅REa��h91�zmZ<2K��c�mK��Ps䶐,3�G���0c�~ei�Ƀ�3�� r����_��pv��&*�.�;��N4��I;�0�Fy�T�P��]p�e�DX6�������]��Pp@�b����W��f�u��x��j���l�sw1�ئߖM�Zp5՟ Mf���5�\�A�᱇�k�n*��_���`FѦ\d�8V��SI����q� �������>�XF�ڽ/@m��z��N��9����.
s�bp�KkN�D�R���Q6�yNd������W´�&B�V]��yt�U�Z$Ų�X�@S�*���W�g]_8J�nt�8� �o¢�{+�p�7��Bm
��]}B�"z�ָ�y!,=?#@ӳDYy�4Ҽ��BU��]�(C�:���洭=p��t��R�UH�M<7�!53Os������J��DQ�d^�rR��<���"��r�#�5��Z�R����CC��R�U2���0�j����9!��I8o���n�?�?�s����N2�n�"֬'����!0���!��~G��AjIޠx�{�d>5�:L�xh<���+xd+`ޅ��J����#Y	���b&E!��P��hܽ3s`��+d�y�2q���z܊��;��O5�fѿ���w��g7��_l�dV:�נ�@��J+�;���{6該��e�P)�dZΰ�M��f�b�w���j#��?�h9<����ł������ ��� �2ٿ��W��ev�Q ���be]�mv��T����	��2ŉAg��5uͳ�n�E^z;IJ!�>7PJ�Ԟ"�����F9�ш)�e1F@� ��#�s��bqv��)�:��6@
}u�V��r�����H���k��+䢨���cVDOR�y����{�'B깭}V"�ڱ���Ω���egE'��k�չ&%?�k��X�[�;2JD@#TY���4\0=O�9�?�Ƕ�bx��^vJF_Xn�'_G���u���2��
���5�dW+??���S�/g�V�R�4�4x�&���)�Rc�H�8.h�'Ts�����E\�3���l��J������E��b���20S��&蟮�w"zm�[OR6@���'^1��-zO�J"�w�9[S�"�uB��l&�x��z�
���g;���K�ۋ��ζK�w���R����l��|�����%q�U�	U����Zd	Pa������R?��M�w�����m1��<	%�tPp���z�^�R�z�wC�q��1��5�6>�!��8D1�7�x��=xje�A��u�oO\�Ǻ�0M�O�]��L�=�Qm��VSUl�KiN�y��$S7�*��D��.��£#�3�
Y�����x�2y��(���M�+��0犊�D���{,y��N�Ϙ/�%7K�͛��I�qODѯz�:����?+Ʀ ����6Z9O�ީ�&��P`��u8T\��Щݢ�I��u��4fA9��ݷӘ1���f�[��"����9�_4��|���-}4)E�ך|BR�ԪAF�J�fJT�����,ɩ��[�7CpK/��vO�$`#Ү�#�JP���R>Wlɘ�b�H�$htü[��C�n%�=��q��ݎ��*�>��d��^^M
]���ͫ���^._�	E6g(����]n������lHڏ��K��M�d�%bF�"���:�QG�o崓{G����'����n7�g����j݉V��
vj��=#�A���K��ٺ�9v���>?�`v�)s��*o��)�%�6솏��@�(���t]�JQ�Mڒ4W�[����<���6y�̫�L���ty���}N�ŢP��fq���Q�5�&���Sax1@g�+��O����c����΍�>6�wE�����2D[As�"��;Oٹ��U���裞]KH�0i�1[�mS��M��@y�'��&Lز؜H"��d�5g
�BH�P�s;��������y�z�t���ih5�6Q�'�IGD}��ٗ�����M��d*p�Yh���O��2��߆���c�젭h��ӟ���0�1-�sV+n�2To�R���n;��a�f�^�m��Ň��j���ĉ��`�Y�)��_QHˉO7�t��4
s�6��]	�ɽ�-�д�C�ێ�Gհk�s��>)���"�Ƽk�����\��o