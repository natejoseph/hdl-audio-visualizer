��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ�@o�G���D�t4�M0G�R-(�`�1g^��rf�מ]���`�?��P�/Uj���/����`�
iW��'l)���Z�hމ��9n�h�$�� ��Ϗ�H�F��柑L��}�X��Z)7F�� �D%�?��"��M�˥[v�2�9?I"á�/�E�Ky��g�G�L��'��N1a���̀���OeU��ٜ� �a��`X�5dK����Q�=B�l�8���UZ' V��ξ�v{ҾN,R	~IW�9����Bƫ�l�tj� {�v}�B����f�Z�_�r3:��p�hJ��E/���hꔜ���D�O?��%�7D�L�z�.`��E�����Ճ�]4�����F�ՠDv%�T���Xp3 A�T��SXBX���R4����P�t��%ߤ_��x��q���t��
��Z�_))`y�p��_�o1�{'�B=HtY#Es�̠*����(n*8���^+2�c�d�D��s����q����P��3�_@�3Fp)�n�p�I�s�F�?�F�[������n�,�%�Z�$�\}Pg��M:��D5u�k�EB�a��3�nQbyBt����%Nİ��Q7q�����?���."%M�r�܄�.#"S]|��'�Q����I�l��i�4qq��q~�ᖀ��`�/Bѯ�R�^"���I�.\d,�vgO�p}��i^Ñ��WX��O��`K ���y�O��i�E
���$î�^?:��Vi�k��K���acQ��@i�+A���s�����B����7s������'"2�E�2�����O�����@�r��J��ݳ�֏Ǚzi蚞�kMǔ�V1������@V>]!�a���$p9���n�ɵ��P�<[��k��R��O��y����=!��sBf`����Xp��]��e�4���F8U�[ʂ��ْ�3Ÿ�S$tmJ�D�&v�{;�����b�x!������O��ՙr�=aR�㯮X;�+F�7�"v���Z�+�%���TPF*1]~0h�+���x��s�\7�� Z-�,�a��&k�	C���/�a�-��8�>6y�:*M�|Sc�Ik��*S�\IZ� T�[Je��X���������R�C�}4�x$E���5�<����1��?	��9�ʷ+A�;�Z��h����'��cE��nB�x�'z���b�X��5iE��HNF�� @9�Eۄk�=͈3�1�l"pj\�x��P_��@���k��;���v����i�)_����(kNe2���k��?̐L�)�����[EC�6*g�e��ג�e�"�ذ�;��!�6�H��E�63~��J�&
�O���H_T�C�ҵ�K�G�v�@[�0�_{�\o��!�_40Xyo#��=�3�{�y_9�)���!�ƣgx2ҳ1�p�M�\����ƹ��*,�s�2���B,�le�]eQ������)��X0�:���Wdǂ,�'aRa����	g =9���g��#��t�8&�b�/CP��,x��JgH�	@�|�����W�{��E�F�Z퀜P1������V˪�$���3I�(k!���$��UU&e_J-I��#1�j��B�����Pv�i]�x,J1l
0�2�7���ؠ-��|�C7UD��ȁ���H/�﬜k"[���Q�&@GeT�N��r��KuKDN�A��3��t�8x9RJ��|�&_����GR��y���`dC��KHY��)H ͒f�׎8߭�k�q�_Y���y�)0�v���9u��D�cτT5a�t��T/Λ�0�IbԶ�](${�ʱ�\B���[-$ꝁs[<jYEFɜ�ن4�d_�jl�<�X���|g�&����|v�z2.K>�l�Y��З�zy�,dZw��b��LCw�Nz�W�]ah��2��b�j�3�+C���q�"?/j�I�٪h
�G���A`����R���sM+�`���N�K�����O�)�L>ֿ
��?��:�\A�t3B�f���h��)@Wl{�E�b��{�辬O9�8��������wjw���|m�|]�gS�_�v[FKB���t<8X�k����2T���ʎ��"��{�2�<d/y����սZ��q�+�� ���WZ�ѱf��M�Uϵ�Jgi�f�kP$������,��o��'r�øp�8������v�2S���� �$��(�wK7�FV���L��'n;�ܬ0� �1j�p�y�r:�,V�׵@�w�L�(�� L�,�]��u�Lb(��hl�l$�s����gT�V�B�4Ų�x��`	�p��n}r��S������ ���W�*���mH�66a��n�;.�/ZI������n�a%$�ឯn��u�ụ���9�����Lyu��a�r �X)C� O�M��9�iH���*z�)�9��W>���a;���-�� l�������C�0�����
���OCorʊ�4Ы�n-��Q=�H��w\A)5lST4M�1�Rm����1�mC{i��@g�! ���w�l����s�pHy�GE ڟհ'@��i.D�����c5�rQ� ���W+�� ��}�To|�0�qI��]�f�l��3��s�� So�%w��+Nl��Rr,Il���$H5�ʸq
��S�,�V����_�78�6���-!�Y2.��������B	S��5�Ys9�� x�FM8;e����Ϣ%M���j�/y�td�Xp�Y�0����i�nBKWw�ƪ��%w[
2`��'PQQ, �e�o]����|y�[TCpt�9VY��h�����W�0�Ce�9�`E.9���C~���,�B ϮN�8��:쐬�/w�Up�����	�eP�O�g�����-�;CSZRf�	jJ�i[aB�@������|N��(���obX2O
?&].��Q4)��54�C~᳤�R�M�����֦��~�/1�����j,\Eٰ��$Le��5^��|{h{6��>�.��x�f����*�����2e�p� �	ӗt72�O��;t=�l��Tί"a��y%�@���{� ��,Aqʓ�آ�n���'���&3����b\{cZ�$��e���cawd4�eƩ�����'��Wǜp9+��VaǗ�v�ϊHyDh��������I���	z��fܱ�9�n���ˢ|Fl鞧DEy���5�<� C�U�OE�����龟݃��Q��.�uf۪U������6�wb�[�������w,�eԠx�ry"W�˙�,�����3W�u&#�X -�j��v۵�V�N�ጋBA�j��7	�B<����vǞ�RA��A�Ђ4] vʘ3�x(h��ۨ�p��[�^�7�Bc�ud� l�+�m/z��˩O+	�5y�v=��i��� �8�Pm{�$\����qL�OO���f�>ܜf� �{sT�B�G�Ʌ��W��f���Hر�PS���Ǳ0AJH�2?$����	�z�)!��J�=w��`N[����)Mt#�ÒjK�k�e�ƳK>�爳��/rp���`s��Q��9�ܩ[
��>"���-�a�����k�l���l�>���S:�ZK��r�Tb�BO�-ۢ��ت��<��'��3�Pw�ڭ��M�p�ą]�U'�Hs*�$	|
��L�1�JC�r=�i�Gil
̰���Z����cCJA��D�Ѯ���E.��R�z����� /��(�1�wk��]�m�&K�ih���Z�6�\�+��j7��׿ƪ�-7��!k��B�o��a�S�aX\R3F_0��r����
�w � BTYw��a���j�ѕXx��&�A�qwQ�5�лێ��t����$�|��3B�P�.ODhZ�����>`��|"[9o�}�j��˽�.H��5Ȋ	����sP���{�_7Uu�EʣEC�0RL�N{�@��sl�\�f�t��l�L�q��3��FE�m�з�|6-V��%�
i�oJ�,*�aiU��v�8�'���}��P�)�������Ϻ)��<������2��<�n��_��Y8`/No�R����g�T�}���G�f���!6I(ŋF+c9`Ͽ��a�,�6�%NFR�)+��-�N)��h�:���f�8>y��ҳ9��SH8���Č�tVO<��΄=1��X���U��������U	G��|j�!R�� ���2�A��Dz�' R���s&�y/|w�y+��j��~r�h��n�G����l���1�&]*���q��"ݱ쯏g(������!R���Z�%47�zE�Eȳn�]�a����AȀ������8���[,���/��"W	ۤ h��E��lǛ\�1�����\��6_������N'��g�G�Qm�ң��v`u;�FH[�R����6�>��?�v����U:h������Mf0�h�*���A\���lU��܈�z}�I~�� K���)d�Y�	��܇W,s���\А�i�ө2���$�(�$�g�����?��1�o��6D�2MH����K�|�T�W�Zd5�Ú1��E6�H��i̕��$����R�����A�¼�
���5��L'���vu�2>��"���D�}�IN�[6��̷�N���͠*D(� �0?Z9uk���2g�>-�*�_�v`>�$�Tħ��)n$H��\���h��0��r@�n�����2a��法�Ew�%ۜ�b��RO���'�þ�fu��{�e�yE͉3�V,8�ڞ�a,Ny�Ԁ��ɷ��y�I��i�d�5�*#F�<����˭������'�׏A�ǋ��}�oIc��rF�u��!�	qа��r* ����_��=n�A�똞W��O�	Nѩ�%?}�������0�iʊ��4Yм��*��:e����~f��'lG/��m�D��4mw�a�w �D[S��>�t��#	(1�ҼʍtB���	�.z��1��cWu�v�W|������֘v��Gu3q�"p�3�8��T�a�E�p�5b����-��aF�����t��_�c��F�id;y�ܱc�u�[�'��d#۽�T|�P��O�s�yU�"ʮ�.�eR�eS�D���E-�JA��������ku)��J�	��8�3e���6R��J�$�ԚE���,t���� 5Χө�PEQ�K�1Z�D�<��6%YS�Y�pYF}f� ��/У2��?܉$x�����鮊�9mj[��]s'5Y�C@#:����m��2����R1�(b��/X�C%$�A�	羾	Lvazvw��P�M��@��'���d� Zg	Ӿ�.�臸Y0��)��rb��$�r#US��� B���6��P�:@�A�[7{Z� k]�?��+����!+�Z ����l8�i��u�E�u�Dr�=/x<;�w����C{}@�Ѽk�Pm������SPoL��oD��Q����ߩJ�,�����'����_m	{�q�Gv��sMR���tU-��Ҳ��И�Z..���O��o�3|�Ъ����ϬFonb2���ސ��'�:M�l<[��Hp5�'�:�*����j�bE��C��dB<�!�p�ɝ �w����������e/&v&�fvs]�=�8D��˭]�o3�V�|Bd_r���&{�;�퇛��}�!C�ժCڀ�ѥ=�����0�������$�j�K)n�O��C�.�|P�*�ԅ�>`���[q�?*
��E��������߱���G0a�F��⠔��'�1�=���5����q�+?��jw��	�4�U����kĬ��?扳����a,Ù�T�q�F���N_����*J����h�q�$g5�$_�(��|%rЪ�}!�M.��;cȭ���6���?]����f��4�
[�u�X
z������L�hH��L8�Eb��-�<g\�eڑF�:*-ڽ��߰۱���N���H����<c�V�i�z��Bxd�C����20QR��
Z�D�j�����P�9G\(ς��ɲ��0�]���	 ���*�'U���#BǏ�)�x��;*_��w�(#{�j.�d�qJzȜ�x0�e�@�z�:�,�Y���ɀ#�� ���w�ԏP��-oT%�zؾ�yL+;"� �;��پs�PI���O�MɟL�!3Of�L�w���4���~0�\g)���Y��Bw��xV�,J�z�ӜD�wJ2��ƚX`��b(�6�=������<�NҺhtЀf��u$��aT�ؙc��h��|�
˕EUR�7��|B���K~�x	�L�a�]O��{
P�H	0�Oj�Μ GA��PQ<�f[�/m��Q��JB�bղ��	$��\���}Zz(:
$�_� ��=c7F)ن$��k�)դN���u�M�"%�� ���.���]%��#�Y���P�Et����\O� `n�BM(��k~�u��z���2[���n"�X\2xG�@<�;C�G���,o��cF������|`����g�׸YR��
��TM�n�V�j�Sb�G����οo\m����+�'�ccO<�K����5���s�ra�`.aC����n�@;�	,�Z���\��2�:���lĭ�K�px�Y𢥎��(³���Ts��@N8O��Adَ���RZ�T�z��h�g��R�"�|Xv]���Y�?Z���Q�Ri�Kp��)d�
[�7�j��͠g'�d����P����ʮ7cY�LI��by'_��D��uz|[�z �[�j��:���&]X�>��$���|���N�G�r8�iBf�\I�������8�V���i��Ea����u?}��I)w��䣥shZ��ĕ��K<З,!
�olr�,Ͷ/�'a���i(�헿�����scO���%Ӓ���N��o��q�O���u�o^[ �m���H�֑:�;?�m�-,w�u"�7��N�*�����w���;&�P�`	�-[>c�w�8b/6�j��?;�	���4��"�$�&�2�Mp����F�>]�{�o�1l"١������V�4�\�]���'z�KgY��u�5�#L���ͅ�Dڥ��o|�>�Vģ>HF��!s�vA�H�\,��b���N�U��\���uM����xsT3�ա���#N �F=W�!�[��O��OE<��=�Q\��W���!��!�^&ݛC!�׸���,����q��ѹ�G8�� �����i�Uk�Vk�7)�P��� /#�ݲ�x2Zh�Q����;���[��=7	ܫ;0��7;�����!�I9p���k}4��Y��th��$eNu۰�A`�"�{��+$v�T�K��җv�����K�<�ϵ�����uN"� ��1����na�n7<Ĺ��_��L�Ř�e%�1���Ԑ�0R/�)iw�t�I5��tW���۲�H~R����f"�u�����a�~�Q�������s�^#�\L��6�L���G��Rk"M�������d���v>�o�#�r��(��ݔw��vB�G3hӅ9�5踋