��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���֚/�뤕:~���.�>*��3x���{"=<�������b���*p�Л��u+�r����ߞ:�L����"W&P:33��+'t�%��u��T���#�2�`c��m2� �
��v>LE���D6�?��@�a����F�1�
��vS��Sl�t��`�)����<� {�e<?��9�^�V�SG_�.@��n�:粀r���G�B��bY����P�N�:D�������(�YsF������~	�W��DL���@gt��Bq>���܆���E�"��;C
ޢ��#�t�/�SDK�<�*=
��x��ˑ���RU;��������L�~&g���7�>E�LW��>��c�Y��ܼI�y�<�OO�\�_�� #�-n��(�&A���m'r疭Cov�~�wC�j�*�)����O���ߵ끇��$�!��(���/&^���U����Dg����ߓ&�:a^�rQ�I� J�k�D����6{���+��b���e[�E['o���`�H�@�Wj��+g�d ޻Z����%A�t�H�3��	m�f�h�!>ˍ~�Q9-Ǒ�6U;����a)8'L�)�T�y��J����|�O%�/�ؚ�5��RmJ�wÊ�G+�*�V�*�y��dÞ�ť�Z�>zI��{YR8iʳ��;��w�o�����B�d۲kB:f^��¡8����}�	[<����H��H��[�A~��k�]@mI*X��Z��$� �������ͯ��[?.h�1.�<���b�3�<���9c��H:W�ܾX暄�C`{�9p�B"��E��0�4�2����~IJ��]h�/�����T��C��U'���)�$*ЪD��k�X�.	��L�' � �\�k �����#�t{w���3������ލ�W��^Hƴ)���Vl�_ɔ2����Ɍ�3�G�Zz�|�@E,�����i�8*�	|��٤� �
ݫ�6I�XP������jL^����݈�}��&�NM\g��s[P�������u{�����y��2�|%_z���qwT����s�� .���C9|��X<��'���b{�#���޺f�ے��=�H� 5C��xХ�m1����/Y۫��t`�b�^$����)�^�n.r�hE���������}A�a�K�B�p��t�k=9�^َs/V���p��x%=s��/����Y�����Ol�p�I�~؏���-�Y/����^����Ǻ���A÷�<r�).�hWO���,�멑��ꅢ<@_�޲z��	�0'BD
���0A6�
*rh�(���`M���
�������r�l����M���=b%	Z�M^!x�ڞ�vZ�y�
<�s|���p�<�N]҆��a�0�"-dǲ�NIJ尔U���?h��?Te�N=fN��A���N]Q��zgvt��ա��E�y5��dI]������L�L�:G.޷�{�Y؊&Y|���ߋ�}Z�,�p+^z@���`QG�&�\����#���Q�q1hUH��I�QX>�C���g��jg��nb�WU���/ά �Sf�7�E�x��1�7��x)`���w�1 l�<a�]æӰd�uf�+�ʮl�Q�I��$�9
��u-f�[Y�2�ـ�R���#�~���ԒF*%G@WsY@di�s�����5U�a��>A��3]8�Nt�`�?���)��*��s�0�~K�@F,ys��j~�3��z��v��������h�ʦ��уurha	����Rb��+�[�����n�*����~ʍ!��͏�5\@�qZ�{�,��BL���u�$v-�%�_��,Ÿbd�k7��V�&�}If�`��.k��Zߐ�7 xI���	(^W��Y"�,�������/�^��5SU��ؕҫ�+�m��E�i�b	�ٽ*|��4����CKX�l���YQ�@T�_/-��.��ts�u���A0�f�:�n�B��3�oДJX$�gqeQ�!�Im\�K�h>�5�����J)����(&M�u�R�J�"���+�-z�t#��pn� ��"��7��E����|&��>C[b���B��	���a�dŶ�\S��9VDg�ak<CQB]�����79�p��
��ٽ��~�ǳ�<B~�[�|�o�7=I7�C)�z'�CrAټ	�`���zN҆�����L����ȯ��ܼa;>(�Y����g�zr.�����x���.[�i���[{@��0to�9�#d�(S�7�߷t��%�j��fa�Y���ˑ�+��& ���L��y6URx�I�S
�X�tS<'���	#u���"�-fnf�?��~��;{j<7����Ǔyi�U�x�(g�<�^)��>�����7�u��?F���x|"��a#L�vX��Ȗ�1�ʎ��:g�Pע��_4�`��!�z���Щf!��3;���T�h��}�i.f���}��l�_��K��UBw�M�r� ��k:W|�xq�U(/{�hM�Ũ�g4�l�ֱ	�V�}���O�LE��Q�3����������~�) 3hP�Kkt�N�ӈV�P�?�S��H&���S��(�/|�0V
��LZ���c Ѱb�����ebzb�CߢkL0�,���[j�V~W����w,��3G>{K�^(��r���E`~"1�.F�����o�x^�mT��ᄅ�%��Gz���WҾ�~��!/���"���w�c1fS븃s�B�`�nQ#�5�r����d1S�j�|V������%��<���ۢ 4b,g�"����>���Lj�bzØ� -���=JP��^5��[	��iƶo�VA0�'*��!H!�dh��cUf�Y����ޏc��<�S(�ټ����ۭ��Z��`�я��l�t��N�)����KB�� �`�\��c��qX�9�
եI��A~0��DW>�ߡ��b*��T�ALo('?N�Su�JvftD�\Ռ���Ykg��m���q����O�b�P�>�.n�)�A$�%�Ŀ;�����l'�G�|L�ο�y�p5�ˌ��-0��(���FyJ���V���j~��H	j&�в�r�-莙z��R������U�LE"�֤����P%y�G#&�~�9��5(1�p����	J�5LkXin5OGr"��i�D���q���ϗ<�K��$^���I?@�>ೠ�M��2_; z���� cU�����;���`��ҽ�h��1��'�f����i6����a�y=c���?�	��=�L�ҋ�L�w�,�}Z蒉�$܈��3�����@|f�S���cC5-6H'����X�d�ؾ�T
r�����h_H��ヷ@�./׃_Ͳ�����in�o��(�Hw���;�pka������X|R3~����I��n�U�cQ�ͭF��ta�IP�}�<V�~um�<�d������S�AC��x[�E/%g�'��4'�&#�,D��1�p$��)z�0��A�@(�K�3n����ʀ��7r�'%F�`�Ռ����o��O�5]Dy��jS/Kvs��4#�����Yjn���B�B`�L��Y��?�;�7^��Ì��$��Ӏ���?�%ܩ�YE�K6��4���+cǞ4�p��tLf}��jɳ'�,޻���5�4Fm��BT][`7��KqA�S�D��G�]� �)�$.�x1��ŏ�+c���;V����:29�;�M4�Z���@ �N����D
U6�gz�Bj��*��X��g�{�yy�U 
�{�ǜ�9�޿>��,���[b�zS)��Nalp�M�<���wE�8��q8B��>՜��Y�\��?jѹY�km��oыq���L�q�(m,d�T�LB�r�A7��r��T�vtD�!b.t�1��$/hg~k�-/�H�
.N~;x02�RD�@�T����M���9�o�o{�N�#%j�
>�>��Û+�/��.�s�z��l�R��	S��� ��"��ãPJ��$���E��<�T®�'n��[
��h�P� �Kc:���;��O�0�8!8�l3V]R����f��i�QPP�x�8b�����N��D_׫�	�@ �L��oR3<F)7�G��{I���RxtI	{BWm$�D<F�F<!�R�<4R��UB�&�i��������H�s�V[�����L��M^uMD­g=��_Q�J���\�[����������D��9t�8	\����%���i�1k�Xp�;���;oS0au��VB>��|�_N,(8@��~_�
ԅ\��'+�]���I �maŵ��_�so�}���|}+V7�`l�+�O]]/��%ύ#*���G?��Y�e.@��Q�&�^�t?*��9j��3�}��sIXR����3����D�C.]��j�莩*tFd+���!���]�q8i1����%�����%5�r�����;�9������.l�f���B�O�
a ���Pm
x	����Ā}X_�"�����{�o��M�l	O3�?��4��|���6��V٬~zݲA���v`���_��Ίv��fі�Ŝ;\|��n����JVc�6Y��z<3AԠY@���f���T�k�cyϴK L�}sIۉ�x��q���JV����#�ͽ��%j�B�Ҏ>,߽���Ws�`�MJ�3(1m��m�^A���"�R���*t{":������r�~����X���8O4g߰ɿ���Nt�n�<�gʜ%�9	I ��q㓬c�Z{(��[4H#
���>՛Ga�N�^��z�΂ �y�z��L�ަ%]`0�f'_��ӓ�w{����Q�'��uE?+��AiX�,_����|��j����YW���4ɲ)(8#�!�h�.��N"E��]����pEU��1���Ù�}���Hv�B}C)�̈́P�X�X��2��*R"O8EG�I�0���׉���u��@鎃��A�/=�-�qyF�6*�&1m}9�Ew.�6?��QfC~��F	�&��P����.��`�� �g��Gk���E
�Ġ�I�/��J
/!�
//�W�k���n�X>w�Pj����J3�c�/F9E��B�%�|%T�3^���+�t����r��>�ƾ2�!n./ɣ�P��s6��oT�j�Բd2k`�:_Ǵr�Fc)����L7Y+���̊ߗ�`#a��C���ƑnRn�,��3���W����Ƀ���F�J~���*�\
LCo�y�����,�f��Ѫ�/{J��7�V�0	��)-r#���ˌ��F�-Ys�.�MR^�1�os���]�]N3����e䆠Y%��re��Uݲ�R�=�׵Qo�A�<�(08������d��i]�m�yՅ���m`��������-��i�(#��P�nQ���yR�<����.��M0��P>m��6��[8PT��A+��	��m���x���hD��`�������8X�rm��#/�e<�y�p� g)�gk���z(d8[N�e�AJa����T�����1p����N1���f_��3�A���y�I��@����^��'<=�N`,�t�Kb��ɼ��{�&�^C����0]`�ƁZ�"sL�(��o�t}�P2}�ʪN�IW����*�ɯ��<�<�8PC����0�&�ю;��=aNT��$�a���Xc��E�j�(��/ʄ�m� ?X��6 ���+e���,���-E�);��*vhfre�#���1��R��n���]}$~e�㚎�����u���"%ԡ-�1.��Y�� ^%8��yy�͊�ĉ` � ��.���
wS��A4����i�1^
�&����Ew;��E���KO6���rR�.=��L��a�4SXo�t���p���T�M%�/H<����$��B��y�ݕ��Y.oB�� ���PlÇT
ۀ%I�z���cǸ"����!������v��fS%W��&��̝w�1���������Z� A'g+�^PTx�"+S�݋?i��6��=��A'Qo�����ٶ�G��ϙ��0"��^Wi�� Eq�3W����Ϟio�p���M}z��sC��pp3Sb�O/A�ԃ5'x�< �����u)]ZK[Z��V:I	�5�����G�f�t~��$u��!���8�"�`gD	1#ĦI�'��p}�2����AZ�����5ތ>�/�$�+	���#9����0i���ymubƱ8u��k��p<�46ӭ
7�}g����� ��G������[f/�v���L�Tᅷ~��&��sT�ӝ�d�<�$���ѫ{sW�%$�.�+x�g���_���d�iV�U������Ȣئ	j줞y�t�p6�����u@<�]-�D��5�.��k�ô��a��l�_;u�r��4%#@M�9ˎ	�E,�6��]���4�^�SM�Q�[J��؝*8�T��M1T�c`L�Y��˽J�y$a��Ww�f!o��{Ƅ�,*4q�ZT� �2r'�UCz��8���#t�=���d=���k�~JEz��KE��1iБ�5�ips��&P�h1Eb�M=�:����8G�~�5tH^������r�cU�m�e�7× ���������3�U)C|����Z~���K��E86�(i��l������^P�=�yݰ7]A���>�O��g{2J��t��`¯���8���	�0�ώ���uE�M�0�]�x�댙��r�n�A.���,����Kd8�E�% 8'}��W(������8ܶ�$ćbEi�Ɣצ�{�l�!��b��4�w&�]��� ���e�1��ty��#�IJ���m�Wxi�������u0Ы�N�fa }�*��ɠ���>%�Uj� `��&Y�Nj�������"���z�c�5fG�Oa�A���O�.��ە��_������(HC�S?�sgyr~�^#���j�'��&0����]�>֐���� E'��L�ɷT�B�u�k>4�f�Sxb�$��2�
0����v~���If搣��O����͎wk�	j�[�c5��r
��;X�}-O����)\�0 �ᘨ�[te0B��zWM�2�)vT�j�_��/�߈`�(��0K�D२'�ґ}��pfFچ֖�	�9z����U@��i6fWI�	��Y� ��C
���8k������a�Ɵ��r�u�� �u�R���P�q��5��#C����ZGh���YwKWP�U�o&c��a�7�k����p5�l\�Ho��^j�-��Q"ht�ir��+yn����G81��u%����[�	I�������cGX³�>I��_M���|�Yn�_�����t������o�Sb�"�??��k�� :{�IR�C����g 2�/s�V����{�򿳰@�k"I�h7��}�D�d��ji\���+w���??�*��c�0�ݿ����+;�9���3E9ZDE��FD �х������z~�15:�Wc��M�;����w\3��T�`Hv��J��l�j�8��E��N��!�2�AVW�r��;�����<�Q��lQXІ�5Mv���W0:��sw�1�a�b��I����0�x��?O���L��,Њ��$;�e��N\7�ls���\�����|5s��ܑ`�SW�צ(�Y8���R&�;��L\�+�!��[@��G�����H�c��.:X�;	z����"�O�	tT�E.��/\�����)Uhr�n��D5�����e����Aw��t{���>��� ��=+�ľ�@�j0���d]�����X����!j�(�Q�D��>��[��-Mn�H�E��5X�2����@	��	|�߂�"���#��M��G٥��BD���kv] �k:3j��tW�[?J5ی�q�n��M���6�O���K��%���<"��ꗺd�ۛ����))���i)!pf6`�U�[���R*f��0��̆7�a%�,$��$���J�[l'%n�%_��3A��G�����_y@�g�c�VE� �U���}-�:�(�c��0���5<gֱ��I⥷��E/cI9C��E̎��9P.OZ�b�`t����ܰ;ҷ��Z�^����#�pk��\N���
�+��)CQ7��}�Aer����Q5�۠§���0f�2�`�)M��4��@����|j��B���e�`S?�O��*����S�hB����������Krd�=˷��t�u&T��jOBh~�Ni�{C|�g��g�Wn�!�?5DZv��4 yT���MK3C�Ě���Q�7y����d��2��Ja�n!P3pM���z_��^�gޣ-S���Įb%t�i��|�6ռ�;#;�����w���̒g9�Q�5n4�n7 ���:�k���:]ރ^�R�!z��b��G;\{���O�%��ٳ�y~��"��-Z�(��T�~����ݐfiv�2�r���d'��ziy�&߂���P��wj���Ӷ�gdC6]�������IW�W�
5\N��*q��Q��g���.�Em�O��_NJ�m��k��dp���n
�Ǎ�8��c)�aH�E�Y�` ^�s��GO�>�~���p{��rS�)?onE�9��'���Z��(�o<ƩX��&~>~������h�,M2���w��HJqS���Ry�=U��b�������Ǡi���n��v<��vK�.�N}ߛ��̈��Q<���|Ș
��q*�������F���-8S�(B�90X��������b�j�_*��>��Q��ʹ-d����,��u-ő���>�3~��Ѧ���[�`�[�����&f��O聀m"*@�WT*�-oα���4�_��<���M�MJ����yz�T���u��#�3�>�1e=L��r�=g���i0\���~?k�P+�2Nòq&�}����P'���.�*�+|�@��,�O���ן�L�!j0���R�7U��y$��3��}�ҽnw���*� �*+~NB�9�cc��0c�+��RF��|�W��׮4�:zd��xl�a�w�
ˈ%=���OMd�
�_�U�<a${S�
h���ԮQR�-0m��Qڂ	���&;{$^9��O��4���ʷ�`��a�5C��؞�H�*���o$��I�w��7��5n�b[4,k^3x��a_��D�VԵ�.��(\�b����|6L��Z��J�lЗ{��)7Z�����	#P��}[�dlRD��9�FIH�������������������[�֟"Y�U}N�X��S�R6�p�XZa���X��e�|u�='�Ƭ'O�L�W���m�W%�Z��@(��i��@+Lː�S���H�E��CB�5�J#�&�6Gńǹ�靴��=nW��)�#�o�gt�����&�e&GA��%�&V
���#�
�֣�m��M���
908��Xr���F������)C��P�T�R�F�}������%%.c�<�������5���3��J��E�����j.�ﾾ�$����fg�����t��I��*��ps3u2��E�w�p���{�5蜊$X����v3���|�~/Xѐ�����J�0�	�^�~��z�	N�>b(}o��.Fh3�����a���OX�S�'�$���-�{dm�t^���B��@�N�����?ӻ�$	�@��6����Ӧ~~�u��Ҍ.k�!Ad��<妭!��	J��#��TJ4��t��u�[K�Lه��cc*�����~g�M-�G�+Oq�Z7�����_Ϭ�4�uKr�1���p|�Ii��7c|�(`��U��&���n�6��ӛ�� �E����Y_lk����=��Z��� T�S�P�����&-�����T�$rccn��� W~`�՚ƥ���lr���^��n9�΃�*����%{�X(u���~W�p>��U��=�x���y>��V�{�����T��.��QP/id����|9��� ��ӎ��J� 7=m�\�t�"~K��q�!�g�!��lg��SW�`'Xs�?��)��o�i�3�&^0vI�b�t�ܧS�}N�!|_�,�f+=-8��K��R�=k	A���as�KtO떈��Tz�2������z��0ݘ^"#q+�g8'�i��	ďCP�M)fȈ NG[���"��ja��8�9}�lh���gx8Z�F <���	G���cڋ������<r��w�B��r5M@���t�p�d��|ϬX-3a�p����NA�,��X��H
�*��p�x�<��+d�Y7��%�.�Q�!x�^RA<�����RRhp���^8�7�ݥx�_�-�g��+�`�S2�v`>q�,豅�U��M�^�} %�:�+`�nل �^0��  �9��r����� I�{v5��Q�ؓ����`X�rܱ�K����Z�|�'��U�tH��8�t���z�����q�,6b�Q���ߜ��)��=G?���AaZ���e�)	�R!�h;�hN�YHZ(4=��ދ���B�FL\��x-)뇡�G\�Bt|ț$R?fcb�! R�P��4ʧ�z��L��f���p<�9@��|t8q�xcn�Z��>���(1�+MC+�0OEF��r�Z��XU����fs�ޗ��0�i��d��o�#ܭC�ٚ3g�wF��N�\�w��}�� �ln�����uGfo?�$�����Ôi��ZrW�f;�|;Zea�PE�zՎ�e�&	�5�GoŘ2����ӥ���-a�'�~�\�@��i��׬� ?e�Ն������o��P$lۚ(�ƃ�Ͷ�זċ��c|��oZ�.p�6�%����^�d9���?{5��d��R�ZO�~���\�H!2����5Zݑ�WR�W2n:�B�F�o[,P#�O}b�y`��_�U|o���"X.Z�Z ǟ��#>�]ܘ�8M���R�e%�]�c�&�a})��N+^�֜����m� ��D��
�b	��!����հ��Z�d�
�;~�$X�����'jM�/Ǿ�:� Jը+0�b��ڄ�QSƿH35����𠞉9�p�*�$�9
�*!���Du	�፽��lB>�ꛯˇ@�|*.�� ���
����E�j.P�$���x5��c�� �T����Ŭ�30�B�'5B�	>5_�妨�UA��&�YK����/6<$���X����tb���x�|>T>yw�BQ�Icj7X7���X���W��H����U	�/R��k�تix��Xhѐ��$�����y:��^�G�K�I����L�LȔ�M��94�Bo���9m|8�:��nS�� \,b|�~G=�[�M�i�z� &���s4�f�M�y!p�F�T�w� �]kЮ�:�رi�k7�<CΚ��3�����~p`(2��!�ڲ�V�������_��L|�z�0Ǚ�e�HU��ƈd%�1�p���Q�2B�g�hA&�2�B���˿5�$�T�5��a��=��`Ȇ�h�h����J ~�g��e����=�Ē�������L���p�?8�L����VR�i�)|x#ihScR������Xc��e���E��+RʟOTR�7!j��4]�k�ɧeEj�xn��oy�^�]^��V$}�]lG�x�,�̇f��?4im�8O~]����D��W�H��?����o×3U�X��8�I� 5��-C�Io��5ށ�I�(vQ@���V���`$�H,(k�s�������Pܦ���]y�<�^j��W���˧I�7F~_��V�fw��o������.���e��ɱϷ*��D6���e4],���I�۔�������<mQ�F�q�Nk��L�P�D�D:�R�O=��U�T^� �{JK|}=�J��.��$�~i� �%�Z8��lO�dN,o��]i�I���;�������y%��m9���J�7�!���p�7E��^����� �5=awz��l�hN��܃�mhF%c�+���b���6�ޢO&���c*��'�������|?�H+=4,���5���2	M���G���8J�%�J\!M�Z�ȉ�������.U���,����>���m�m0�|c+�P���BT\��W<�ӝ#d+ֽ0��*v
i�(e��G�����/&N�úP��9���V��Ɯ����o�`��Ŭd��O@�*���,kJ�炽[1(*�fzo��Q��$�)�g�� �N��/�RC�w{��tP�?z\H�W?|O�6���`�z�qWK����9�9���:�5�Mn�G�BcC���p��q~��p~��i4�~}���\�i=����һ���P-D��3�� 5�����K����������c 	b�ے�����P�-�����6:�[�⌙&���$BA\x'� ?H?am��aƂ�Tސ�Y&K��w�Rѻ<���A� ����h��O��@hⳢ�SKӒ�G:c�_s���\��:��/%KSi��/w3�<3�wVF��3V�����az0	�HQ>�mK�!��`�F�EkC�.��p��d����N^����NC&�J^kS� �u�v �s;�H��*�0_�pl-،�{7S�?�9�k�bl\�1���=M�?�$pa�N��E*��%
<Ǵ��m�N����$LԳ�	B�O���,�Dy�3���cc���c�yY��<G��n��Ap�N��G���s��}	�������+cX�\^���ǜ��+��W��{J���g��O���q�1�H4X~-���u;Ħr���>"���C}x��.+&z�LyY����v� #"���3� ��+���5g�b�q��=��\�i)�r��	�v^R�8�_�!���
���1�x�����'�T�WTœ��9�E�W#ō��1�R[#����NoU��{�>�i�D��ᄅT;��
$\�NF�]h̹��*#صBu����!��4aj��~	c��(���lY�7���Vp�8*�<��(���l��Z����n$�R {�4H�xcn�f^v������P˜>Y�1����Vd���U�>��?A���;�4��/��ӭB�l/����{4�,k�m�.�m̳KJ���>Dʭ7�2zs
���/�n4)?��?Yї �i~ȇ?!w��TB�zG�6:�WuMb4	q}iN�?5h�{*:ĢX~��	��it��pQ*����,qfB?XE��2V���T����P8���Æ�C���H�G�W�4��[�����SE?���Cx�Wt<Ϣ̅p=dý ǭ��q�`&�%�ʢ��G�0�jY�΂�M��upς�<p�|��d ��h�f��	���ݭ0�
lG)s��V~���$n	�����%j���y�B�o�H��@\c\΅�9Uzj��I�GS���e]ĐB��\�K N��O�`�����HX�n�>�P��c\G��?������fE\���	;���±*�(Mlx�{*�`fN��p/�SV$	Ɓ/�B q|6Q��c"iu�h}�J:;���%^�c���[W| Z!D�o#�c� 3��t)�����<�\<����jj
f�ٺu�5U�(^���;�����:���'�]N�d�L�3TĜ(C�h��6����$��@�\�,��ݍ����"�Df'(�r���.M}`�D&ނϓL���<q��f��EW\�?��CV(~48Q[�����j��O��g�s6*�>���^ĵ�7��_�^>$0@���Ϝ����v�Rv�gxs�:Y*?�9]S�'��}3[��i9�v�@o\X��K��Ϋ#�f�e\q�'�A�f߈��a�)v�9@e�[G�I�/i[��x�	C��g[���f�6�`k�e�J}[ї����e�OL�=��xN�_�NFI\�-V�SR����쎅L��e< �g3��*�����	$��B����P����&q2����q�x͟Z��e}�)R��Ȼ/��la�+��/������; �)@
�׭>h;HJ�)շ�1P�qX���I	
O-"3����	�����7w�O6�C:1�����������G�a�rR�0����)Z�� ]l�H�6g�avb�W�����_0�QNG5����8�P/�Y�0�$ܳ�M��1E�����)��]K	ɤb���{4^Թq��7u�)#?y���L���:�LN���n��ձ@�~�$pp���'��%�&"�-����!vh}8�'���9+��+K$�B^V�8���aB	��N�F@P�@���Ie���6͔0��i���Y�<����.�S�0�c�fߩ�_�"P��gB�B�P�
*ttQ�\�af5X�uE�����g�4O5������6�f��'�Þ�lHy7O�ĝ;�z�MUf���I6�*Z
����+��y|��d��`�S�dS8_�L�w�V�X��ڙ.�h�]X����dLu �^,"KJH���ڨe��W��/�P�[/���+�7�J���\��[,;dxE�&z��EP�g���߈}I�sk�;֎S�
���>�*6B�13�C>e۷YP�x�Ÿ�#W�šLÕ����p��ƚ�� �L"=�:�]\��t5"��&{��=�t�����?M�!y��S��������E��ql��ߎv��'@���i� �;'���g��H����|_|���4F��5Y�a�I�Y��JP��y4�t�}_�gΖ�'���	�N-aR/W�r����K���SR����������s�^����W�
����d��;mfy�6"��#�6�Z�an��k��T�kKVv����#������*Z��Ѐ�X��e��@��Yg#�����?�=5�D��75��뿄��Jj�\�,ݥ~�JA�	��|"g$V\RnI��%���J풍EW��,�P
/�Yz^�>UX�_�Q<nþ�p8��z�&x[�M-��\�/x;ǯ�Y;��
�BnU̕�S-���.D�������?稵��Y�*<1���v8�W��t�M�#_]Kc
9�-�Y�������Y�B�u{m��S���m~�g�@��_d�?Fpw�K���� �w��@ʫ�}�3Ҧ)��K��!�3��
�=O�Ol�w0�":�8�u .�BٵwP���w�͈Ho���8��uxBi�iٚ�ݍB�X[�Y�W��_
<�r���ߡ�����݃��!�.�賹}�& 	L<��q�pײE�J8�h��19�>> ���W�{Ɉ�>i�{WL�ƌ�����+�;JvW#�J�>{�w�dCi����A�!���+ƻ���c���5�o���u�1��+�E}�	 �ޥh$���ޑ��@�e/;� n�[����Vl��� {�c�����j��m�zS�IS�m��\l&�-�m���IH����.�JrlɌ]�_4��,PU�\�'�֬�k[gY/������ˠ��h�
u�9��5`��l���0&�򼏯��(T�fϳ*����NX>�O�l���2}�7�ѝ"NTR��9�]��{lk*�.�c��=A5������y�����\�+�HRϸH��b/�U��a�A.��X���%�c�q�i�|����ŭ��E�I�����}�n�$G���zp\�gBo��)
��#'I�ub�H�C���$�[���l���m7_8�p�� =�w�|�����[��T+z` �`g� �����┵��TSC
c�������H
�:�P��ѡ�D"t���iQ���R{B)O)�\3c?��t�*�!�X�8E���A��n����2�9���ڼ���>X����'����E�����2��٘�i�Pת�8�\)���ܫ������=��v��A��c�����/+�v!��ϙ��f����N�������0��;x�U�,��/#ɘ��Ũ�dM7�O[�M2����n�{�4�bևH�g�K�ɍ�7`�ܚ�5�1!�$�|�#!7y^
8�1c����������l_L
!��$�h �'[��0��1WL�.�V�E3�L����;3.6	����ÍF�ff�G�\9{g���v���x��>_����L����c���A�˪|�����-��0�TSU!s���f'U'rp����}w�D:�?���i"�_`�z#$.��d��m��)
�[E��׀[Ѧ*@ᤤڳ��%���|�¨�ĝ���s@�Q����F���&� ����'�[�N�;�	������vT��Lvj)c\��5���#IE���%���h�m�P�������"�'u6����(z��4�w�uO�^�H���(CNn=�4�n�2�m�F!rp���$a��l;�(mș���iS>�y��˘oZ��]��x��l-0��ꚤOd�+ ��|������1��4=�anC�?�Y>jlA�+&�m�Ǯ)Dd�i�)�,ǵ��\�G�X�p��$�'3����\�\p��$����g7�RA��g7��Ʊ�Ҿ;���9��{����8G�1t��]�
5�f���%"pgP'�U�R}��s�^�p�'R���VT��"�2b�}/K��9@t��i�ĭ<X5�*1�6�r�0t�X���^.j`����RHfӁ�"'3�;��8���5+�{�+�9IN����¼��R1  %���������*���(��81�P�Sft��z,�-�*���%�q���2Q���!�]�
2����H��]�u�U(w�-��a-���iXp��b	���Y�fl4�v_OBm.�ko3� �@y[Z-#�I�*�Lf�].өw�����<�Sd�~�PYcdX|�i��3^���댁Ly�����@��1q�;4�k�jAG�{�Ʈ�=������L�@j�R	��$sU� }����-}�1ks�VP��o�SW�#u���7D�w+�+�Y��rŬ��^�Qy�U�P�d�N�\8�x ��ɢ�����I���P�.�8�z|����6��5����7��;�+���0�S��)�Вy��ߚ�c�f85�$��QG,�|�0����߽�j���0�M����V%4���h-����~�s�K x�����X��<3�Wzg���ؒI���s���� �ח���6�����#35�6��:fvg���U;w����]����������N=m��0�%!Vގd�W�Ro�C�d�^��!�8ijW>���8tv
e 5�?"���"�t��h,�x
��7��Ƽ�-���5��>j�����`-���������֝�;˧�:j�HS�T��G���7�'��P�!�~D`��v5�+�����p~ ��#��nj`_�_�d���x���ޛ���Է7�>����=��v +�gZ��"
桨z=�gc���3��@Ct
{�����	N��Ws��y��b;ڏ�&�7�C0�����l��U��<&lJ�j�K�J���(EAa���#ݝQs�a��anٍYa��1=sR�ډ�^Yk����t���a"D�2�`�n��q{�r�\������Y�P�Y�_4�fS�l1�H�M;�8�<��|��~t�U�:����B:�)|�`;���]Ĝq��Ģ�v!%�گ�!hX�¦��V�G�6��ӫ�]	�{�M�?�5�}*�~}2����c�����D��7�Mߠ��v �%�����܈>���k�,G�������ZG���L���	6< �&ҥ�$�l�w�cok��W}��F$ac��&������[����b�'��v7����gn/BVg�u�d�)qE��P0��1�T��m�����{�g�DV^��|�W�|"7,�~r9Sp�uJ���	1��~��'��R@h'��՜� �T���
d��i��؅��|C�*�Y�3Ǵ��?�����#�R�y�̈́qtẒ(�z��H�4�V3S���No�N���年��N;[�ȧ�>%�᦮|��m�ڸ/!
w���Jr�L\s�>��jqp��w��V��f�W�E�<�2��5�qn�¾S8w�����B� ��HZͽ=�j�yn(VaCI�:���dO��M�D{c�|�R�?r9>]�-�:V
C�*l?_�}��^ώ�.�y��z [ P�3�0D����>JF��k��%u�eF@x<�qO�7#���XVRW27��R?O��ly�rJ��`]�T��*����VY�M������5�d�!�f�������>z�³�tTc�SI���c�݅�W��y�C�!���*��pK�m�o�G]�%k�����>���G��;*�N��O�^b_�m� ���I὏���w���%p���z��g���gǃ��!�p#Z�9��g�q1��2w;�jr;N�R�}@���I9��`!���w�[կ��{�R-��� �5��[,�2���ǲ��gU��C���X1���˂�%�o����T5�]8YJr�(P�����1J��
�E����3~n��0'B���EE?����}�� 輇υ`���s2$��~�F���	E�z>�����`\��6G���-A(UJ�Kӎ�s��@r[0 c������`$s9$ֹ��\j�K�S_v\��I`�Y����'�>>C;����=�8�Re�0�#�h�_�V���7��T;��h��o� ��*�G~T�����if�.�k]L�k���u�v�	��@�yz�O�����ɽ�)�����X�q�Rzf'��9j�;ܟ#�To�j���@�#zܣ��qq/0�-ǟ&�f<��_#gT��S�$����%Y�$�U���f�zm>�&�SF�+O��,���TG��X�Ɓ1F��x�@B������h0�z[��2��㜍3��,�B�k�-���d�E�g�&u��;k �݆�^kN9?Tn�:Rwx�Wb�8���΢,�U_��~����!<i&��bvj؆����)�����z�ۺ��
��"�����7�).�:��˪����-�6��b��"]�%�G�i�g�'��&a�A����a�J�xQ�T!�zs��Y���sJ�T��l��Zs�9&FJW�q�݂�D_xQ� FL�}�aؖI#�UPCm��ݝ.�90&1i���O�B-ŕ>�1��.R��@�0�g�R�t�s���.`|��t-� �`J)�:Q���\f��~�5]�����'������q��%�BC	E%VG�aϊ��%�|�������;�