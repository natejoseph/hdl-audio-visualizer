��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CG�ʜ�S_V��HrG"���v-k<�	��	0�������'g��}�,�_�E�n�����1�w�C�>n�� цa�N�j� "�=��0��B�ȩ�_��_�Qנs{�E�
�R�%�E��T��/ ފ���<������C(Ks6yZ�K_��ࣤr�'7~
���\%l4G�Ȅ��a¸���I))�.�;�qFل�P���s]��w� q����Y��W�h��w�X�T.��ڛ��	h·�*��d(gJ]���68���<�3��)ī�oڍ�<�ă.�����6	��Vث�MdS��7]z��Ă�&��Ԯ9ҕ���za�(کߋ�$U�)V��^�*��_����(^��7�[��^��`�U��ٙ~��p��l�ݹ���F��ͩx�Bm��y���bL���5��֗��24+�r?�7Y��a�9|b�C��#t� <���?����Y$��BA������KJ^�/�&�OH�c߰��h��x� $�Ɯ���Kx0'�ܤ�C�u��vc!0[�ɏ�h��쩝����C�\_%7Ou���Ŀjۈ���ۚ�؛�nu' D34I	'�lurO�6�$鐿.���0�eۃtR�`�=\H�?Y:��!&����S�dlC_�>�[��칼d�}����@���$�x��d�z X�q�����#��)bNݳ-���3]�yؕ;�*�^k�$_8/�+v�"�m%�.V�X��J۵�V�q-k~�4c�>ɢ@&D��x�Au�?��������My���gǟa��x!�+N�y�CSҫW
gƵ=��']��W�����DU>12�΃5I�w,���<̆�O���t�j�*�˹�0
�Ѵ(�U�	�
���{ב�b���tq���N�<O�q!bZ8{-��S�~���������c�ɥ�wT�^����7J��j��
h��hʵ0�M(��AJ�i`���;8�C�I��7ٺKr��/b�c8J��m&s�2iCM�?�zz �fԚ�/%r:ѷK��R��Ta�j����	vHU�Yk�dh�.Bݖ�w'�2�tI� /t��>����qñO�@���Am��L�ӉnN�]�<���ʁh����6�+i�+�
W|ϡ��Q��d�CfxX~�E��}+�c% |^*��磒�3��˜�17)m�~¢�A�$�b����8l.)����4��v�X]h��L;\��������O��d@��j����Bo�7�#��Ϟ�᛻ ����[�W;xr'w<Np�3��"Q��]�K��;>��n������4�=��$T�#03g��gR6��5���k?�d}�^'NI	*�n�������T)kVƿ�.�mW>Xi]��8����3�\!��'E;�����y�xТ���x��鲇q��Ԋ&�rl���.ؔ`H��������Wd%��SP�KV���[o�P@ +�i��Ӑ\�ޜ�Ȼ��lZ�� �k�5���d��V��
q����(=7������j<tk%=�7�B�z�0��*i�uO��uu�9��̅��0)M�Z V˦��x��wRm�Ay���r$�ǯ?ce��� �M�z1 ��W+ۋ� � em��SM%���PՕ��W��[(8s��/�\�A;٣�.��85������nSG@�!1�҄+WJ�Kx����7�Kw)+��O���"�=�E�q
Is�W��)�C'�'���񻟐���99��[L��z�n5\P}�e�=ڗ��)mj�i��Lj6�O��zr�$���4��x�XQ2T�C*���u<N����!�<�.N�ȍ��L�<Ǖ��QTZU"����ȗ�Gr�)�2
�l�o$��{}]C�6�	^����M�ѓ����R�7���A��o����9p��@S%/�c�<n c�{(�K��!f^-�oW ���ЋYaIn�Z���@0�8�*�f�sKzvWUNtĄ����ӗ@��x��,�B �	�7�#_�%R:� �����'x�}\��cu����S�g�.�&����n�h�Y�V��t��:��+�.�'i[�F�Tʯ� ��-ʇH�p1%�R`2x^�e�+�3�X���	���ǝI��)@��F�=��Q,��~�a57�<n��)v!�0�> |��75�aw�^�Ym`O���栧Ȭ�-\�D\��:jt�<���j
!��3J�.�3��o2��UV�P �){^4F���{j��
+ټ��y2Z��G�"�X�YRxu|U�P�e��
�J����a���%	�cs{X���|�öw�u���ue隒a��q�kb��.���/64[�C+עƠUF��_�P�;���䮺�_0J�2��[�FyQ��צS�g�lF'Y� '�ifF�~�h6��ʑt>�yF{�!C��9���o��4(�~�Q�:v�ay�ɷ����J���	���"�8Q�^=��=P�Z��\�b�"�"����Y��=�|���.{�d�X\��o�א\�B��?W0�Q��.�ѕ���;���@C��i���sfT��<�=`ڕK��o2������?;�0�Aڭ�� u�Ns$�b��s����F��{���9��B�"����2T<��<�/�zD�na|U졔UUz$*B�sp�,\*6v*���?�+�^�4D^P����`+[%�	?�j5��5gZnZl�Ag&���8���mI��î�h@���h�Ơ`
m�������h��h�Ì]��}��M��e���� �=��w�������
K0˜�A���+i�x�L;�1�M=�p�`L�<)����&&�D~��V��F:e������xK����E��񷴺|1<�!�m����R sK�6�ziHx����ج,̎[Fc[%��[C��x�(ûß��Ry7^{��d^����i�6B7���~-�{A+:�j���.�b��\{b`�p9%�Ȃc�%.��s��;�q�S�HO�&Y�Bm��0a!e?��F�Z �P��V���3�֚�M����H{KD{�Hx�,M�	��ݩ�m�k�ς�&��w]p�'���^�a�S�4���s�7vZTX��ɷ�����+�������-Q�7�3odc�d�#�r�#(���jkw� a��=���*S�.�NO�'���Wv�	�ۿq{��d�|xW�՟��9�(��ukh֬�j�c#�L�c���D7wQ�L65��_��Sj]+�e�SY�#�\�8�p����Wc����J���l����yK�/�J�a�?�g�ܓV�/GŠ��	��J��ڳ�<Q��ض�S���1����;,�E6����� ���^��r���i1u����V�&�z�.��G�]2u����hI&	4�B��a���;�`Ӣ�4��N��>���ד��>��[T�����L6~�����T!�4~PI88����bW�m���k�疗��
��\�h�"'!IG^�i?�'r�z��Bf��ar?����9pP5����c��E���p��x�G��vJ�����e��!C�`!/�����ΟJ���~\�����,L��\�^h�#V�i$ҪB��-A:�Z�I�4���D(>y�(�6�N��S/dAs�=��[|���Q��"<YJ�O���cg'�Ƈ�꽕+8�	O<�=t�r$�\��쓝�e7�����-HM�H�l�
m�a����1�1=۪�C�F�e�����5�;b�@�)��>{��V(~���1h`�E`�|� !9|"$c�U����N��M��}1��R�W?����ȢW�~e�h=��vo��q�ε��7\d�gٍ7���r��'߶�g��ɞ�K
Oz�yv�uJ�r٩=wO����k�/J���j���ӕ���S��O��a���14��eLa�KV����8C=�9A~ݣ�+�o����<�&���t�Llo��i۰�'���l��P�w.�g{ǈ�k��M���_j��3��[��i�	��
��-e�G���k�#�ޥ� ��)�#�yы/������za�&bc3��֎K�W��E�yw���{P�5�qI��V�l?��9�^H��$<`�{��s����:�fM``��_k�K��}��:�.u�c�{<r��B�?�I���a�56l�>~CtU][�0�Kɗ{^�i+f�j�^�S�x"���{LW)�jVW/�$w)��Z�.Hn��G���Ku�[��B�B},*y؉ܻ[�-Z�٥�b:k�3�<����Di��h;v~�~o��;�kk6fFz�я��z԰x9P���R�%�Q���C�%�(%^2�tZ�h�fs�������aِ��m�&z m	û1����#g���m�q�l�&��Y��DָV��vc��ARc���r����̍T����1�CrԞ���h�a�i���y���n��d�/L1{ԇ�'�b~�}������C*�)ya���t�葪W�L�#F�_��h2܂`��`��nc���k��^��7�uV� �C��6�ܖ�z
�F-��&�蜃	[�#_��5yI)���Tͨ@è �%?~�cp�"L�8h���z;Ū#��y��OƉ ZV�l���$l�Qul�؜�j��~�x#���Q�����w���O�H�Tۧaa�����K��^�Z8yV�*��(|���*1� f��@��k��[UB�3s���┙�ow��U2�	4�|~�a��E���`%�	dD]a�"E��V��3�&����T�d�6i`�9�}�Rk!?|���.��uʋ�#z^�7��#ZMi�jHc��k#2�!~J~,�WM]�FQ&K�|wK����?�&�9���p���� <�{)Àm�I�i����?%<S�����o��jA�ʎb��:��qX� �Q��W��7�K���[g�IQЕdY�9��wD �t+��&�a�˸z?��ޏ�4�����jg��V��	�-o�Є,iw�2P�x]�t)���ڧ�����-�'�J�֝C�����zjb���4�����"�r�����jL��W�[0�\�JV���\Y�*&�3�E�Ǜ��[��w1� l�ұ<q�Ǿ� 9P�Tȗ��T��i��>΃6�g�1��$kJ�,��ot��D0�����J�!�%��RH�t���|�c?�ĎU�$+��\��rH��R�ևȲ�\�[#�ϖ���gV�T55��I�����!�Wx��I��Vb	��ns^��J"�|z˷�5��5/��_)�GK��7��]��0]�e�6�U��Iu�g
����	t�[hW}�����5�7��9R��;�^,��=+ ���$������#+^���3���H���_2�Ŋe^��If��+)I�8Z���ip�#�,��L5���� =n��e�2$d���z�,����\�r���,���(���=h'q�����U�>�����>Y_db�G����^j�Wx�#r0��A�\C����Q(L֩�����b���R��%�E��AL(��9g6�� '����b�-�j�ò��p
��(z����o6wW]�N>�K�0��~&J���دF�pƱ�κ����m�pɁ|R#8�B��)�jW�8�~z[� pЕ�Jgk��=N������=g��Y���x4K݌M7�@��q��2��P���29^�Y��^�S�����k^p�Ջ�ٔ?(�e���Ay�H���4˩��h�<�F�.L�u-aV+'B{���Y�X�؇4��J��@[�>�0�y1�\�XS����U�X�6MS�p#��@��o>����^s�3_�>il|�E��W�j�Y�e�� �7(�)�HK�R$h��s%�~ ��j���}a��y�oT��~f�NpB�&�H�-��la���ev~mSb��4߃�Q���0����#ߍR?�~."x������:N���2�ݹ�^�]����  y�gAb m�i��x�<5x3��&7���?�.��+u�#��8o'N��k � p����}���M=��-n�R�����R`^�[��&M<k6-����q�k���Q�(ڊُh1�W��@���)�l2��2"��\2� `izJ[ ��w��}�lC� �S���Z�$��$Vg��=3��Rb"���c�h�����0B����GNAs�v�b�z�&���Lh�p:�t/�>\ڇ�M���,muS��	��]��j+��a�@J�3���ek�X�@)���k���D7�w����E^x�>v�������L��΋�4�i���b_c��8iG�ڗ�&n_u`�D�0d(=*յ�Ӥʔ�5F ^2����i�2�R� ]�}����h �;�"9���c����~��]���9~<�'����3)��
'5D� >�b}rF�$Xm�u����j:��������hr�?��	�����z?yy~�EM�����N���9p���K��b���X�&g,�`�	�;`��K���c�/�@-6e������> ��r�`�8I�P�΂@�8�R�?�+��Q��N���e�#�v��NŊm�bB�	�ZP�TH�AU����{��0�Ց���og��!+arN?�1= �����]��h@卼��o�-Muw謧ZM�k�=�7}<$~�"
݄Ɇ㋚��M�&�T1;
h�����n��5]��&�l^|��;�4�>B��)4!D��L�0Y=��݊���<�#������T�.4�y�
���#ٝ���-0d��䘎|�5� ��OJ7+l�v`����������{]e� � :/����$'o�b��|̻��Z��Jץ̨�� ����=�ǉ�T���Z�F1���mdZpûN�����L���x@���2D�РT�I�Jx�g��F�6�z,�ډ�ۗ��^���1�k45vU�mVM�>�4�'�J�>u�����͑�U�s܋��F"�9/o��\[%�����)T+\���5Ba�K��8�Zc�	
Pu�Z��5������}
y˜�f�B�[v�nu�h?���鍗�9���Y�f,����֒�����o6�y����k��{�4H�B����>D���-�K���(D[��b�Cu��������-������>�/ s�O>w�e���t���ţ<I��͖�Ww!����Y�Mi;Z�~mH�Qcr�I�;�>߭=�� g��i�3�a�+�Ҙ�G���ʚ1��7��ŀ<ݼp��+YY���Y��'��6��E��w�*��A��[#�9�__=�g��ŗC����'��t��op|�Ȯ��Z>2?v
d�^Vi��z�6j���v�Maɻ�����\�Äfe;a��`�����k�( P�{���4���K�êDG|D�vT�B(� vs���O��Q�$�a�A�p�qT��E�F�6ͷgV N�>dU�E��5������#�4��O�:��B	E{N�j7lh�ј�"��Re[���}����3py�n�}2#��y	�W�]ݍOd�_��.6�E<���8����p�Ջ^/��N�~��s�U�̻�]P��P_G����W_�ѯ[z�5�\���z��s��#��������N�O��ϢHG5���Ѷ+L
�5L����|g��K�5�q:��Uż��@��XD���S��^O|ʠ%{v�}���=0^��ͭӳ�.��;�7��p`~�Z�ަQb�~��	\������{b`��)�:���G�|�������?��>q���A�Г�)SK)� ���ԩ�ǘv���`d3jL�Q�h�������>�����l,�FQ����#�{���op[+�f��9,��cg�G�`��;��F�~b�M[F��$Q�x��1[��`��Hn�a�G���$p<��v
�S�,�\�C��P)X��
�Q�4I~Y�ŀXL�)#�D�ܖ�p	`��<�crR���f�0f�δoQ
��5 �Z��2��f�*�!���+���4Y4�����_SV�e�ވM��c�'�%���a�����u��}�r�vt%M�W�bDCX��f �W�A���@�|6g�~�>f��Ϣ��=�:����[��Ί��c>�^��`���-�u�?־�jW�l7��K�Z:�&�)�h�������v�v�#B��ゖ��P