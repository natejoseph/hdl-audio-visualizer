��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g���`�SF�Z�6v����(E�ݻ��<���� �1��4Ee4>
*9�g�Y�� ��3�I���mw`��ڸc~;V�!<���F|�Q�o�;�1�Ϝ��'۰�8n^aU��q�� K�y��l��㱫ry�B��x�!v�h�;��&!%�x�b&����_��P�,����A_2�	\W墺&�+�Z�t&q�T����!��a4|_	']^"�d�ys�d��[�k����ڦfwG�Pւ�$��%tCc�� VSq��g�����c�� k��y>�D|�#/�L+E%�*x���������B��H̼ú���Q
HO[����z������`��K�O8˖���3�ش6��Y��6>_�e�U$�0Im�4������!NM����7ܥzyX�T��2ζ���Dz��ʃs��)�H����Nx�����=�r�zn���ƃ���|e�ߧ��Jg�ﳌ]5ŀ�٥�� W!��*�0{�&X�1�R�����p��|����߶[���.�x��3Q��y"EU��� �at(�]&;��;�y��\5A$ ���8i���N��|�����bz>l�-��+UX�
H��at���pe�+��E�)�����L�ˑ�ݢ� 2�	�������B�z�����XH/B\w��⥷�F�j*E���``8YX g,��v�R�W���G�yq_��2f�9�FM/�'� ʩ�Wlpn5����ZR�T�Ơ@�K��z뎫�s�CBНt^A^�0<-��$�(V�s�3�V���z;��1f�m3�&�E��a���Vw���}�E=�a�i xt�T��]�5��r$�!�����E50-ҩX��˽���Bb6���N�j4NF$�0�vϭ8n���oΓy�֥\��������)}I�e�Q�-������Ӆ���xC��g�#�����fn�?����[�-��k3��'�G�����-�i�%? ���H�7���r'  a����� ����D�:A�����k�Fx�Py���#W8�e�\�� ]V.���RZ<A��	��,(����� bW��&���>��U�<?��g��|`���
����y�	0'%������r�X,~�]#S:`������7�4.�E�8z :?�U��J��/�׉�]��C�\�o;�h6-`���vE�+H�1��{(|��N��1Zm�Z�l�0�U���y�����<��p!���zhv���?H\Ի��:�1�SM����D<�4k�W'��f�ic���k��L���G-u��fnn7��c�h�\.�JȂ!����[���^d���c�/��gYY6<ѣ��Qr�����L�C�+��vtn�$n��9���>�s���+��b_�0f��!��s��ʷ�#�t�o��=�݄���9�3�C
s���^�qi��)&3i�M���)U ��'�2���㗧�N�������K��'�_"�TtEΒ�5��^����E���I���M����5�0&5�D�Sj���V�S�"hi��;�lׁ&S<���X)�Cr�c��`��A;!^����ㄜ�с#�X�+a��{H����L�m���t��*}�hI7I5y�SI�D �������p�<X�J�CdW��ԯ��eT�.IiDԘ���_V�<�2�N,G1`ujyP�s��YH�̺`Px�ZC@T�!�7y���ṋ_ʵ��`�)r�5T�r����pmrK=(�S�G%�Z����#8���������RF�I�0,���'�ӝY'
����6�\t����	���a��:���8�����@gۗ�F�����%�o�[��]�pMf9{��O�jz��H�u�'i�,T}n�4Z�P�0���a�|P|fZ�����&�"�hS�*�%��ې�7�u��ӔM�C�����ЃבT�~��m���q�ˈ�g��0��2��!G���	U�ܝ�����:�c�=�����}MG�#�y:r:@��O5�!���^�&j�'���p�:0xڰ�KU[S(ID55q�6�G���^g�I��ۜ�m����G��zϡ���~bx�+����Q�A�h1��+��eS�1!�l�V�zgH�����9���ƫ�6J�eE��NG?̋��'I����NF���{um�������d�7-D��O��16� �P��X���Ό��o��c��C�$�R(�^� gf��&XqȯQz�,WͷOd�B�oo�� �ƜSh��m�|>���"���pv�6�����Ke���#���}�Bz���Sh8����8�)�n���ˤ��FS�=h��g$:�3�R�{D�ݕ\�1K0����X�~�]�:�E;�ȁ`w�o�y*����R�ދ4~�4�������P��۶oDMi�ۙO������"S����1Y$äoXk���UD>�\t�$+��<)������u��S�fO6�;��@`�o].E��(�S>������fLM���O��nHͣf�}�%��5��ό����nx�c�Q8��'S?\?MB!�5D��rQ���@�w����)�RL�w�Nn�jg��R׷��5��~f_�y�tb�c�A���g��3�<��I�}�մMV���H=��u�����P�rV@�Jh��Ő���F��
\��X+�GUzXIuڦ���@���L�r_v�,R�P2�K04O@�ϷLhj�=a�3�oW�u�����O��	2i����va���R��i�C�_�!�e�I:�vH+\���L�kK����tw'�]}���̮���0��J��L���A9���F�T���#	#F_Uj&G��"�(�[�̆�t�H](�h�h���G}w`�7���.�q���B�9���tm3lM��4:�lr	L9Z'xߡ��a�Z�N�h�D�����:,Ơ��1�v$o���'DX�4�@dJ�gq��j�YZ"�O�@U�S�!"���$�S��Ǳ�l�w>wf6s���(��.PsE>�jCUZ��M�^,��pڍ}�����<"H85���j��1L�3�K��<�(�2ŧ{�J�\�{�!�%G6٣��x�<ܛ�N?Կ"K��ʧ��Le`|�'Ǘ��S&N�W/Еe����l7j�+�����V.���p�!ɅB��$��������m���`�b�D4:)���B���=��V x����]	�����ߧ���SUC���e���@�6>����*d��l=^[R;b�� ț�c�O����'�5H#{s�S�`OU�HƇ��$�X�e�����bO�5��B0O�V�\d�4���@W���H��Um.(h"A����
�>���#�S�YP
4�݄�L�Y�a�p��x�C�M�9{'�|�U���ިo�
>�	E��a�I������{/�ӑhRΡ��@��Sۚ$�s���<݌���~�E�	E�C ��}V�Xz�	:����R|��c��$���b�X�3��Tn��	9�����D�&t|e{G��"��7S��)���3{)��bI���D�������2b�܉�$�mrA��5S��,�X[�$�/��=��ՙ��q��(�:հ	����xm;f���t�ȬW�CUUa���ˬ�L�-|D�u�H&�'�׵�;��G���F�O������i��$�����޶����"
M�����g��]1r9���\���7�	�D&g3���'w.�EK:��4Fէ1�<V�P��������1ToT�˸��bu��TA��6.���b�ٺr�Bm�sW�dOH~�$"Q*1wLh��WC{�PF������SQz�+пUkaj.q���ώb�޼{l��6l-\O��z]�c.�sE���e�"���4q�zǥ0m-�K�M��l|��w�%���Ŝ�Adv��|$�=Y7ht�U��8�=8b�|9�OM���&w㻽�g�J9k���[V���*.����;(�af�!��'��u,H�M),#�`zv����qN�o�']�p��"+s&�i���+%]c��N�Ǟ6�bP@�����<�%��J#�fH� kH�-�5�I,��i��i�iY�*�4;o28�B��|�+�������qw�"�v䆽��w�w�.�I/%y�Z���=+��r{��j�##�'�]�t^�������������M0I�C�H�jT=�6�<+CF2ѐJ�d�JFʮR��b��wO��%�*{Rig�i6���Q�c8�!�
�,�YX���Ẃ�	T��S(����P��,���T(�u����ܴ�DN�L$��&Dt�V)�5uȤ�r�a��""�,�G�Eg�a�g����I� _��?�t�=L�]w!�TĈ�Q)��W��I��/�\?)כ�x��Jծ�^�+�z�H=��iE'T��BQ�:�(Y/W�U�E:н,	�6�i���4ƞ :7,���i�Bפ���Gwl��k�U|e������Q�)��<2��N=�)�������`�/��KQ`딨��G����(��ו-QI��^Ui{���R&���_�bϪ�f��j]���e�p�^C�16����k�H�� g*R�1|[>f#b��)�#*������&л|:IV����B�$[Y����e�p	 mD�e��J١h
o�@S�o�V�2j�:�"lu�Hh���Z�e�!�te{���
�
���nz�w�,���X�2���?�v)L�Y?��?��'�s�W\E�o2�'��}j㮣�|��<�C����H��hB�9Y`�X"`�1�lr@ȲkY�0Ncnߍ���s;�a��#�
�6t56�HB�#Q��#�v���qJL���Zթ����HX�Ђ����6�a;O��#qw�8��3���0�r�m6tOӺ>E-��p��f��7q.�||~Iʚ+��u¤�A�0�c��1Nʷ��n��j�Z}�����9*�2��*�W�����$�~�+aH�N���q�A��x_,�X��H��euԀ�%G��T]$<iȿe���&R�Qg_KQ��{��	�]�yƮ7N���VtE��wQ�f��Yb��p�se?ߋ�;Iҋ�q�Z�9����mc�v��0Cl�z�A^ߘx�h�3!���&����X�&�DPS>�d0�g�^��c҇�{^v�k1�����_Ƀ?R�]u�
�ݾ^�� /F�� O	UIQ%݀�yy���g��
Fh���2��*��#���"��&A�,Az�#*�\u]|d_|�s-k;�i��5<,̍>.��j7���O�q��]05�@7D��d�Z?��]�����ɑ����dhĤ���ձ��v��oO��y[�M��y4��i�����i_`�#*�[t%!�ĵ������G����N���Ũ���[#]W�(e�|�>�c1 0m]�/!�W<�G�+��)C�/*H@���`�atߒ5f�l_x$��Q.�c�X��+GͺZ� ��Uo;����i[Y�Z��%�� ���X#{�h;�^㓰�Ԫc���	��t
_[�=���U�sV��,������Y]�Э�����x�b]f�G!�n/��<�#j�Ѷ�8lL�<EF���@|"��Clzpo���ϳ��e�D��v��㮓��~��Z�~r�8OR�"���Q�{p�mF9aO��	#�K�����T
�xU!zz���[\~��f�Hh~J���$�SF0U7�Y�߮��z�s�oZ�6���V,$|�0@#�E�"���")j���ں.Z�kVc3��wgH�X���	a�y���B2�<S#{^�K�ٰ���A����mOT;8�;�a.]���A��
�ֽ�1�)oBu�S͏A����������D�D`k�3���"HDΛ6��,�}�Z�+�t�~xzN�՚9>���1��B	�:��n:����B�����՚�Y��A��di�?��%�Vu�����w|�,�f���sD?�y�F��>=���=�Q
P�v�/�t^����⭾A��`
��gN8m*����\��_�u�8���2ѫ�&h�G�w�g+d�}yV��ĳ��,c�]3.�I3b�$���~����IA
!?��y�=d�ɝ�Bc2�P��,AB��gmWpY�@����B�'������B�h
�^�����
�pH��=�
�!�w�����,ޯ'}�r�P\U� 5 D�ٛ���֔z%c��ܔ4YYЎM�eS��݁��Ҕ�c���nV������vT�x��^Gh��>2Q��%��lӿ�6�12��-9�Z�������$��eogq�u�u�5��X�?J�zB$�U�?�𜹢�4�S�<7�[�"�߫�։.<�?"�\IG"w�Y��z:�H��w)���l�3?�`�Rڶ����5V��+Z �^C�m��!��h/K��,�(��������΀�ȁi^��<۳dD]D��)��$F
*�M'N#����� �x�F�Q���q�>��F[`�ޝa�_�kl�4�[6�)����T�G�N�M��;��~r' ��Vǁgf9f�3��	&9�|���#�"�;�\V���Ң������o���PX�@���U�u��a*W
p/��#���ʙE��������u"x�@��������Dn�+@�k���F�1�9 �DR{h~�Z�J�j�鵵��ﾭs�U���;tX�T�o	�]&��ēK�_=��]�+0���ɨ�EH��m �Q�t101�q%dήh�]�~�ב�q���n�Q
�V2���?/u����Ë�<|:��(J>��ES(�����<�U���,��'lsrR�9�ӌ)?�u���)GD{n�ܣ"P{n�$$-�785�$Dmי��>��6ὼ�nR��t��I%M�J��z��սX�V�a3-��'���Yo�-<ۥP~�w:���W��]2��
vAZe�]�/Ѷ��a�p�_��n$���4�-~U��>��'&b�d)���|�s��D��91�Ӗ�$�]�<,�j��m���#\>͑(�ұ�Aѽ �{�����Q���¦���:�&����>ƻ�$#ݚ�Sg���6K?� ���/+9J��*�]�2r͕���o�J=sf?�z-;ƖgF��`a��VY9��q��v�`���YR�t%waw7
o��)8y4�@Qׅ�h07U��Nf���OB� f�涔�`QD�i]�z�T}�X�ʉ�˖|`�,H",u�V��Z����e���r�"��01�!���[�CE[6�`�C+�v�g��7��X��b%�/��S{c����g��\E v��y��h�����~Cd���MO NN�԰f�%�Y[Qw��׶�.0����kL����0WpǏ�q˄uwӁc�����B�3'sz�[!�������ۈ�is^������@:Ne_D-Ǚj��k*g���2ʼ���@=��:s1�]T/ͦ�� S���vB���_)�@����u�u�l͕3�J�n�h~��0m�償�wp\^�/���V�,}ud5-��5aeZ5��ژ�"Rϝ����Aly_QW����m3���>���o�����P|���
(��#�(���<�҈�;�� 8Bd �|�M�B��<_N{)��ٲ�^�6G��#^9+��F��=�kN���1p�	ߣ�f�{���jΡL*vd���;�;��&u7<u�N����M"1�Hm_��+.�@_���cC��S%����N����2�
@���d���d$�1} �M��U����vߌ���fήyO;���Dg�Qú�-tu��}Mj�V���\�[���6�q�<i@�99㉾=��|G��`W��7;�`�t��/?�'�>2{���v�;"E"HXO���,�����,L��	����'�B�5��.Mq�3lH�*}���ͯ�%Nc_Y�ذ��e8���j�o���&VMq������\�ü��&|?�N,Ion�ۭ�<Yk�C��Я�:�\�6#�UĪ:?J,��?�h=D��|����L�^�<S�-��H��t�H��R*��-@m���*kV��}ҞYf����˳�۫s��Enޚ���l�G�e����ƺSz�i��d[�v�4"�`w���W���x��wP;d� _x.���9�A.2��D���3 c:���z��=^Lp�T�Q%��R��P�0��t�C���`+buo�����Ռ��e�6_�U��Flګ'e�;�팓� �S�j�GqP1#�'�+�Mdy��ŀM^2XN�U���6��ׂXD��C����O~�v�A�kӫ�j���L����6~�'*閕�~j+�s��+�g1B�� q:F����W���4J����Q۱�Mi��t1/4��a����؈��C��AMU�O�\����@q��>Y-D�'�X|as�dc�E�d�l�3(~��0:��C0�t�4*��.c�s��'��:����<A5p�z\�ux���X� �OT�Dy����'^�'������+�;C�{����1��ȱ�����Y��Ք����8�|gs�n�go��{���G䇨�%�����B��1�(ry��:oa�Λ 'v���,]2��7T�#}Di^h�˳~��U�e�p8\�V9�ݲϕ��4o`t<Q5�:}7�"�S����Gѻ��Ӈq}gF����^@���f��G��+y��X��V��.ҧ��o",B����gͽH����bne�W��V	W	�<�2�~�][����1����	Y0s"5�����ɐ"_:�p=�؄����C�Ho<��"Na��Å�
���(%X�b�q�iK�ٜ�y��J�)��Ro��cX��tuj�-H�	a����r*��9��?6���srL��H�4w�i;����c����)�����<�c�|-I�-�	,غ�N�@`<�C�>h��c�Gq��4�2s�� =���n,�>D`���'��}��^�ŏ�{G�zt�:K��z$��O�9�,̅^��-��B���Ut�ꈅ+-(6N���SX��r�ԫ>�.x��l��ѥ�4���W����M�����;5z��Y��v�C1��h�J�P���Cly-7��9���r�L���\�C
�A"��[�k�:���`�8��l�Hbr@�g�`��F2M>�V��pXJ��Я�#����������
ӯv�4��+3Y���!g�U��i����^��+�&���p?b˳��k�_�՞�F�z��-�s`r</&w�`Y��ޓ���ğa�{̲��0��
.���FҎ� L�蹧�w��2_3 ,wUw�i\I�G�x<�u�S�r��s�B_E��C������1N�
�4��~�fU�șq�H/l�E�c��¥�4{�S��۪N��T��,8��+��C$�T��DO`�Xd�_m�ψtS.K����Mq��עvőK��m��Y���&�	�g}��P'q���?,�/���9��%nߗ��yi�x�;���M�����)��1�k�Q�����ʥ���Q`P/�)���d��?�i�M�b 0K�N�L�u
��ꥀ4L�����}a,�K��x�W�H�0BzRc�L����ڈ�`�nΣ�zf�1�E�?l6Ce���;3���{�a4yRw�79/W{�g��*�emͽ�1�r���0�����f�:�Ԙ�h.|���8X�?���p�H��ʍ7~�#��iJ͒6��xy������-����|\`_cz�.�(xa����n�-���I,�[�6Ww�I�"z���O��f )7e����ڙy
�M������M��:�&]x9���fĹ��}6O����-��/l�j8����v��ئ�O�$W:��DfǃSO�R�}m4�i�k"xh��_�i��׉ wB���'�~�Y�y�t2
j\�/�d|)��}.g�����h�������ỷ1=���u���β�0��5������vw���U�;��%͌��/�Bk�d9�1�U�s��.:��"Ew�QV��f�Cy�h���f" /�ӧa|�dH)�L�FΦ͞&x~<�a�ʋ:��6F�߾�p����qf�E�o0݂� �l6�S'�;����_�r�q
��23�L�����^�',4T���_�j�SJ�L�i#+좄�6��3�2���%(�/�w�lJ��+�� L�0��@x*VZy�ʥ�g�]9������3����?V�yP��۬k�g�P��Q'�;���!�b���#x��S�@���2pu����^���?�HhHr:��E@��v�����֋OR�q����
�b9B�!����(,�l��CH�Z�-���"!6��'}U�v����-\]&3��u�����oB���_Sxr�Z����@J;�l$]�`��d�7�5e,����pH��!�z���xɭ�Wؓ��
��]!!k����2q*�-�J��f��'����Ym5���LOi9q�ms��R:��"jM��#0���!cDm��Gg�V���%a�j����A:H�O��Fw2H�mΆ�6���N`�^�|㔜�,��G�r���$��QdW`�yR�����Z<KI8�D"���|�ʟa�����VY�����.��c�H������$��r������xs�F[Ch�� ���Ը���O���+*m^�%�~�U=U���ю��!4g�x�c8M�+��.a����oJ�`g6�`n�v��8�c�r����ېNᨘ�����ot%�	��
U���~��R�}�`I�5R"���|I �|���F�;gٓn���\��!
�?�� 7]��J��O������w���N���Z�q[pW��
�@0�U������	�|�A�[��X�\����D����[���G��\���TL#�R�Gj�=�$D��k�)`|�yl�HSԻ��c��V��������ϢM�`#,7F��g���/ڢ=���,	J�Gkl���Nj��[�9*6%���_��^��n}��L���A%�`���K�h �u�6�zJ���Y$����H�I��Z%j���L�^1Q����1e�r=s-I��t^�1a���$���^�mw���ӭ��,	��/m؛g:�S��)G�5��6�}T�OS$�2!W���hw����rk��y��a��K+i6�e�F�g��o��I���TS�.�����O���F��l����c��ˤ����Ӆ�1���� �T��D�,]���)Y� ���=��``H��%1s/�����1�~(����DQيэ�]G?M���ƕ�l
$|m�].�)"����C@[��,�m�PHNA�.���
4�W�yrz8C��_G��3 �ڼa{tq;.���AD������DFhD��&����,�A[�/�z"��Ǖ���FhA@�߮����߷i�?2�����/�2��Vy���-gBWU��d��+��-� �`BG�ξ��\�E�f� �^��u��A�-Jz'���R����6R������R�5p�o���uh�ä�B��L=�5n��������Q�'�2f�
}�gB�<V���Eg��l�NL:nw��^Hy�A�H�v���s�ÂGi�e��b=��I?�#jx�1ԥ��~3>$z��p�M�>��U׋�o����.�����dp���_�e!� a�A�5��U���uѸ�_Ӽꃷ����N�u4O83��	�3�`�h�6�;��c��y�CG���W�@�YW��@���5o�b�=t]�nb��[=6(�u4ߝ��RƔ5.��u���Ը���<���b`�<�13�l������3��q��l<�����ӁŶi�5p��/�p�$F��R%�,��0���[�'��w�Y[(��4��h��h��� \���G!�OnӐU���)�)��H�ӗ��?���&�D���\���.��*������?M%!R��G��Vz�5����,�7���nǏ
Q��������Ň�`�}NYxDl^���e{{"�>P���彐����plM�7g�a=dQ+k���l�=�Z]�D7�,��T��:P!U@�*0��D30Uo㼗Qȡ�b���"�8��/^�a�VG�i�W�70�%;����~|k]��YA�$q#t�%�������9	���[p�
!��;"}=J��)��{8����L�����8�x����C?bü;�!��0I=Εyf�������9����O�* ��l��hd�p�m�zEB \:����*�PΗJ�pX\�ଽh��Lz����m?��Ȯ[2�6].8+���g�K���2��2K�Z�"�Û׌^�1ע!pY.���<�:��}V��(����q7�1��Qa.�.߂�8= <�Q���w�7�6G-�]�5p��n�X"RV$�<�*ݭ���M~p�y`U���M���<3�b�pSC��$�z�!����׼ߢ�h8)R�	c���x������xq�Tu<�Se��ҝ>/�5{�Y9|��Jj��m-ο�����}N��aB��*���W�נ�Ə�"�%4k��π������Z>�nt�UQ�s��J0[�)ke�=��%�rG����$��BH��������XqDI�����0�Smz��΃1>�+#��N_M��O���2���Sh���R@]�C���7::�K������h���O��b���D���E3��#�z0���,��P�;����K;��CA&�u�(�HM+x��r���j���X����"�T>�t������N�Ƨ}���'�I��܎���y�����1ܓ�~LX�e���x��
��fcQ	����e'9*�<e���N`�-�ع�i��o�|5!m%�(�-	b;���m$eH���+���%V��m���G��P��{L��d��f7g&�����߿?���86/�cпY ȱ�8��F	y#����i^[@L(��/m�9�a C(o�u����%Ui�.� H�L[\���/���Ѧj�Ҁ�#�ڐ�]��dr��~�F�kx]��v^�#B}�-��K�q'?<�Ɏ{ÀURqɎ�~��>�s�Ӱ��5��&h�;My�Zc���O �����1��p��M���PC_ID]���;� W��\_epF0���h�</��y�u�;Sj�����{k&a�1�J�&	"%`������
�jV|�o�l�m�����+p@�C'ۂ���p)�/�?�b�?�!����3熑����s��衻�ɵ�b���\������D�1Ū��".L)m�T�&'�>8Dw�?M�*�I���q�p�j��:Cza�2&nb�g�p�`3�ܼ�䧫�����o���׺!2��0��N�j���gUmƬ�̂;�(�������T�U���:=�Bd� ìצ���/�O��B)���d�m��t)��3�X���⥡X-�B"��G��B�y�5D.�W����B�[�� N�*��j`���%�������:�tQ�*nv����]M�a9>a�מ�c�)���xa.ސ/��g'tг��$��\YC�;70����L����<���5��@�,���N��Hn~
�>	��`�[% �t�v�F]�bs����8�A��&�lh8;e�t�B~LMv��ɦ@k<���D���*��Pjc��U�d��ʤ6e��IzL�-��ߪ��3U{S���L�����8(աے�27�p歍��o�?����>��F9�)��T���QGh����:6����,;�^;I�iҀ�<
$�4s���,p��z' �Vx��7�}RMQZLW���>�G@�dI�����&���_.�^g0���hWD�}�}7��'`�����_��WKZ͂��6y)�G`�DI>VgL�=���E}����l�zro%|$7M�Y�v��L�����6[��5��~5i�U[���'(�q�ضߩJ�85�ăBW�1H=4b@����[F!F�J#�8D��rM"� 
6\Q���� �I"��Zj�t�K^�h7Q+���i_�86Z��#��'m&��ެLd÷Ȁ]����D�fn�'G���<*�>�ڄQ�q��W���%��ެ�^�-��#�)>6��Җ1k�ֲi�h��:����W��{:Z����9���'���J��Zw�=}w��.T�T���I{�+uc��<K�ao_�,�K��w�a�d��������!�:6�U����oۣ�6��a Pկݹ��#���=��V��2&�Y�6*������^t��w!��P&�浗�N�9�6�׌���2Y^�zRW�}g$v�����#��b8�&�,���-����ʿ%�@��/����ė�`^s��͒�
��T��4����{@������A��
����c��L �F����o���9�=cO��(�UV*����h�|f�]�x���ܗ��hn_�a��*�)6ȯ�
�*�o��a �!��9]`os�u��o�+�^�hia�M��0b.���_��;ZzY]f���K9\���*���!@�3�1�O��I�t�Ÿ�z�z5e���1q=+��D��0��x��`��5��H5�m?*$�x���N'|PVE^VJ�1����c�7Y�Ű���2�Zk����&.k��\{4��u@*`B[��w��!����'��s�.Sw쟧 �_�aSs�Qd�!�;��D����Uo���m�d��	e����P��ʀ�:Y',~�T:V-&�t���w}��)������U__�s�]�7��me�?.o_g'7:�|\��<H�ٗ��UX�?u�0�O{��p�rӵ4g�W��G�ˡ�_�`փ`r��V��: h�ǥ+Ȼ� ������3���!H�m|v�Q����JA��0X{n���- ���Laze<�yE��V)�B|峄�����K/<G��,L_�Kq�&�CI��t�v��u��%�/���\�)π�'�d�ʹ����ݴ]�=�ˀ\moק
�SzXI�F^������In�p��S��ᨛ�W���&5U[P��R��<-\����B����� P��4�:��<*K�C��W��{|�>ߑK`��脸44��N�i�A�P��e
ߓx�'�²jS�`iw�i��L�!��K��K��9Yc��G�鿠�S�������|}2�\S�P�|����;'��.r\zþ@
Ag�]A�$����k2E�>�(����)�I&.R�A��i�Jm7�٪Ԣ������]��%���	bc�6��o3����&���I�����	\s$*$V8�Q�œ��6\V>�
a�o	��)37mH���~���*<�x��90D�k���;F���'���{� i�$}�Hn�r�^ؐ5�x�6A!�ؐ#
ȍ-R�Wg���z5Z^���z��_7�˳<�|��^~�I@�~4��h)ӥ�� �����B�W��m`�|�?�O$�@߱&w�ܩ���Bg,X���l�\�Ԡ.� R!(S����5$@RD�_ߋ�rZ�!D�xoo������m����P�6��:
�;�6&}^$���^�J}���CL}ׯ06$�C�M9��B,� m�����u@�yO�|��(��o#X�ĭ�q��"��E �Y��JKg{8�1�e�ma�^��[�H��=q�/�g�V�ZaNT��X�����wh�c�|R�!a�B�}��6��b�D��*8P���0��つE,"C�i+�n?Bgc�2�f;���E��Üۉ6A��K"�^~	���Ŧ���b���(9�c#~_l�(��	y�0�(�Y#i�9�$`.�L6Τ1���&����/?ף�w	�a;@<2����|}o��R�`��7�+Hr����Fa���mRv~�[�U�ڦ�Y��!���)�=S�\�V:v��if���5w�����F.,Jo��(EH��	%�;T�rj������0�=i�T���̵�iAf�hH�L\�k�#���R����`�d�LdiǬD�CׂkM�C�X�0��)�0J��ׂ���0y���}2N��������҄�Y;=�`1�����$z.1�p��Y���f��L��;R�x��tH�6�#�!*���j/��[�GWS����K�Sǅf�Ώ5��ig-�:`1�M��6<�E�x�l{YU�#�!��k�'�Z��5� �q�(a�ؘy��{6��@ -��X�؝]?Ӊ7���E���
�!:ك����HEm�K%�����.��s7�n������a�V�D2�����Ш_�fX�����]��,�]����p�$b�|K�H����	��J8�ԊM�<��� Yy]U	꯺0m�����$����L!j@,'_�����.�"w��u��F�T87��5^.)pp��xgr�����&e��A���)�"�Pn8J�A����K䍆iiǵ���,��p����uL}��,�;��<�Nl�Kgɛ2 k����3���8�G�a�$��<-&:��O���<�_��#�"?O�Ѩ�Yo��^�Ұ���I0�ԥ,�5CQ_�B��-�S���� �h�5=��\k
NQP�}:��ڤX&b�,[x,�	����C�o|�a�գN���d������@�����{NW��˼��=�Nz��
�7����{O��|!! Y_�ãIPV���Ge-�tV��U���.#C���x�͸?��:��Z��o��y��s�ȡ��SC�����|���1,�w����?�m��$�eJ�:GP��f�S��ـ[\W�K�`�����W~�0�� ڞ<E?�um�ō�m�Cql����ԯ�.����g�� �GThi��v�D�r�3�����k�κ;Y�h+s��5�g��sT�\�EY��F��\��e:?=Gwu�,��_�����U\,
�dOt��(���o8s�%��4e�$�.���V�O��h���� ������y#�P��M�xy�`*�[=%0I��?���lN��}�.���-o$��')N�^��q��nkQq����qV��S����C�}
�M0�,�ʣQ	jr�c�Ǌ�?.�ǛU�@P҇	X��HnҾ�Z����Q4�{�l�G��{��t�	0[�??nB�h����?w�!��%������+�� S�Z�͂Ѓ�C�h������P��O#J���H|��6���O����1ȓU+I����w��0��G`\����͑�i�f�ľ����0ɭ:`dm���$�Ce�W*H�E�3���V���M�z%��[��A}�j;NO��N�xH_���D�^���K;M��ה���[R�ӓ"<��|c�G�?uR���D��6�Y�A��]���M�q�NI��@�cv���� ���9q �}e���J���o�)TB���+{�%Mp
�3mX�0��%m�,<��^����0��&	���V��]��C�I�wO�b�u�B��<�J㾛�̧�[���v�V�f�ld��2;6X�?_v���|E��Wt�]��舋v�k� s�� a�\#1f�Xg��M���t���H�s��3;�����N�ɞ��F����~�A`�c�s6�!��j 8��~��3�=?,���=O����C�7�l��)��N�E���d��U��b+��a�~��_��Z �q�W}r&ݮ�h9o~�HQ�a����s臃�1I%��h�X��mU]���j?��\C��F�M�:E.��. �C���1������Xq,�xD�Ͽ ���iG�$%��OT{00i�B�� jxnX�ݝ��j�b�, ̓�.��g�j�A�6Xmk�g�ѻ�d	��M��R��o��l�y��9=�eUߗ6yW��cp�+&���.����˙��cg�ǳ3��$*��L.���ۏ��S����F�c4�s5\�J�l���'���iXHd�E�T��k?���Rws;�#�++�{�jUv�<F�#Oӝ���ZjA6#F�����PA��g���F�l���rs��*�B�A�G���+y2>��Fi#q����:��Í��S��8��4ɝl-U���H��� Y�-�(�vR����`�| B�+����#�� X,S^�J�yጭXY���Rs����% �k����rz�ęo�;~
uq���6�[@h�,^Z4v���n��n#:>_�A��f����>�s���0�a
�+��M*@�6�����4�c�!ED�o�;(�Z��"���~�������b}�i>���@�����Xp�%����R �~�c��1�$�1r�O<��r�-�w���s�ˌ<x�!��~7�O{�8�u�c	�u�=�����Fi��#��s9�/tB^Ԕ���x ��@�j`�+_���ȁh��x�S]���dB}��tI7�����x^s���af�7�o��a&�j�T��\�➾�9d�X�:#|ϓ�\��w,�#U�����ݕ�iUX�K����&W�̄ưaC	R�mZa��)�@5��ֈ=�[^62B�p�.�5�.��s�[�50�EY�S�����g2�Bg�m4�;��������
�_0�f�͖�?��%�jj�BM��Z�����D���	X����x%��p$�\���f�rDn����Km�D=���&N�(��y��b���SW����&��Y4��c�;/����4���߃^��ԣ������4�`��F<�@b��Z�[��ibsw�V�2x�xD,��88(�����&>n��u6Z�J���~�>:C�zB_�.E���Z��3�9viB���x�M�Erʄ`�!Yw��I��.?ET�����f�v��k8����%n��uv��P���ζ��r��*˔a��錒L���%�yh\j�����[ǽ�=�;��Y��4$��4~�b�������G��bM%;��Ngq����(����")���/�i�_]O��0!{Ŀ�>���}-9�l�Z�.&5���A�JFr�ueaA���#,��5I�������X���I�߼v'��kHQ�$yڞ��Ⲓ�`�-S���m#A�@ޯo�9�6��݁eO�o;�GM�h������p2Fb ��������N�"7���X&e��nΟ�[b�z�9��i.IfF�L���p�/��sr�N��9�����=)�A�J�LL�,�M� ��N�m�˘���\���W7]n��b Q�?�*:L�&�����}�v]r��ɴp�	�%0�}��9bV�aS4Ya��ā�.�%�����'l̴������ps�VeS7�r.����,i<�/���%?,�"n�ζ� ^"q2�k��x���|�9�����g����xf�ǗՖS�ݮ�Қ��=�%����QzE�$�z����I��e��f�(��K����#pȁ��X�a'���&?P���=��ӈ���!Z���b�9=�7����99��Nn	��U���Z	�r�Z{�5���_������&�ą�X�U����{�M��;L��ޱ0�ne"����5�YD����c3��1qH���'a�U��U1��R�P�"�l�S�3i���t��&vt�ͩ|>�xę�.uG��/�����E�[]�*��XiE3��JǱ�1m9�?�T_�+/��Y]�?P4w�nY���sz��[|ٳ6�w��ZM�Б��c4��.�165�����œ��%�[��4?�H��Dfݓ���l{����@��)I]��DB�ኈ�)
�S�������!6/�a�3a��G�����~��9�b�H2��2�%'�S�R�f���uO�Y��,O��E#���h}n(�`o����-��
<R�Sbh�����O�(�<�d>a���Ĕ݌6$Wh���
���ނ1���TL�=�īK����� 0wC�����N�-�M�!���OQ������b8���m��PCP�EV����q��/�eÇ��WO��g��"kEN��C�ļN��(�.e��b�u�3��;Gz��n�}ʃжU���;�W4[�*�VS�Y�ϰ�[�Z�y�N�N� ���sv}��Z��Oѽ�J�Ն������!ef����g|���Q���]���G�i�/��O��3�h�ac� 'a�ǒ,���䆱�׿˾	��;���!`��6�N��\��%}ѽ�l2���?����`���g��ǿ-�#�چb=�W�E�+���v�:|�ᱍ���	�z�9][&.,I1|�� ����<A��F��'�>{l-�z_���VL�D	6*��E߅�U�e�/Kk��EP�x�@��S��g� ��q��S/��$�4OgJ2��c��ʲ��D���d�Wx?،��W�1����^,�+)�G�L���u$zk��MA%����\�s�-$sԎȘ!�i����
6��;���@U��4��2l�������&U����d �c�9Fˇ.Ouv�E���z��B2;)��p2��,��D$�Ɨ����� �/��@i8���(�P���6����+�e��V`��3v}��	(�29.B:>9E���G�a�h@��m�s_�M���x3�E�<ʱISw��k����%�VX�W��#2?��7e-�sP�B��A#d�}���W$�M�#��x^[.4/%1�P����aHiή���&�(��uyWP���&�m��!+���qZ�l��@z �o��ko�q�&��V_����hd�ک$����,�b~���|K�Y\���t��`���BQR������#Άr�Ę����>3�����#�c�<�m���r�imC�y4t��Mq���c��É
�u��'VR��4w!b�}-��Oܦa�ԫ^3��6@��&Bh�蝠ȍDN����K�M�lW.����X&!�a��~LW���Ƚ�o&����*<�������M�� �K=I��O)��H�3�V�3�1�7GtŅ���B�n&�(�	�����e��Q�dl��o�x��87�:1�YJ�s����~y1t����m�b���<�y�w�n�k�l�N�&J���L�j�R�f��dGX�ãMOm92E|/ ���dIg�/�87>Ca#����ya�����j�9x����>��cm�dg��\�H��f�F��9ġ;0v?��q:&���?b�8������4yF��5�۝&f�~� da����� 놩��������-=�}� 9�D��#;G�eUZ�'a]�Fg�bB��h�8U3�1�O[�0h����h�k��G��>�ʋ%�n�
 ���d�d�򳏀-~ q� �.c�K�r��Y~��^�"L�'~�'�6��|�tt�4FK���'Ze�Nx���R9s�Ad�& �[9)���[w&�E�:˞&��n��u0^e�1�+H�;d6 �Т?۲Cx����{a�7*S����<T`�)j.�>����P�(�+��Ԝ���X�h�����z��wx2����2՗�ON�}$-��������J�B��e��;"��<#���\l�(�������^�X��!���I��r[�1 ���m�)�<R��k_���	3S墙��7U�'U�O��]��Y��'3�Z1�s�J�tu��͈����,����t�CZa$�˻/������'�{��@-�4�_����+�(�Q1b��k��Au"ۯB7�=�����d���Z[�i��;��q�� �8�^6��ܡ�`�q1��΋�+�7r4��>�S��-?�E��t�n:�ڼϔ6>M���� q��/�1��[���O�/�#�����
�I���e����|_��j
9�EW㗰���+����`s։�ɡ��9fM��6:��h ��?�T�4��O��R�J����_�=�M�mϦ�@x�%9��2qͮ_VL��?4������F�5��l��8Aݴ[e���Sjb*'�Ne1��Ck�]�昅uVj[P1��L�wU>��Tkr��"�ZAw6�Ꜫ�r�{�苤�T�N	g�'�\��A ���9��hm�ͽK0�%��k�͓�0�ovX�v�Ȑ�A����KG���1�U�U�}l���Zw��m3Y�kl0�R��ا��W�3A���1��=�-���m��Sz�ǅP��%T�^/��S�ޥ%���$ju}��4,�H�0,$�,����+3#��2N��\��`c��t�%����c��U�U1e�Yѫ�A�7���B	|��熁���{�a��Hm[{p��fP��(��!���
*�02�!�O��5g��rS�*N��J�,��L�Q�YD����'cx#Ɗ�����rm�D����=:��d�����ق׻��ht�& W�}��}����߯`�&�������.��T�Ǳ�IԷ+pβ�WP�W��^P:q窙�԰q+؉>�)
݃��SxG���� ��v�K�6 �>�@�6�#�v[�_�y�7�,�l�{�����;EG�N�U/�*��؁�����tLw��c_,|�ҙ�����d��VS�n-I�r�NZ�٤�W@
�=�y;%םg)+D�~�t��- 
�6K��k�Ds����>W�uJޙ�Q�L7�lܰ9����(��4�}�A���
��F
Z\l'"]SPm�>��ܘ;V�	��@���K�2�_��<�U�ؽ��􂳕��!i�̰]���`�����D�v�lIP|�S��C"�Ja60	����JZ����/QW�?��\BTecsV�ݛ��q�������ۥl����c���^?���s8������Y��i�����ZSt�i���O���w� 9c0�������f�{)�`"��6r~��s)TU�-/�7���^��ؤb�R�'�)f�(�\��MR��ۗ$��Tp�i���bL��z�-�6��pQ�$�ېD�F7���)t����"j繞�<Y�5��.��Df�X}����҈BD2�~�Lc��h=����VD���)C�_�3 ]��,���P�E���^��k�]�pH�Й�m�go9k�AwE2�P4ޘ���"���@�ڢ�̼jM 잂=�	�%ɔ�{��I�~��m�6ѬX�Sx�u߾vN{S���L����<�����>�T�B
�"�7>@�5�4W�V�ّ��"���	��2-X�����>���A��8�ϳ���Z^}���lR���(���]�l�)��*A�ӥ�$�K#[_N���Tot�[Y0ӈ\��L&�F�UC¬s�eJ#�.��t&�>CŞ뛃w��e�m7��{H��	x�FdNd��s9\�s��-H9�ʋ�5WC��Ô^98 ��X�T�^\�]g�%F��E���Z����"/�_���\]ZZ�z;����4�ZBB)`Vi��CE�S��:��Eg�E=�?y�����x�����izA�񸦷��xx�j������#?+�G�ן�ǜ�k=�8�V�0����dO��ΠV
o�ָ]�*ѧ�c�� 	�$��m�m��~�k���PqN�+���g��T:�5��0������V��%�IOa'���k�*�r�ݐQ`��Į��g�ʤ%�9����"2�0���P���Xׂ��G�?L�oi�� �?����O	����,Ȏ�Y4	Q����%Rq؏x���ȡ$.�7��	�A�JX�:G�K�R�$C�X�X*�J3�Z��X	5 ��c�Q(�pym��rw,K��~1&����e��m�,����bGl���%�wU&\�+E�ᓇ?��jOwF7AĂ#�0�LTr,��r�L�S���n
"�%g�t<͠3r����-� �?o@&8�U:d�lpK$$E�9SD�C���� 8�f*����ݱ4��^c�����:�Ry�s0k�ᡗ�1�L^�t��+GɌ�bH����Q��#'b��v�D'1��`+�e�):�cR�j�û���	��Yw�Ì���I�q6s$~�rU���L<۲���p(�:D(Z 7�˥ݭ	�Jx��Wո���۪��D��߂�_�[��0�U��D�!�R���Be�H�Z��Jj�@�
�9eb-��@1p4�y��G:<0J{0){Y�UoY�o��q)��B�_�!��;�n�Mq�*���|a|��β�ڦB
n� ̠�V������*���/ n����Q��!��Z�YшK�o� ����e��5"�_*�7�|�n�^hg�;�ɚ��,k)��:!麃�z!^��}G�����(��8\T4,h]0�����	uzy��&`Ձg�tCJTП�~����,�O��5��"���Y�!1Kr��>(���ˬ�r]8V�~������h����O��F��?�׸��Ɂ^¢ְC�F'rI�g�@	����˩ָ�m�#� 6 {r�k'�ur&\��#&����X��l��9��Ip�J���y������Q����Q#-�M�w$@������x)�5�čcn�A��f��D����v�k��������b|:�nk��O)RP�$���?Kt-5�k�66�ׄ�p�����>���K��{������G����S)��짎�3r˚l2-8+�X���2"'X�Bi��6� �!m��V�m�@�����ux�����9T�A���[f{�o��!�� ��]����fF�gެ�AM��t*�m�8!X��0�m˥R�HR3q�f�v-��ƶ?$W�����R�W~!����ci�j�Y�f�²�_'O��\��G�Nt��򋄐F��I?	�Y���$��X�[N��@D�P��Fi�~#儓���Z?����]�0��'X��ëҡ�x=D�}H0��x��ܛ������Yޑ���+���h�3�fB�!AЭ{�T&�V��&��t�� �Γ�hV�d�<�d�9adfR�f8Ԕ�P���*.y?�(w����N����i����2ߑ]D�x�Z�~Z��1�Ac��-HT��x�q G��[�mN��͐����MJ���,Ч-_��s*~�T�^6�-r����B����T�=���7Ux�QV��Cp��bx��]L�bmu�n[��G�H�ѲHIU7��q�/&���.���e �"#���u�Չf�6�q��2�n���v1h����|I��3�t���
�1S�=��i�.��%2䘩�¿gU0�?�ʪ8�}��@����s~�(F9��h?�>��coX�3R8�lqO��9/�y\N�u�؁p>�O�W��h��t���a��㚿~��� �7{<��!�	�7�<;����qr+�=����X$c�T��l�5��*[�ª���9����K�ڀ�����"��A��#(�����;��)�bNf����Uq�IQ`���N:�������V���m�/���UvA���Y�Ǩ/
D����( 쟇	ٲ��(
R�C$'�9Pg˞Vi�s���C�?�d��`�<ǅ�w��S^��E�b��xc&S# �r����<�#z$/���vfut������d@�1z���1�E {����2����%E˖S��XC_��E$6�u!���檕 O�k;$��KHy�Ƥ�g�'��
�^k���6�����3��x/7�������̀|�e����d{�A�u�다�g0٠ ��B9��4�֮}����Е���m���޷X/���YU��F��<������U�A��AD��o`H��Iv?�"�f��g`A"x��`��|䇏�"�BY-�V^����Qv�����ǇH/�%���0��E���.C�Z����G�lKG5�:�(������ �bCx6٭2���#L��D�����"�ʸ��=4���֣�őo�A9üP2�q��ӛ�'&/8�QԀW���=�ir>D�PQ�U#gpz�h?��qTSnƅ��oS�w	z�F�q���_%�l���r<�/E
B<٤����x9��O��'���DJ�N��Wt�m%��*@�w]b���,02�!%Q����![GZ.W,�WG^|A������� ��a[iK�`�%��x�� L���!w��q-���c��t�"}�&�g�%A zR��,L,���MX���h�D
�#c"�Wq$���y��A<f�p�3��%�1���X����!��kF��f`F��҅d� Hn	3��g�)U�Mw�����#�C��R��9�Mg��-f�HA���ؐs���hv�7	{2��9��3B(ҕ��.����Fi!v�wiUӟs����u�4"�:�uQ�ԀU7��7�ww���՟е�9�Ob����p��|��#VF�+�%�8�i6�u�4pI�i��p�(Y��gɇd}?~�s��\�0)��-@��u�h*
5��������Jo$臬��g��C����zO����T����xz����f��U�6��U`��5%h�:�4b-/�SZD�!Mu�YX�p��_"�V.����>w5��`޼:�Ӽ I`;7��[.�%Ց����Q�,m#�L�ɕ��������:�
�Ȯ�3�!#�1KՌ����W1�`B�O�dB/��1�Wy��D"�����;�!�S����{u>I#����a�i	j�.W:E��W���z��I�E0O�P�����ޣS�S��"��~ �Ӂ�F���������X������=$�VE>#^�@�����U��l��DZbp3~�b�o�qV��7�9]*(wT��g��_�)��K�ͩ� 
�7Mӄ~VF���3 !_�OQ�|�dF�n�<9� 
�Gm�R��r}~��t<���''�s3`���$�B�_�]���EM���1r7Ҙ�D��]�cWy���~haY�q���w˹��}y�,�x�z��J�����}%9d��h�U��J��-HZ�<���@�k���*���[)k��B�꛳�;��W��-�6/(��ZFh$ǯbL�錖���C,?��-�}j��ڑ�˒��a��J�s��S'���Q�2<[��1�H(-�������f3���lH����>��@��i���a�*V�V�W)�V������E!�`���dK���ƭ��ۛ�Ȍ�W6_RA�y4K.�l����O��N���Q����xiڕhȊ"Z��W$rkBC�4��/p���[ey���wL�'B]�,ۡ��紏x���L��&�Y5Hҵ�>CF��cԡ�m�4/�6G|���B�b�R�򻚟O0(h�*�Q���*f|-�f��z���$߰��_�Q|���S/$e7�T	ީ!�1�]/md?��kM$x�� �)�)��%�G���Q�*�Ĝ\��u����n��w����Ԭ�y�53!5"�e*�0�CM�>2�w�o_/[OZ� S�Gw��e�dKp$�&�x8U~2Kk�|�}���M<z)��˫==����+�ix�#r�h���U�86���b�v�¹� }���s(�)�^�kW� ��1�WG[��x[Թ_�����ޞ�5!/xQtwt����^K��(�rh[v� �(�޾�->��������Av;!	�ն�r��[�(+a�F� k�"�𔵟"�ʦ��-Ǥ�WR���#�r%�6̩��w$�]�(`�&�	G���^���7>x��E����g֍�7���е��1���������P?�7�%Ӵ����s�!������nw`��%����l6���ARZ�u�w3��>a=��P�(���׶\�)�w�7M��F����h���0���=m� ���<�q�5��L��J�D׆��_�Y�a<G���+|>2�uIW�/w-��������j�+ݚ�U�xP��y����y��İ���]����6�d���g�h�V�[�M��H���<�M[@��^^�UU��R��c�A�I�^-no�O�!�Fv��H��SCN��q�
���s��W���I��^�rc]�.X��m֓nw����ˉ=w��H}���`��;�-�a��-9c�0�гUo�r �O����EԼ( *�+h��gJ�E�}��l�XE�q`īX�ޏ�G�S���`2H��=�0�#�J����g�%k�>������b=�����it_��C�#̦Y�ܷ���Dh�Vsvh\���8���W���LS�����`�]�<	�{<Gƶ	����P��BQ9U��_Z!R��61��;V~Ƶ���x8������Im��9�)��P?�tQ ��A��FYL���C����� i�d,L�9���������"Z�y��泹��n��Ơ9+�]���*���/8@V���=OF������w�T�ze��ϛ�p��2���b�D���O��j�#%<�S��Ͱ-�h(RLѻ������,�������u�,��PB�1�� �zz_K�	��A��!b�s�+#���S�8�rmF��evxy��g��]:7O�՚?��gx��`�I�W6�Lz}�9�n�/��tX�}�,�XT��.�������h�b��Pĕ�c�ƿ���o)��|t��`~A��$��� ��Y+]y�Fc$����g�n��J3�w��,�F�G�?��~O��	Ǔ:Y��S�"��x��?�w2y��&���>y�I��*�5�i�B`U TA3���?�D�9��1�[E�ؼ��9�=C7��'���ٽs+/���E���Ӣ�Y�4!��Tȉ�J4 �X|St4��,��,�����-ہ����H���;3�I1�������L�n���Z[�KO_�u_g�p�(�c%C���`��y�p�\�����`cW̘�=_6ә��+�Mڎ�F�2�`���\��p�*�4|���iFA�����Kg���~:��xu1�ˍ-�[f���YJB"署�*s�tF-�������xudQ�=�Z\zaQ�����N΁���ȍ�ހ����{o���Wڃ�Ґ���>�LG�c�#�����ė~KvH+Px��&�X����C��A8e>�D�6�`W�i�C���Z+�KU���p����oj�S� �������)�v��d'��C���
�����lV�#����p
v#�/���!iQE#:	Oި�a"7U�H�;zr?ݷ�J΢�`�tTZ��� ԇ^�5�R��� �KK��	kל�s�b�)��#��Rs�/	rZ�G��
P�ҡݍ����siJ���L�f������m��N:��K�]Pp��y	����Vx{���+���z���ܣ�4�����d��3�P�4�d�G����`�h��Q�_�5kI�܊�Wpʸ#
����e�:,[��$:;���������ŤҾ�4��L��������	5����j�䙗�w.��ƍ� ��R%�5
]?��#}����A��|�g|}ċ�;�f�����]ˤ�F��0F]
��cp8�����^A�n�k�W�5$�L�ym��9��� $��H�����K���ټ��IDl�r͛qAO�r|��_u(�U-{R�"�Ԋu�q+cv�DK�cs�<�>:3G ����>�#ҁmqZ�@���	%�H}>��l㉰���xn������P�!&��9i.��-���{�?�x�����M��(�_�e���֕'9�ێƩ�	T���7'A��t�0��t3���&�����B?�J[@w���Ԡr�Pu�[U�&��_���-�*���5=E�����d��+����a�k�[l�R���Y�m��ǜx��,N*~C��|J<�j��e���KeN�\~X�B���f�t$&FVa���&�'Z�8�3M�QT�+��5�}_%���O�[���@�_�� ���������w#@#܀Ny�-e��3�^�X�C�܎8;�ػ�ؤ�_������/��b�y�}G���4`\D�0ڜ�&P"�}B��b�j�"x#Қ�儌�f��4�V��&��Z�+A��x������r���۩+Г�{E�\sƾ12���4p*D���k�'��;L�$�u��.���6`���r�To7e�"/��	�5��5x�є{�Ci��텯���j������.��L�܇z�'$:r�\:�KK"H��;�ߑ�V��|���*�Im6�i�e�g�|"F
F��`�����A����'��x�f���Nd�.�������7�c�����z�� M!���w�n��d�0�Gׇ���qZ(B8L��>���
��U�KE��Gj��)T�q��O$ur)m$�*�ឤgP�Fm�}�"S��J�-<X�sr�w�AI��D��Զ���`�ĳ'�n�A�ε��*z�0��l#�ȁ��ZWg�I|oW�}*?���DӤ�ww�]����1���X	L�\�� k�0�>f�\���a��]��>�a�J}�@ZF��	R�_&Њ.�f��W~d�lQD�;����#�[��/�0��|&�M!�����=-�#�xҥ;���9�#���1a�u���xZA6/vob-�7@�1�G�� ������SL�D-�Zf����
%�Ax��PR~�$qid��kؓ5< l����������TiU
��E{���2P��C��zЙ���Aj�H'V�q��\��0�������JD�c���J�쉲:R�_�˛k���k�7���Kva(����Y9r=��Dv�B�p��m;V^'b�7,;�wM�0B�������6I���j�G� �Z�e��BVg�)@��[=�]�%��}�u%��40f��˅��/�����:t��3_GR$��Tx^V�[�I�`F��_�~x�6\�GF�h\}�5�O�R�����G�I�o�5���X��J`�f��!��71����*ZU�=���t��"D�	_9�u�,e
�Im�4|$��*%�⬱�PTq�EӀ�F���ǣTT0۬�bx��'<_קHI�B�v�������8��Nٴ1m{�l#���q�Bn^&�_af�V�=�/Ԃ�nL!tg����{+\tț��� ��ǀ�H˽�{���՞��%M��ZB�X^�Ň��#���kH��H�y_A�� @	z��,tQ;��@�;���w��ya~�t�R|4I_�Gi��'������7W/��ġ�BW|�!���e"�m��%8K�ڶ����ZPC$`:���$6V��50�m�������\84����y��Wo	�)ͳVm[��d�M�V�L��vP�����]���h��Yշ��Ӑ��o��}�$*��#�*=����N�R�{�UPqC���@��k����ܢ	;s#�,�T��A<�o��&oF�i�5�F�q�|��E���&�����
3�{�@a��u{;��;q���>�����AxQ�1�}��{IY:�"s-���|W}�'��F����qN�hU�q�3�i��#������z�>ZR/�ڪ�fs���Q�Y�P�T ��Z_]R�Nn�/�w���?Z8�p�Q-а�+�F�?'e$n*U�9�t�9�bL�H�؋�X�s�	◷���b��L��*�����R�rC�}�_Q���'���l�
DnKR�A,�Sn1����g�+�ZyE�E�A�tā�m���Q��2��Y�d�^�La���z٦�X}�`�O��}��6(���	�2ڀv;�&�;��TĤj a�Twx���~�p[��9C>�!�dV�d�u�ܫ�%s���f��}djQ���7��	�W��(W
e�h8�A؇b"Q4oQ�dOդ�H���'�n�v���Ĵ���sń����i(-�|Ǯ|����H��跔|3UT�񠳳�|�\
!���4|y2��:����Yo�F�k�`�.=-Cn��Tw�ܣ �[?Y��y���#���p�� ���X�M�@��]��! w:S<y镆�|J���#�p������-ơ�"!��x̬�Y�];AQ�z�`����w�a{����=�MU��^�l��j1��T�;n�l����� Ol2ck���N��K�V��!�_Q ;�sM�&F���U�T�1~�ɛz�׏�c���\��lZ�Ĉ�0y��7��Q�у~P) �,H8)?(u�t��Y���l�h�Ē�S�)����H
b��������9r�,ع�P��-���;�������U�tA�C�0{@)�ǔ�ݍ6֡��#+��h2���Ԑ�6�M@�F/ŧ	.��Ԝ4@)O8I��ch㶀u)�Zޖ��s�Zw�A�M'����b0��5�Qq(z��
o5#9D���$+�}%R!Ɍ�����(���r�9�^��&elذ�Ӕ{����vs����Q7���N�����b$�^ViII�:s
W�HO�<e���W���/e���lP�ʁ��(�Z��[�����̫�1�^R�����U�ݳ)� \�M�?]���ZABε�
��ɍ�k��ܳ�Ͽ��^M�*�e��uV����(�v�nE4�y���rf^+W6 ߇�	��}���&���Z%���m���w��d1P�_֗)S.;�\�qUk_PuK4�¸PLNEA��o-��{�
&���^;UN`�i
{�`_�4�j�D+�_P	�5���\���rj���#[Ը�*����C����)JN]~���P�U��qj����ڲ#�(���9��s1���u�ē�6S���?�tA:�m���6Y
`]0>jٱț}��Fz̠�˯p�ݡ�.�h	0GR��������4�/��ro~uz6I� �ZF_L�xN( �È��;���ī8S6�#͈�zܗ��[%�BGe�b����PEN�S�>�Rr�ɍ7|s$ΒO���B�����D�" prkp��b��	i9G~<���'��P=��;�4B���Q`����Z�����![y\�Vl]h~�͑�d�,N<�:ߔ}!F�hH�I-:����%$^4!�D���;,�$�qm�W�K����V����Im�\���������)�z�y��>BY��`ڟ�'U2����0Ƕ�Ug��l�<ʗ�G�H��a���k-s��{���}��#H�+g�2���d�`�"6*����|����7qv�;m�]/2\衵)HW�\٭69��)���?]9�#�R�BC}ƺeA����Mu%����eW�ɍ�>�vo��8}qo~�7v�FF�U)���W-n�u��U[wq�<��N7�0 ��Ph�0��x$qj�%0�+������|���k8����$�U� ��Ұ,��m*U�ר��VJCȭ�u;Q<���@��f�z�o#L0fQ��b���������n'���Rk��~m����a�hy0��*8�Ѻ([���cr�Ih.��ZrMLoi�K�ޣ�=��y��7t����+I�pY��W����������큮N�b��� ���$\���f�A�9�j������3�ZR��dl;^�����nT)T���O�C�'�P���=<����(8�\�Y�fJ0�DV�M6k�"���������(�IBG),���.;�gnCt�h�^GYD�Ee��HGo5f�ń7G��t`�Vb���@�E'Q�P�Ų�~_{�/h'��^��"*ӱ��\���kU����}n��y��*OcYu.<�sx���źR��"�8�Ҹ=��ṝ��jCɝ*��jn��S3gG��b�V����<�rr9�cZ�� ��y���~�W�� S�u��6m��I4j�e�	��ᚑ�"�4κ���>����S��o؅�P6��KBZ��j�#՘���ވ�g��LY_Ȏv=�Qه�U5̸���H�g�ǩW��'��buSJ�n+��d-���W�h�A?�{���8���Vo��5z-�F3�\l��F��J�ղn,�ԧ凞���=
�8�i���9V5@��fy����mTc�5�n����{=�v�z.��%��r�st0�l�R)���=�Xd��o⹞�+t�8
劐�V/V�4m��K�'`R�������,���9��G'����Y�D-���뻀vY\�
2�]v}��pѪ0�<r�m���/U7�.���zW���E��ok��Y�L�Ncv!M�DZ���k� �:�|,�&��o�U��W?!f�(�_�>#D0��>�k�����1��5}�%��$�ocL�L�������=H��oO�3��Ԩ9����O
i������1��l�P��1=��'�,q6����%�|=P@k��B����J%*�Ѫ��m,�d,���f_ZM_ݨX6u���	�*��|��f"h$|n̙�Y�������ܡ�L3�34�l	|x�-��[�+�l�u�4�����c���X� �� ���YQ������nБ"i��1�to���!�Ý��ǖM~��H� ú��<D�x��	��RK�B��QGU��tr�w9N���mU�Z��B���l��,�$�����i2S���0s�����p�i��I�Y�����h��p�k�Sm�5�yr����Cw���!w��.T�ר��c:?���Z��e������<��$!'�`���T1"��?CW��9c<V��Od�k#4��#AQ�;ֽ����2.���vYл>:�����n#���7q���]}��ʡy�a���A��
��T�"��e4S/z�t�{Z�b靇��|j�O����k��p�ꔌ��ӣ�R_�4zu�R�x老����c媌-e�50��k�Hr�s��"�H!5W�)��u�)Oc�4縡�\sz��\ #�hms�V��#�جT6�RelM<�-9�V�3S�����oQ
Dœ�,T�n��؛�crP�ݵ���ݎ�$0B0=.�wN7ۙ	��K���X�`�7���2T��6(���B��* ���Ga&���B n�r�-z��n���K����h]�ұ��Q��y�Ϗ��%�W�߬�d�4D	]~�K �;���:0�`f�9��4e���H�{���%F�cy])��nF��kqd$up��HZ�̘�c�0�tv�$Uq�\b������e����j�Z��!��~��θn�*ޙ�x����d`�]�R�̶K������np+7,�Aŷ�`��Eܦ�]�(���'��Y^�uI5r+��O##���W�7�����������	G�%-�Wo�`�.�^�PH�^B��5tѦ��cqa��hWL���L[��X�u�z�W�5ˋ���(Vq:�۸㷱#P�&W?uZrE��!�9�~��S�}Ҁ,��y٢��V*8�u�h5ˋ�K!N��H��'w�cVٯ;��<���WY:����0h���ŕ�W��:�Ǒ5��e��R�U�-�;����W���70�����:���d��fw��ϒ~�W����t8$	�/@;0��2r����_ht�������j7+�ਪS��~s{�p�2#�ݸ!��
�>����[�!��iW�`m=*�_L#��?*�҆TB�AF�E���4W�;h*{x�u|�!���U
;��n[W� ?(�LF����u��"F� ��rMEľ�SC�a�B�=�#q��~�D�~�h/'������&�߀�-� ���3H����a�!�OCW[�F���i.<c�^ɩ.����	�@�xI7[C�z�M���)�n�mJ�����p�5W�C�8�[���JWP*�	_��dkHS�p؈�\>���rE77^T��/O2R��"�%�p����W����G&b��ɕQ�������Cn����5���e��Q�vK�c\�z]u�|�|�<٥�s@��߀g$p'��&m��i�� ��0��[)*\K�<�1���ܒPL*�[r1��ͫ1Ymo.{\�H3�]���\>���a�`
��[-�6�|YYȫ��0|֘x z����YK1Q��$&�U����%�[��s|-� ��PO�4#�Ș \�����W�[��Y�k҉��z"T�Tk6�Q	�AA'S8�~����� Hk X�v|υ�:���e�����o�ME�wĖ� B����6Ը�F���n#�ߺ�H%��,!5������~�zD���?��	`3"��"���o謹+�lW��>,ʥ|r�8^�(`G-'�o��T a�%� m��n��{Nb��I�~R
��KX�T:�g^���Nq��.��p�ݛ�����_L�@���6S\.�W� c_6����J���宕ލ*����GW�Zb��x6oAOu�涋N�:5�W9�l��-�9�!�*�Q7W5s��}JW�2�l�Oy�1
	�c�"��U�<h����Tu,>&Sla	0�]'�v���!��!6�z��EX�?�.ջ�i��%l��^�+	����#�6NG�{%�^��!��,���gn��s����F�&�y%/��@���!��l�#��O��/�Y�����{�P`�?�k���� k�B�����_�H�\q)�����d�`�����:K6��s��7�/ n�U������r�^~I�:�zc`鱛P�y�B~GR��g��a-b��n��\�E���>
~�� T�6�[l�eU	��a}�ϡZ`�����ђ�|���}����K�X��� BMւ��x��}Ԇ�7�մ�U�Sл��mjA^wA���*�]٩X�΍2����(�����;r����c��Ce�����������B!�X�r��x����0��M���>��h�/��}�O�l�4���]��̃&�l{��O���3�%4dQ�Hv(H�*�U��SI���V,�3�~���<L����L��^�D��
�e"�Z;�\����yhI�ď(�n�)�ƚ�ΥeJ��K�w=�Z֏(.��w�=7g�����B� 1��Qb#-���Y ~��G#jD�z��Pw)˾��*ck�-q�5.�<�8�0�����^-�&�	rh������Ԋ>�Ş���c��q����� ��=�3m9$���=�g�t�7ݣ�e"nU�q7�B�6��W��N��U���J����;�����}�%fk�z��%k�z���0�`#�&�0�k���� �Z�� ����x^�(FYG�j�ؽ0��倊���<���6'O�Ei��ng�2��q2�)�Nk��w%O���ٝ 5C��xh��1C~)�p����mSn���R�"�!�h�FS�� ��ߵ�O������֥�n~5*�z4xk3' �*M�-{G��ė�\6b���Iʍ��qpL����_׎L���$�i�6�Ua6ƥ��'c�BÚVAh�	�xUg;�x��h	l �>�q� #���7u˴m�hL��b�t�W����ʴ��?8�߶��{+)w4LVӫ<��7?Y�Q��5�R/��hM���EOӹ��8�9��O$���\k;�����}.p�;JGR舰�������^�'^	� �j�e1��_%�&5ӝx�Xn) �����"=�\��d�˹��ԅ=1��������B��a�7��@w8��@���jè��kJG?��҇W�)^-�~O�����I�6�ADI�$w���^t~���q�d�M�HTv�����f����8`1<q6o{����Պ|�I�Ԥ��Ot6���s���A��������G�vy�p���v�Ll���u�r1i��Xx��=�t6�ɗ�Ҋ��ec� �&��ī���B]Wh4�	�uvR`o���i��Z�!��Uxr �U�=��I6{"�(p
W&��H8�r�sty{�k}rm�l3g5��Q}z!�S���~�����C��B���ԉ 0�7�0�C/����zEH��"���/�x�~cj��Nc}D��cGL�����C;Ư�G��	���<s{����2A9Gm��Y��UI���Ш��!���ϲ��[�	R�G
:�S~��L[�\�Dp�PV�=�8=T`PŒV�X���q����j r�Tl�
u����E�o_�⓳Ɵġ���RG�p���d�'o� 1���h1�����=���)<-�W�{hY1�W(O��������[��|�:��R*�����Uq�р��H�K���q�����H�����<6G.�\K�.*��*r�$��h���)d�	��������!�zP`F�@����
ߎ(�ۆw]�;�a�y|֧cƙ~���ZAsX���)=c�kui�Ms8{�K!
浹�F���Y�a�63!���șCdꚤ!
R��~(���xr��ndR�~�(Z_)Ĵ� =U��8��B(q�$�L��n(���>���m��� ����&>�M�#��p��eC����v"���*��Q��QA�����+O���D+�k���SN�Û�W�X���zp6�*1�� \`���H����󜐪T�WT����I�\|M��3%�7�Z`b��柚�t��HUw�4�%�f�e#�������īt)���"���!{��|lm;�F��M�vW��_ʹw���s���G�]J!�z�	G�`�I�*}��QX�6�(�F%|ǭw��kJ��]�	���c���w����~�w��T>���>�<�tp��0J��U}�4\��,�4�9Bvؘ�?�H����,���y��[�*�߫T�+b�yJ6u
E�η�v5x�� R�4�K�R_來����¹b�,�|_c�./.6����r��]�Ә���5Ъ��WW�B(D�*����(�w$�g�)����i�K�
Ay��_��.+WAjcp�Z%ĕ4p<Gݽr��.����R%%G��i/���C��s�9^^�[�;Qy NX��A���; ��Õ�ot[��N�Hu�8C0��4�H����X�c%XD��("���&z�ZQ3��̅h:���������h�����0ZSI�߳hՇϙf����l��d������^G��&@��0����@�;s�"���-"����!�%,�͵e�K(��g�r��z��"��W��L�tWp+�MD�ϻ�����~`� ف�̍e@�2n@��T# �.�����Y�R�0��
 �F�<�.��Q;���,�IC��_6,
�M��I�M�?ޚ�n?�Iʵ��5�Q��F���NU�CQk�JǠ���R�wR_|ї�i��R��ܤ�z��`���\�
a>���_lA���Nj�O͈�F$��M���wv��#�#V��2���P>���D#f�&O-�Z�����0�U��N]��*m�a�+>���׸�(���Ϩml�芒����F����U�q�{� ��B�"�р3�$�1��˗ԯă[��@zꉴ&$dd�y���]W�4Xa?.^�	-nUE���F����d�@g4g��w\m "�ܬ�dO�'�մq�e�CC,��%z�[���u&Ӷ�n�g�]�]��n��4�֟>�qVm�dƌ����^փ�P��]b���ozN?Z��w�i�Dڴ@q$�n�:�1U;�*�C`�^1xWN�1^G\��Xa�wH�ئ)<$'C�b-��ސ;ݢl䴴/��1 �r�G�=SP����[V,�Y�$���g��D��9˷�<�a(�B�6mzފ�󆌦�?eH���I�B����8:�꠷����j��O��a�M�M�g&ħ��Vd�|j�o��[`Ku �d��7�������C3y��>m��)��G����Qe��#G<��iM�Y���
���aa�F��'�)��n�k�mL���l}�3cM'���W�2j�6�i�X:1���}��V7c�5�R`�Vr����4|�S�q��;d�a"p��p�oδ�;q2�$�Bj2!��=�@"oL����H�.�7�۴�7�ϗ)�vs��M�$��ł.���j����*���C������H�����+�T�7Ғ��0 ] g�q@g�K˥0~�C�(���K<�p�Sg�V����S��mo�[5�8���m� ���L�,y�J����
��1�Z����)��$��^}��5ɳ���S�N��l��?=�L8Z�5�G-d�%���$��}_�\p%xA��lu�9=�=n�f�h}�3u/Ӻ;�}�����Lv��`�P��z���A�[����ˁa��Y����R�MI8_$��#~����[���v��.�_"]��1�V�uQ�Ïć�ހ��BkY��G<�y3�9�J�x�3�f*ߑ�0��/$�b�)�1�(�[�UL�Ke�����2��JX���vt@8�,�P���%�n� _��b�e�B�V�A�;�͟�y�k���6���x��?��~'�&蛽r�����;;`Uf@u,��>Ԫȶ,|ȵ���\K H��)� �ӷs��tA���=&E7}Cp���Etc֢��'��d��I��q� �����3H1n�'N_���?I�ί�$���|T|7��xi�K#�)�j�GＣ$�SA�80���`TD�=y���f)H{�>�1�ޢM�s���1ץ�d�b���~�G6�+�B C�f,�{K�\�37��q�\ל��e�-Q;�E�m�!m$YطR*,���Q ��">gW
�Qz}y�j�Ԓw�R�� D��d���ɞ�H� �B@�e�ZtbE�����X�J.^�{�r�rr>q�c}ˢQ�We�{8!c0���w7*�>�7%ZNJyvJ��Of�����O�-_�h�܍�P�< ��)`�j�!��.�m�~�FZ��>EH��hͻ˶����5�pJ=�ĥE�^x��BA�	B��p���7�f�f�5��W��ZZ8����!��D���G)r�k*9�$r�F�~W��G����s/�i��A�ix����!��FU���|h}H�w T�ц=�,�;�G؜zqB���,d��G]DTʍ�\�,�;Q(�u�_W��2���1��ؔ��m��0�M ;�t[������q��g����H'��AqU�vb?� S>G`v�jkm�F�'�:0k�ǥ7��ݻtw�4�*�Ŋm�"�i�-�j�#;5���F@:�qD8�H=y���)�C4��=�����+y��:3�JN���K��ZG{F(�ٸ����>��Ĩ=m��ó�{h�뾴���j������@���f�$8��{�֑i����'���������>�dN�]}ſ�ߌ�ZEtZ��$���~PS4v�D�����w1�?렼}
#ل�^��uC �J{�.�ҋ�cF����t��=�.��SF��u���1h;J��u� >������Fd�7t��k�c�C�j͸9v2+�>��C?Um��Yī",�k��%1����K��U��&�����5]eͮ�>��$�2�,��.��4 �{��}:GUD>)N�}�V�T��5�`�v���x���))��/<!�l���~_�$8|J<���
��+��4䵘�;ZnK���N9?�t̴\��dh�)7L�[8�5jQ�i@
-R��ռ+eE�������W��QXG(�����{��z��=�X��T'W�|&�^e�sN��?�Ԋ$�e(Q�3�+�M-�:��l�۩�d�>��X� �w�L�H� '/�ʙۡ��OB�i�g�\���)�x摎_���x_#���e�Ǿ�ܓZ��-)���D�wtEC�IH��������tГ��[U��<c�<��H}`��7�T*�� �� ��N�����O#B�	���	m�L���E�p11f�������n�!�׺��M��
[tKe�	eI��#�̚#���aS_�0	Ƨ�lN�>��1	��rX�Ic����}m�gr��	X O�W���1��#M�;��B})�*"�k�x
yE�����.��juQ��#?�dO���IU:�"3enW�n����B��v��X�������]�45��0�5?��{�>�J�I.��� 5b:>���0�@da���ٶ�K�b�w��̾&�H<n���p���a)FPz����U���m~@f%?���.�[�Ƿ_�~ً	ﰙy�p��X�Q,HS����=��T���<R���/��5�#x}X��a������	���o�|D#B^ᰗ����Ni��>Tvo�'T�4<��>J�=g�ڸ�l��t��vU�3)�g��"%����`���"��8�#��a:�Gt�����{g�	kd_9hQw0���
ͤB38�c�C�p�#Ў(��������R�c��C�w�-���v
j P��wi_-���c�.{3c�LH�*��@%��BX<����DQ U �$zjd+x�8��Q�z�x.$���k��.���h�X��97�����5�kh"�8*�݊чP��ʀ��S�W��oKߢ��XJ���h[���W��y�����o|�y�o��}��	
 #Qp�,���ʋ��*2it�d(�8R��_�&��u٨��~�:`	��Q~p	锻o/F{f��.W���qd�&�΀��W�٤��ʼ�r�3�/�C�]�򲑱�Hؤ�M��+q`dsL��	�n��<b��H��y�V��ك����s�+KIs���
�$�i�J�_D��i￬P�s��$��w��?��mT�A+�m�/���H��q��?��?R��$�Ub?����S��5��I�VZS$��X)'�@�v$\v],�ZBLb���_�� �y�a��g�K����? �k,��@�55�]7bi��o%����v�vL����k'�c����o�0�CU«����hQ=���e|A��^��.N���~2ꇚ��),V������c�m�m7�2�x���?P��߼��G��3Q��fp$�K6������A����u�g���t�(06��[a2��5BO1�H'��S��^��ZW��tp?�-b�o�t^���`����1�;�NÂ@787{�ӫ ��3Ը4��eK�I�*X+[F�1����	5`�箪��N���d�0����r�E!w�r�zP�YZ�픈��x�~���ߙ�AYX��ћ���\=P�zEqbZN:i�g�>8�C'^��$�L�h_l7>k�p�~�z��z:�tC��#��A���L��aZ+�2�W�Z������-i���a����Qkk�Dv��p�/ͦtV,����BFo��C}�"P\�� ��ht٪���v<PAul��G����<��Я����'�Z�������`�˄����]�T������N���d�_�A�~cqG� /�)Y��Q4����I��D��+������6\�jQq\AF� �ر�6����ޗΙ���+Z0 쫝2-����0 {�^�eØ�J��6ǘ�z s�A,��*��sz�Pߚ!�����=Z�MW0�c���]���� ��Â\?g}���<�契����n���v�MdX�V<M�R"'�yQ>#�02�8k"��?�(���Z��Y�d�N|��`dL��W	��lFM�_�ϝ2�vy�GvHc���k1����B�����!�9�Z"��2����I2�����l�pu�ހ´�#�����\Ղ��/�R8�[��ܲGD�o��.4�����߀����V˴<���"�4��:��*X|�c���3}��v����/ѸTP��u�U�3u���/D�_]��x�# P�����Q���t'�՛$���O
�b(b,/��)b)�y�a�^��:�w]\mr�B��C����ǿk��y�d��:ːʁ$�,]﷤y?�f�h��Mf���cΕ)�:�wb�4�c:$0���	��G�?pi����Ĵ���W�ە���� �Rў�w^�>�@u[�Y���	�+�������o��C2�!�.����#�L�ldan�q�f1Z:�y�zJT�@��i��]��D�b���~=�I�2I㤨�*��Vja�ޙ�m �9�O����s9jx$m��ʊ�<��<�B�XG�El�����h���ShGB���'���rL����7���Y4��\���4B ��]�3���T�~62I((�O���T�����!��˕Ңͮ��r��=�Tv~�P\�`q`9z�Q���El�Sv�"
�T'���Z��v�n:��y���ߴ�"���Y�1�pH�4i�w��&N� ��:a��h�9���(P$���x�)5r�]�
u�V���v52/�%<T%W����.���Q�������-SV~@O��1{9��	�D���慠��l���"�È,3�j�0'@�0�v��= ~�%�`��Pjp�~] /���'��Q�*pg�Y�̫L�)�y��V6���X��hS�L��z�b����n�@�����. ��밡o�����|_l"0ge?�{����\s#�㷣��kBC{�1�ve@�Q���A/�o�	I�G~���?�% �Α�<��<]�
/�Z�
�{�W0���yO,u4k	���Ry�"�bho�-h{�i	�OF�iM���I 7�]0�.XS����܎�\�%�>in��x�C4@�dt&?+o:z�'�����^yH��l����Ѩ+���*�����D�Y* �N���d����c�b��#�i���P��-jba��c�UqP���,gI�3��P~��K�9I4��[)i�c�D�U��!�8�Bξ�ߑ���{��>UV��06F��`��%�|�z���t^?0���7/^(�t���E��������%���%z�#^p4�g�dlO�
c�,P�eZ*�?�]�u3��w{��~��-ֱ@�E=�6#5�T	�m�0lI��)��)��4p�9���-���ʎ�R��.b���q�&�7�h�j��%� ������ЋW��6�T$hs?�|<^�5m�{�+Xz�;��(ͰY��	IX����wн��6~'��)� 8U.��8ԫ^�a׃ۼTɶB�L\��;�s�� "����5��e{���l$��03vR�~x�_ ��4�Jϥ�܃io��fwħX�t���/���uB�X{|���`|Ɇ�k6���#����/m��?��9�=�)�oU0	���q��E��iO�4�4}�?%ؐi�n������f�쏶�E�Ԭ��>Są�D��i�z��#6�W\꿡�"��DS�U���ۥ��9`��T����_2�~��T��o]a4���[�
�XKFM�K�v�G��\E���j���)"�qQq.�0�����}�*��S�Id�N(O4��ʣ=8Z�.�U�~�����6A�Qy�
�F�d�V|,�Ƌ}�N�!�z�ú�q����Ե��U����;�qL�l��-��E�b+f!��+��Y~U��UK`����&"�m2�N����e�}��keZc�K�p�x[Am���*}�f�� ��%�����ar<r�]&Y��BFD<��2>B�3S���DE�]&Hރw� �Q�U�;����Q<�k��{�+�jv*�$�y�1�J�H��ݕ��t���s#2v8-4ä`�>N՝t����:HO.נ�;�P���PG�6���BۖA�s8*�0/��@�aL����v��Α&�/��A,X'>��1p���>�_�2�0\B8�z�Z�w���<�~�o�:�����`�jL�dL?����^k3��$�J�0�6�k��4���_�����A�D�h���n�)�9E�4��n������`mƀ{.��e� �Op�*�a~���KδKlkV7�9����H�e�&�z�]��A��tV[�}�z���^[�f�FH���eRJ�u���	����K�Q�&� Y�#���	/m���FX��]�Vpِ�:���u�/4m��+L��$f<����Hj����C��A/Z��r��?Yc4�n��z�p�������$��qr>OS0���o '�D�#@�@9�W��6.?��/�[q�l�U"�V�/=����F��7��}�&�ߞ��Z������ޘ�p�ט�O�1́Q�,C<@��b!M�B�;7/���ѬVR�V�H}�VS���h%�.L��=pFx�f��wӽr]���%9��D�b_yW��]�f0�5���ɕ)��������X
.6��̥k��y�3����'���k�Eдg��{0:6��
�{7�b��kȐ�����a+�L���T����T�:{Uo�O+�O2�q��SrT�D�4�9�H�P�z�ff|��B��m���3a�
�Y�H���E��y�������k�r��4I�W���x$�b������&]-���.u&����t�<Mg��wX�]�U5�`�F�˴�`[���T��%�&�\n)�3/*�A����= Ԍ�X�J��lu ����j���Z����+;(�]aP  #qc=V�e��+m�U���|մ+�Ƙ�i�y�]4Lzbc�6>�@�5!Ǽ�#���m��͕����V�d[�7�y������f�1h�n�p�J$�1�j�,�D[�w�$IzP�|%�+2j9G_�����!��;�I��y{�D��4; >�PC,��ǎͽURԖ� \	�C3�Id��s�N��T�/��/勒I��|瞱h`	��20�������s!�Dx����4�o'gF�1�PΦ� �Y�*�lm�x��l3[�oX��X�b�s��c3����p�UMfn	��D�yƻ�p�J���m��� �a�����OX;p
��T�ݥ9uGH����ֈ���.*&�>�8T��/��s_�:0gJ��Q���;���c��������
K'�츼��Rs��9o�`��M��U6	��c�B�!��!%h��++��Z�A��r�.�t�d��F�`r��i��`Q֊n،^���u�7�������K˻����A��
�����{�0�M�Je�N�F �x��=N�7���!ڤ�Zv��0�0v�#,�ԯL���x��_��e�;��;Y�Z	D�h����E�e���q�<!n �ޝ��h�ʵ���Bu���"W�˽�zp.��c�9�{��5:��x�5���{9tI�2��/�]�a6���8����U<���~�#��QaT�Ҋ+�t�;t��7��A�R�[�tg��:���N� ����3.H�6�g��*�Z<���*z��?��?uQ#��t���d���*�m"ԭ�>o=��y�!Ǳ�G
z�B�����|+�3[�HK"������{Gh�vߙ����.*��. )��+��b%�ȂL���;o�%X4������c"�B��i��h3z�J�&�!ɸ�E���EY6-�Ԟ�M#C[5����?L�83���3� �h8Y�5{�I�C�7
�Ț��p���ƕ�KI6��Ζ.I�1���Yq-<�j��g���%��7hc,�&jwp��lFׅ�\��*\�C0_��#�kFG��=�y�v����v:܄�p6E5T�cɌ��\Q�R3x��Xڶ(�${��η��̂�����(8i�=t*��K[�E�6�V
n��=	��+!r��n.0W۾R�0u�F ܱ���{c*ؤ�0/@b�+�R��*/�}g�y߳M���I�m�K���k\�p��;w3v��3����*��1/7�yb�u��._rK1�&_]IQau�gr3/����$9Z�V���P����ьU?��皏e����d�� �����Z1gf<�b����!�_��������}��BBL�?��X��d�VOK��.^����ln��yBZ[�\����?�E�n/��bg��ޒT?��Z�k[���E�G�<���)��IY<P�ұ��+���l�4>��=A�P��ow�~� >i�G��e��}l�"��S�TjU@����� e1(�%�jN�OتX>6<�;V�d?P�TD����4=T�٭��6�I��9H�i�oHF�׌���$K����P����08�I