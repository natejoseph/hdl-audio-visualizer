��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����;* �{pBԢ�Y[w�S�Έ���+U����������{���Pqm�y$�T>H܎}$��6,�W;}{(��CTZfW�|�[:X��QC��L`�t�b�$�.^���a�*�۪������Lș?���s����MT �y 2c
dhZ�̀ʛ�L��(����G �l�������0�@�;�X���Ɗ ݵGD Ɓc�"��5(���3ǫ��Zʃ���;U�h�U60��e�q�a��Z����G�g�TH~���w͘!E;�.�Z*!e��:
�c@���rE�o`~bzGa���v���\�e�60R�b���p�*� r\p�¬r���
`���ӽp$��sVZ��Dn�'�H��2������uR8�o�T�1;5?�c�e_J��-�x�R��D����3�o�����d�]�A����LD-�'r PO���5���j��`�q+o�W)ա�n����W��(�db��yPw��Po(E_�<9�ܚ�7��r��l h�fvĦݸ,�����$�{�*~j��̦�vr�C����������f���$��AB�rM����,�� ��u=�g\n�H�%�*�5ydNEhc[o�#���Dk9t@��Y�'i�r0��J�7�� �>F�d��Gw���pփ�V���{�ɧ�cc�!v�����"-\p�\g��ǎ���]aE�3��>Z ��M~�GX̏I��W�:h��7LtI�M�%S��=\i��L�w}��&c�I����k̜(�#�L�"�o-��ˇ	���;�g��2�G"�g�v�ɂAe�*id����F`��k�w��-E��5z֕?��FPG���^�+HP)�q�eyΧ\v��\��a�?�M}&��Y@.ZI~��hQ�'Et?l�[�:�؁�@m0���#��n��Mى�L�g��o�+#�o�c��:W���1�~T>Л�N��)B��.�oxj+n�03��li�NW��`����#�2��-�3M���v������'eQO���%)�B�AIp5����}꧴gLk|��7�ցk��\���M�}�U����SI(�A�7�$�D�=)v����
g�@�39�ea��aYK֔R�ԁ�-Q1�#n
�8J���un6t�&����{=���l.��y�l��}�*L$G���i���}��M�2<SPs�t�'��Mvao>e�����' �zH���1�o�A����9�ϵ��0Q%��ɍk=�6L��'��k}�Ze�WOX�4�1c8K���D۱ 8d �s9��L_cCX��ి�@/z,�;+ ��ҁ�R�y�=�M�̃w1ù�'x7?�����dT]b�-P4��
�I>���G`�X�ͧV���d!G�
�崊�2r��Fe^�������Һ�x�Ac���,B 	B�����1��0g7 6�T��G��ʤMUf���(���Q�^�m;.���*c?��S������@��Z��������u�B���!R�	qt҉%κ�Ζ�����I��G8�����E���Y's���Y�qpo�QQ��6���,C,���
{d��+�m�������I	�-��x���YT�X��$�҆�~����߹����lw�7d�꜕P.�)������y�FU���$P�[A+�zO�?��ʫ��'�ڎ�B��G�1G�/f����FeM JfM�
�>P�!��}}�V���H�F��tBMvQ�G<A�p��(V`��&�,�`n�4�����W�_E�2��R�2�
&S<ܿUwˊf;���F�mA�q]�U8�S��G�>8���?�6zkڇ��A�J�r�khRφ��aϜȣc��Q8�v����������.�K�ބ Sdt���(=ը�g��z?	��������������W m]�`�I�+G�[^�:sU��f��=��w��Y���B�Nm�c����*�h�bk�!`<��ջ�n��+1�y1F5kr�e!��{��m'�9[^Um�d֘�l�}E�3�)D|zd���,.t%�1�g��D�x`�ϛ���,����*Ce���b��t(�H���©7����f6|�<�D����y�s�%� -i�~L'q�x�Z~�����rE�a��)�dHŶ�簷�����>%��A���d�v�NTwl��0Y�#���ǋy���6-C����ݺ/���b|"��"l���lW�Ze/�k�d�&�ײ�M ��"�*7�f&�^���g��W�^S�CY?����0���<-�0r��������sO��:��ݑǛ"�K֎�wݮOQZ��0�9r%@pF?hB^�6l��c癓ی�j�I?�H�[�}���eN6�]T���/�.R,�=��6L���۴ĝ\�ѯ�y�P@O y�b�!�X>%N�bx��ǫ�u���b�B�������S���/j�e}|"a���D�j�!�\�K�Za�����W�s(}�7�F��śq�n4�|����A�'�����7�$�od���f(`���<�}�� ���X�B�b,��D>o�Q�k9�c��#���H�s��v��O���L�>�w�&�\[M��8=(�P*,Ή3���{8(�$��A��OI��s���gq�`{�ti&�j���~Eu���Ur���:��2�Uc ��z�M�	��:��H�_^�����(����tTD�}z�{6���V�|��vt�x�^}͉H㝕�ǒ\1'�}u&�1�%p<E�|��q��%]����w�&��_X>�IY���@��|��������oN������k;��C�qpT2��Y�u�:��90⥹B#�3�ϧ�g�8ָ�!a�>��Ϯ:AJ��^�iP$����������g��$���i��Nq2J	�,�� �D?.�����v�*���wp;`p��$�d���~	��#����(��]D��o1�	�e&��Q��?�]vw.���Д�~�|̧͓��Ye�aQ��d=���<3�~X��&���v�k�f��k;��IhI>�c�2U�.={�p���<:����u)��`�y���q
)��CNf����N�O�
�����R������8-f�*�(ke9�
��.ҭ���=������:�c�4���k�;�@J�{x�nMW�������65D�9��	%�M[����Y�k�c�[��o���cDI�t�TEM����@<R���Z��v)r�9!�a�@}��0�جs�����(�h����82��a/�K�$ӔtN���n\�ݹ�d��x��2cH��&-��s�I�X���H��w+������_�P��@�Cen����as!ض��J��[�Cg]h>IX�ŜT����V��i٤��M/���Ƃ��#c|��o�����Ak�m��L�j�Qt2��^��������v���,g���()�W>�,��}F�,E���o0��	iV�"I�2���q��䲪d���V�W�ԥ��8<"�C�r�47T�qt��TsC�v�]M֋��ȜK� \��e�n_���<�����j�{�W7?,���P�������:k'r]��� �%DE�������CU!�6���fb�%k�>/��C%Um��d��l����O~�N(5Q�8E�I�M�Š�o9J�\n{�4&�J-��#�S;����RϨk$�/���/����"� Fb���t���IP6<
I��nqTG��E�Q�yggu���>�ʨ�fFy�x�����xvv�_��[;�&W#��S�C��*6��dE���x�ڻ�g_dC��vXs��Ll�\�<�K�Y{�P��P �t��������HǦ0PH[�_�j�0��2�8`��	�z_;0�^��[��}ܳٳ)���\= E�1�ծ�vg�U|o�4�l؀��}��Z�#�.�h��խ�Z�*��E	�bG����>0n��x�j�F|P^nF7$�g���yJ��G?��ɺ�&�����I�������Ⱥ�:�2�y�3?f�١:���&Ř�X� /G0&w�J�
���y��}*�-0/�����
Ժ�G�|U)'���>+K��1i�"u~�� ��Ȁx��ᑝ��V.D#J��-��d�֮��T����Q`��ͦ�v#i����?،���E��Ѹ��9D+s^$���z�E �2&g�11��L�8����˄��=u%�Ǩ�.Hl47t�V#LU��{�w&���R���dsl96/N����uߵ�4'v��a�wל5���y5b�]��ʬuO��ͬ*�SR������k�����Y�\Vê'�#��n������(b�j9��r�K6{ ��R'��~c��I�1�2�*R��k�)϶�BBʪ�<eu��T� Ƈ
)M���~���'"�Ob{l��j���C����5�t�4��m%�[��zJ�h�j3�`��R{<��URL��bY �5�;H��Pj����;�˛<B���@���է�U@'a"��b��%̅�K�/�P������RfL�JB:	 ���ٿ�g�����g��W�Ӌ�b4V����'���AV�s�G���Q1�:ƣ+P�eXHW>� ,�N���g�"$�w���$���\���0R�������3�@��s0np��������;Ϸ�;���Ȁo�tY�r�B
א
�.us8�r�{�u#�7�C�ς�+�,H�lb�BV������ڔ�{��)��w}�al���`�9L�u��W���u�ȱJ�%[�	p p,/��S2p�[�Qy8^ͦ_���$�2�X�t)����BiLmZ�O�VZ��" ��SM��*ٵłN�<�\yүgCx�IG��<�\�����K�+�xfIW�*n~�0`N�2��E	S���	d�U�wD�֪p� �;�Nqs!0�>��8�
��\�I��(�d�Ӟ���  '<���%��VZ�*� ޜ��T%�"_[�6�x�\�Y��E�
�N�[�h_�+�K�!J�3�b���BC5�\�Ъ�
'���l��f��*��1�+V�EeL����_w&~]�������#��:�z���	b�m�4-yι�\jQvt%�j L�/��.o�nV�z�Un���U�YsӌyM�^@u���������Sz�ؖ}���a�*�F���!����:8�NR�A�d� ���?���ڎ^o�!��dݢ{�~xJ7��w�yCJ+��m؊��`]�.�8N�%���ֽw�5u�C�cg:����׀&�6n��iGq��tJ��<P@�=9\�`%���!J�	����%��"k���R�����|�刜�	r|��慺�"�H�`��d���Eef� za�Gs1��}�ǋ��[�?��09�xڛ[
�{�d��:����9�ڵ�w%�+ _$�]X�d,����T��}��ϥkw��S�_f 醄һ�"#o*���}%�f����Sh)���	������i7�@oDj��� �4vL2��N����2�4S��3�]"�"?!�Տ�S�d}�`�G:$>Lؑ�ʳ�x���y�����4O�������*++Wa4�o�OhQ��刊�h�#ub*�x�����Wyu�	��/�$��gi\�9���5�yԾ���@��s���?�:Dzc ø�+(�����`���!՞TY��#K��N9��"�����>���L�MX���)�C�_r�.D�v	�{tq��0��:�H��rЈR�����Q}�ɟ�S�sPd�8Y����*=p��W\�2�%�4؏AB�������:[(C]4�J��QJ/��e!�������[�팕:9�������~	���Jn]c��E��&����Ev�o)Id���`C�^q�,n�M�%b�F��o<rbgg�5daH<*|�����g�tާ_��C���j��)��c��@��B��bͽ{��RbNM����R�z#z�~���fUn/���q{��nG�<�d����)yw<5��ט�*t��oYA|}�B�G���	�0K=S��D�Y~�b�SV��R�tz�p�;��\羕3����PȹV���l`#�aEf ��#:Ԫ�����F�老��"	�"Ʀ�4o���i!�61�b�C
��$q�\J��U�A0,:{��\�7�▀Fج�6��*���tI�i��*�'��\�rt�Ռ����k@���:�!�?�"�P��k2�L��.j�eoP�D}�s�w[��D5}b��Жb���Z�z���R�ТaP�S�@�|(3�^�^@�Х1~:�Ȇhqp���. �{F�bw,�t�b�UL�u,��]W���x�Q�,�����a��-�L+ZxT��`h�;�Ԩq�k��=�j����Ǌj��ѧ4SHc���Т��B���_�p4�
|;�-����$,����ӌ�B٧�Ȓ�Y��ϙ�rB � ���ߦt�"�s[^���H��/J����E�E�TqãY���>�����;�MK6� �l[`�x0��Tj9/��ձ �9b�AH8�*-\�{��H���܊=�Q�(�0���,*��f\��%�<m���)D�/�����h_a��¡|�d�SL��H��_2G}ey;K���æ >���la�+eqCدYbQ��=�Zb̨.�8������S3�Η�k�;M��FVȿ�X��ba&�i�E&dy����L��:�$�Y�s>&�Jd�����e�s��7�sZִ473��ϐ��^�' ��}¦0W�e��f�`� ����]q�����:�Z�"ks��Q��︂3����/�:\"8��p	�0��z�iR��+O7��{\��aUloTq^�S�>�nᕏs�y.��-Ž�D�ŋ�f�Y��~J���ߺ-�\��4�ș+��hj���x�ᬤ�:[�v_���e�sV����
��s��> 78rR��e�p!���8Ff�h�7�7ү���"����}Ӓ3�
~a��?�[� ��V��-��:�!�o7=kI�h���p�~��G�w���lgh�МQA�$+Eh���r%E��I�ٮ�=;@	�C�#���c�q��:~o�}�����ʮ�@�lNdg�6D�Z=*U�BƗ�|�����%�A"����i,�q�Ky��b�����RC�レ/���&K4��߶�ŝ~rB�v�������5㮄ׁV��.��:�Y�ba�W&h|f��c��"��Tn���z�~� y�;�&0�ʱ�� zo��ʝ��r��aK����P�IX7V{�
���&�qNR]���r8y�U��J����1�@�>�Uu6�/��3�.�"����HX,l���p�s�U��kF<0��}�?�Uv9�X��z�1�ř����+?���bu�=킢��G}��eRb��������n��e��5y�'�e9�UG�[��)�1w�r9+�y����<2��b_���S�b��^U�4v=�� ^`E7�8uP�#��K��.׭Q{'�w���.M�6�ٻ�H���]����c�+�Fo�rQ���)�q��0�㠲9J}n���RqD+>�d�W�����:Mc���v���i�z��Q�e��X7 ��	P�}-�� � �@�{������&�B,�Ayxt�˪K�lX���C���)��V��)����kG� ��];,"�&�iԴ��n ��7L��0~��uX1��r�=��@��~+�I�vg�:r %���\<���?.ɭ�Gh�����3σo2�CH:�*�w+�G��_�t#s���9`��$~RA�A���<�p����9�"�Ƚ��쫑0�K7�r������03�	�M�su:/�S�����miрk����8�3�����Z�r��;������P�2^����CX �6�:���j�w�|Q��3��:�Rp�u�!��,�ƺ�&��/��92��I����`�S��p�TնG�#���v�^`�Y:LȺ�>6�B��<ǝj#��%){	N2p�*�{��71QiQ8A&��r����zu�k�:�+=��"�޷��g4�}}�ֶx3[K�-�/���l��"IU���=���a�@�p�M?��U����#�9�}d�C�_�N�9�/�$�mƑ=������:g�^��,��c��m�
�X2�eSb(�m��eE��z'1\&��D;��9<t�ZjSs���_��S��ν����c�S�s��}s�<��jj��G^_mf�T`�Ёn�9AI*��ނ��ϳ(L�E�N$N������O�c�I��TҭE�<����ɗ�]���j��L�V^M�lܓ�8�0W>u�q&�.& /���� �D�����H;V��n��� ��Fg_E�%�&$�e��
Yl��M�E<��iЏ\��9dZq��,�g��4��~�*��{�׼y���E<�!��5�|z|���.c�\{��#�R�|op��d��u�vt�a^���)�%v�rdfl�y�q���v��0�O>V��
���p�[+\Ȋ�$�����;tr@�&n�\~Gv�onl=�975z�z�v��d�	#���aǏ�l3f�$!��oI�pr�"�w���ĕO�䨸�c�Z���9-��FZRK=-w��3譫��G�wa�	���L A�����5AUTA��c���� '�����H�
&�7�/ƿ��rt�s9�ӽR/�'[�W)�Q�hϰ�!&�W�LKʼ�@���Q��l��1���hGPeXz�"��B��$A�+|=:�,q��>+���N�բ{������DW~���Lّx0^�ٲ"�f�F :��ֈkʋ�H��H�J�.&��}M�{&E�a��e�+�ä��\��f�q�߂�2�qzgi����f�͈E��j2X/�I~��s1a�PvȡxI[���.nX�/�F#��&7U��es�T	�<�\Lh��Ԅ&�q���Q��C2��pޏ��]A�1܂�4��qNA��P�r����`�:&+����=���S}��!�쿂�<穽�<��")�Y�޳��S7E��iɉ���2�_j��{{^9�U�a��\�O(�� p+W0&�('����iA1R���EֻP��ϳ|���G`j�8wc_��ߝ�tx��d)�TF�GI(�& �m��QET�]��q���Ed�U��h��tх�	���U��|	�Ύ�-<
���L�:�K�L�/�~v�b�G'���b���aK���ǟ����2ؖ�`������݋;u�y����B���5V�Ǵz���e�d^=J$�k�gU3țܝ�-�8�dt�FC9l�n��9m���Kw��~W-�9��o��>���d6ݮ���@�g`��rMg{d���L�}Ҳ�3}��&�v���Z���#�\\Z�?T13��L��U��U%��c�0��jޚg}:�w`�p�K����%"+yvt)"M4m��+�P�j�ac,�}&DP爼����;GА�ؐ�3��w�^��C�1>,�=���@c�=.��h�5��d�ڹ�RR0�gV��I�Mv}.ƫ�hi�3U^%�K�"���@�@����+�1����"�V��_1���o�G�M�5�I�3�J&5��5��7\k�i=�ħ6��Ӓʽ��9_�	�\r��I;�>�d|�w�%���'l-�7i��3xݓ�����`~�V��&��,��{Y�|�
���R�S�����O�ϕ�{�f��ME>�r�2����n?���b�VI����gz;�`ߍ��P�p�����~��Z,��іvۜp�H�>��	F@wY�m&{��@G�)����r0~��/�5h]�uܩM^Z�Lo�J=`���V��<@4zJ37-x�¢H�*���gdu+����#�߭ܣl8S�����<�M���/ח��@|O��1��a�	6�y��if�}G��7�k�m*�S%>�ؤ���C2r��F<}{�({T<a5�!�	��T���C8��NdE���O�:����'r&�֭p/�Y��!r�ʾ����t��]�N��87���^�_5�jfHrSV���@���S��K\~u�5��czo�6[�B����E�Y���Z�N�t[��	s�)kwz4Gj	���d�m�G���M}�
�DZ+Z���$�e�iE:�ISDk3ى�:ق�Q��.M�պ��s�$��0���f.���:�*DrO��h�+lw㭝�MH�� ��jC���xxPn�u7�E�M�SP���%k�  +��0
w1�tѦ��/�[���U�
5�B�h����Ԋo�>�[̒��Cd���g���	+NN�	��΃H�c��7:-�W�l݉�g�[έC	�Z[ [���X��8eJч�����N���@�.���Q�:@����r�|Ao�ɿ̍m�sQ,aY�KH��&��PUԊ�!�
�������bm>�6���Z�ǋ�����s�G��f<M x���5�-��>Ts��w!Ո®�N�uo�3��<���-X��1�lB�`�DQ0�8"xT�U��3>&v�Xq�Î�4Zr�D����x];���
�q���I�E���c��|���p�m�H�*��S�f	���pZn=L�Q�l�|	�8�o���"vՃ�GS?4�7Q!����o�`l���w,��uSN<yj����A���3t�o)��kNY�2u��8 �o��kEi�6�-�#��S'���$���L��]L���ti����W�Ms)ѸW!68qr����˺i�}͇	��4'���)%�
m�lRn�=�2+o���a��\��:zٴ��K@6L)���t�)�&,��!ߵT���$%���z����+��N���[�j!6�:3�c�m*&%�i�$ϊǏ9���#w������˦:�I�3��+_N�~�c#���S$%]����\�`H�`��{ <���VcC�{�j�o���K��B��+��r�ԃ���M��o(��5g}eV��ArK����H߽O���^��@u�ݼiy7}�	�A��~��Y3*�&��ӌ067Ѝ�I�����ħ
�t@�p��ҋg(gHh�9K(#�/�^*<���'����A�m�&��Yׇ �mԮU��䫌C�	l��|Е�)��Q�'�e��UA� �>jr9����5.��z�y
A�+��F\!z(�jp�s�o/7s�����c�����V�%g'>�w}�MU��6I0�Rj#9>W��kr�x�^���6�I')�U���"�D�
	% ��<�*�3�t�pF=�ꁆz������(��P_uf�u��a�! ����q��!jV����!�Pm��:��漩����zi���w�԰7p>E�S��O�zmA�V�����m��t<1�±�1OO�F����d�|lK�ϵR\�BZZ��}7�r�Y�Í�]���}�����t�.xS������M�M`?�t���I\�n��u��qVi9		Y�)��Lcv<bT�t(|~�~ߘ&'C�����TuU�����N
�PPXn�n��,.�ˁ3�0�`V3�@i\���\��ɻy<xCJ�� e����@�tM��N+٩|���=r�<��Y;zy��Do�Ajuu�`�3%�.�"2[��*���t�s�j��o^�z�;�O��²TFU���e�`���I+��չ�L"�xH�W��Z�M0FAk�D@�����=�i���ڲ���J3�^
R\he*�g̩V���	�֙�6�
���iW�q��\5Z�������B�r��Z���.x_��9c���	`n'�m���1��ݛ�D�7�2�7��^��)��w��ŘR��4mcN���W�K{H6l�*�L�]�g�%����"jrߧ�0�F�^��dt�� u�B�-{��m�c�<�k�)}GҀWHɔa��K�7�$٭U�3��cG�
G�Y�7�Qs�LY�kw�̊�G�0���9xH��-
����Z<�g�A��7�ڛ>4�E�wˏV����/-
)��ـ4��&L1�Bc-l#͠�\3I4*�W�?��M��^Aֲ������%s��G���JgR��������a��,y{iz�x��bĝʅ���Ig?gL��2�ˑ�����zQ�Gݫ� nk'pvY{��ܨ�24:���� �6Ɲ�W���nU����?���}`}��f�������́�È��	�!�k��!��T˜�7߬�2a �2�]���4{c�ȃ"KH���ag4�x�[ы���yk(-�rL� �n�d1���UXQ���jR�}M�a��3���db~T�E��z�X�֨G���U�K��R�M���ju��2�G ��ef5��\1���%�JRA:�����008!������"Lޙ�<�j�I�@Q���H��@{�A�3�S�A�t��=�{����˺8�h�!�Qb��Z���Xƥ�A
�z ���|�R����)q2m��F'!�-��%6��%�1�$�����zQ콹�<�/���53_ǆ���㊍����P�����̈́�M����#Vv��ouɉI3�����U��IN<816�R��j�x��N�����0�ew���9*��P1��xԃ�X,r����1=�:I��-Zs����".�ʃ��r�o_W�ʴ���v|�8�͇3�6S�0�=@�yDw���s���nO���g��N��)]����ӯg�/1�_r�������yA̻X�e�*�������ɟ���z&;�մ��w�ZkG�P�H̬��f1 ��G�ȏ�m�d�r]�㧋v&�n��������0�+�
L�&"��%�Wgl%�n��	 8Q>f�#P���@�&��|����dN���?����&5�'l:�F�˕�l��M=�_Gk�C�l@��1�2eyYbV�D��19��}�?��TC�1ķ4	�V㹍�5�Z��7%c���Ψ=�Y��7Β�]]�p�ɉ�FQ����)� �'���yO�o�l�qK.��y�V�ڸ�Ȼ�ޱ{WY��[�5l�Y)D;��zըC�!/�s��J������wȞߝ�dTT
���8��ѼB[@�a��ڮ�6�_eA���S�hӫz����-�	�k��ˆ{z�i���d�$s7a���)d��R�!ҧ��ϋ��=
F�V4m��R�z����#�l����m�B_4¹�D�!h<����rS<��nAbAXw�11I�4�A���A"�Eoӧ�xG?�z��/-���������U�e٭@���q�|Vd��Ļ�����Oٲ���eM��czq���B~���q�������2k[��gJ����".�������$��m���T��h١�Քq��J��� ���D���C{�F]\��K�!�G�1��g%g"�Ai�������G�Jy3�v�2|������C���B�I�&����-�T9}.\v��C�9�t�˾����*L��rn<@9���5hRr���c�<��ijc����C]������M5]�$Uw�Y� X,4$��Yo��v|x1g����z�&�F�Z���iNB�(���C�(R���j�b��[9NZ8�&5(!��n��9剃	jfU��d�Z@V��ݼ�^y~��fF�r�f�����4nF	N��N�.�Y�ـ�tʷ���m�g%�^>�73���e��|VM@؝�y��kM�}������>	��`{��� |�+�z�#� �z28$�9��`�EaQ���(Y9b6��O^�:�QNn��Z[���d`�y'�8�>�|
���}���[;?�q���}U�4�TT�ȩ�X��,�w�nB"	�4��_Й��`O�6I�v(o��\�B
����f�Hr ��8������Q`\z�#��pc�2�v�y����h�/�ҼBY
�ɨE?������N#8�
���\ݜ&4�'6��i������u��Y�]-���:����j�[m�&� ���ј��g�� ^&}��&$A�1DҷxҝZν�P�w<P9܌尚�ᬩً��,��&�t��]ej�%X��{~ k׹T��4�Tr&�Bw�����<�� N��VN���K�Dϝ!�N7������Uȡ(�30�+�S��P]��x~K4��f�R�,�9
�_HT��4wj"8�����`�ב�A���H+ �mO��#t3�5�����O��*�2���r�C#h;�)j��^�����*���<ٚ<=ū��J~��b�Q����V����4}� U#��p��G?��r��>��0��d)�C��?�5����#��#��@�oH�V٤�<��*� �:CG�mD()���K_���5���9j�~yQ>�ƉD?����:k�	Z����$*⩨��L�`�B�s��$m1	$�
H� D0˫�"A+�<Cg�^D;�,�F.��tOj�a�n	������5	��Ő&�#xIJ�
�s��8,O^�{�Ҙ)ՋR�{ڼ��C�ny$A��8yq�eY�����`n� >�q��#0̗�_�f�VS����R`G�W>4���:�!�⿵�!:N^��Az@�C��Ҷ���`�u=@�Q�[�P$�c^�@]*����j��JQ%��ĩ|3=��H�-);��u"�{W��9��(�t���E���=y�w�������5�3�(�ة�+�>���F*��9��L>���T4T%,<���)��yf�M`	�WF<2���QVhY���4�g��!ş�%���v��',�����HRKQ03A��, �e�U2z��v)��cK"� 
7E{&�.@�.F�ek[�h�|���X�zd ��Љ�+�u�ì������ o�U�xO]�o�huuY���M�P^h����+ �wz�[R�p�s�蓔�:y#�)�H����F�_)#�Vv�dC��du۲(��V���;����H�s �[���[Q�$ś����D�����`>�F�Q�)4�����`�~���%�N���Ќ%�z�~>Rr�e<o�'�����g��8]Rjۘ�;��m���U���@B�h�L	�BD#��]�4�(��3Dc6��}�%kޱ�2�ҖQ�es#a���ZL:�N����*�1/�Ǹ�(|�M����_�Nh�-9�<���rK|��􄈇�4J�L[��z���t�L!|�Ȅ<87]��=��Y��)�A�;�����1p�C�6����i/"�IH>d��:��T�d�cM+q�_�k��f������.F1Fk�9��q�����I�'���-vV��M���2�S��ð	��y�����Tih��;�^D�i.Y���O���wM�q��tz�x���>�ˇ�����p�h=����fr�
]ٴ@�9���g�\:# ���UU�r���\Y����(��!�@]؟]kf��iUt����Gp^��,x�>1�l]?Ǉ�5#�[��w��v�jY���3�C���2+�.ϙb?0�N�`�@���Ȟ}�g@����@��m�^<A(/k��yZV�����L����y�O#�F�[r7ZU�Rι���z���D1�ْ�МI���u�>�28i_�ֻp?^Tﵮ|�O�k�&���d�SμL�Ӣb��4�����t��U5�w]�+�r,�mČj%�k�2?J�!���Z�2j>#ܬ4��PY<(�>�Q'��
%���L���tS�u�-j��h&��V�k1�GNZ��b�B%-W��R
��F�"�Ҁ�s��K6Jy���^z�<���K���,H�X��n�Gsk\�},N�C����ٽ:���kB��������8����|߸�$jq��L?f�oV�x��Lc������ qp�5�4n��5I��27*�b��\��^'bwL������ײH? ���#P�D�߶��:�I��A�W<u-n{�WJ��2��_Ĺ�kd�y"�/s�F���2�k���u��NO�}pc�Ę}�6T5^�@�_^�N61Ot�贒~��h<C����g �X{|	��'���Rq����G6w��[��-����!W.��7n[�`��:qn�{�=}�%�oh�ܦ�e�ǲ�����Wm���_����iR����&����$G8W@�D}A'�b-�7����=��[gq*_77#H�`�GS��]�1f�$�6;mb��{�0h/�.�y+zy��o��!�N�����34�P��J��_�c�_�T`_	Y/p�\)Q[�L	���C���+��ՠ�ҝ�ZW&Gw�J��0F�L��^8++���n��A�_����� qy$�ܡPؖ�PɻL��E6+�������i	JZ*���'����qa�rwYب�U�ԟ���N֝7��@�O�>~*����}�p�.��R� �S�R5�F<��n��!]0�W�Er�Nj�lǼ��!������)�L�3������o��~/�`�^#��п��n�{�Vf��
���>ہly�Қ�8`��q {�`���W���Z��k�; �HˈJg�a��\l��,����p]4z���������2��,n����hi-%���"u��5����Iw-�G]�L�4�k��aGM�<�K5���u�A��\��a{�n����b%������m�6�#L���O�����lH�J�m�}"w�����7Z_�PQBLʩ���F�]�0=����_�}r��}��n�P�U�c9 !\����l��1P`����=�$Z������x��e����z�j�[�	�_��Zm��;�\�w����|5�����.��
,����R�{���{�d�H�:W��#��ɏv�kA��:��߿} !�'���4u��]�[�(&F��K>�4&�`)�m�1Gq�M�Q���CW^��x�ܻ������A���TH�D8��}�U���L�mE]$B�����1��`�9�x�cv&w[Z�w�
E�F�V}b�hq|W�O��ܜ'�E=��� ѽ\��ݛ�(��Q(�/VZ���~�˂d��$�:�DM�!r��^����k@I�ag
�#��}I�V�M�j��c|O�����V�%�K�z�Y�yX14LGS��C�b��F9s�k�Ni���(�}L�=�D�Z��M�P@�sT���������h�=�A���A+���e�|B�kțM��7�z|�3ť�����&̈́��x�0���s����MB�?1(<q��;*���x��C�a�]�>7Lv�k4�� M�����ě���� �\�yh����x'�gb�G<	H�
���@�F�c��h�[��)���H����q҉ء���"�C;JNސCߧ_�rW����1� ���͆1�8����F^�N���_�;F�.q{[�ypA��:��-O�*��愅��0����8��[>��#��qz�d (
�M��=����D�Ţ��Ȃ���W�-�!͙$g���J_S��y�C���Ry??�V�"��;�٬�):��1��5�Hwe)�J�����~MJp��1d���5tc�m����M�7Y��Jq��8�Y���}(��� ��:�f�Q;����X?R�vg���n��C�P��@�`]t���ۊ{A��l�YL���NŬbh�&��]�Z-�M���TeAm�n�XζԜ:�|��K�
��@�Cd.�]Pw���p]8�I�	%��i�nN)�U�% G_���O�� ;)�p,�*Sާ�-h(��9!�$ٹLܻ�9�f�MO���_^��c�j!�.�'��S��M���yYx��씡�u>�p���(4�޾��q9G�UV��u#�W�Y���	��ݯ��D�#�C��Me��"fW0�΀0I愄�jd�T�暛]���}��=�#�~���{�9Ar`���L�rLO:g��M�(9w�)�I��}����Oz �W���[��>_t�|@�@};��d?�\���ߤci�H��J��(z(��-�����9o|݌��u�ݤyaCw1�f.{[��@tdxp.�?�`������oG/�O)�ea��:T�FͿ���o}� �՟�.��^�b����)����ԭ��>WCo�o�����w���H8�ЧJ�#�H�]�ɍ.k�Y&?�+β���N�c�+����,��dv'�2�w��>��8B��.��p`�aD��M	��H�b�T��d %��N�o�f�(�u��N�!$��g{�YJ�	Bm;G~��ں`n��6��~u��(b7.�t@}�L�t�kF��ۛ�iA�)xꄀ���i�Ö[v�� ��T�<MϹ(0� ����n���y�ƪ(�jo�r�֨��!�!����aDLN����][�-�X�����r�W
q2�|��T��3L`Oj�n�D$U���&��C�K��j/^2e�s]�?�ЃǏ?؏�1�x����rx�9������ܟ�]H�;,U��V�ڍ>y��G��v��,�UmC2�2K���xis��d��jF�L\M�Z�N��}q�/����o1�H;?#�K@�~hɯ�8�q1 ��!�Gp��#���4��s�v!�X�r�u�)m�sz��̸��D+�v�y�e�p}��ڂU<}�93�gJX�g��
�jT-�k�<��V�,��+��iF�&c�y/��_bqa���zy��s���å0|jc�+G���>�6�&�u6� �p8Pfm��OpI��7�ۍJ�G�._�����Bh|[G�P�A�	X=(�X��-�$����1�'9Gl\���0�p��O�+������{~g���{� v�dʞ �0�s2>=�դ����h�����5�xQ�W>vO[�0�H,eWƘ�cҚ>oҿ�&)��K���5V���lJ�2/gLc��)X���ΔL��^�Nb9lI:N�����=I��U������@k�qP��4��_ oL):��q�_���b���~��/C�kL���M��S�=L?���.=\uW��B����3�U�=V�J����\b�&���4D��uQ���Z��l���pEs9�բ�3��(4O%(b=�!qnȬ��>�(���''������,&z�F'֜G}�3�F�|�'��C�܏�Pb0g�Vj�?h �5��7�p#F�I�����2�k��҅
+˄�km���gp��KB����c�Dj������mˎ��+���p8!A��:� f�n	�|�Z��x�p8�h7���X���b�d4�W��O����c�A�y���1�츚]$�";��0�)���f��?LLTd��Bl�oYh��;�Ɋ��]��J)��*�״?�����8pt��L]�>'%W>������*�� m������Ƙ;���Y�T�?Y�cH�G��*�,�Vv��}=��"F�Ot���X�y������@jYXֹ� �4e$>�7��g��9ȕ2�I� w�o��/�i�o�)�����Y/@�7��p�_���m��s~JK�T��a�ѣn
|��fa��$3Z����nx9ꐴ��_�W�����Ty�[i���둗�+���,��"[,�Dǹ��SU�ڪ�z;�G��"�����)�\RD��=}���!~�����ѣ�������{Y|�d�����xf�(ߩ�����K 7ui@�n:�R�<w$�-ﾐ�WF�u| �� �ɟ�bkAÛ��H����R1Ů8�o�f�}�mFg.���}��9�!k�!<�d�@�ݺ:�A������U����O�2Sq�Zto�'V��	a���Q'�r�P:�H�1��3�
D��4��cA��x�Md�Y[D����J����+�׵���'��H8^�j�cz&ﭗ��B�j)�@-U#��������Q���;��嶩�-J���{��4h]�����ivҊ��K5�u�9�sL��z3+@���邇�Ɖ��t^V�I�k��Rj���N ?�om�])��*���pqP��`%�ꖧ���	��	r�W�ӭd)鏔�Nt2\5Ɉ=����O��_B U�/�L��9�W�q�� r����ԈQ�A��Z�3t$��J�6����|��zW>���fGW�����U��Y�e�f�i�
�v�
��~�l�'to'�jTQ��lCOugFb���C-
b����ь�!(5H0xg��:�c��]��8O[�G.�~~�yӖҳ'
��[
�0'�O�BZ�N��r٘뼕�Y�N������iU������:r�LbuP%��1Z�+��clA�)���m��b�A^���3���i� 2��[W5\7P�Y����?������y����7sQ�.*F� �pCa+`� �o���L�?����zt�fw~�O�p�U�Itz�Y�l�)^��A%������.`���T����-Ud.t� �\��!
s`�.�$fQXY87�7�Y}�{j���oy?!Un㙓�}��Z7�E�F� ��;
K�Gwƺ�=�>p5\Ř�9�&-=g�T�C`�b�?Iޒ�:b�cޅ��"�	��������<�\����,"Q�0MB�>�$���I.M��Ba�z��,��wi�-
<���53ݕ>~Ǫ���yʲ/�v�<�<ٜ�������&��U�T�T��+G�%����eg4����ޓZ���ލ����G[;�13��ؕ��(/�lTt+�4Z�J���h�q?��>SyJ2�7s�wP��
v������?t�e�g\�7֜e��S%O��+�%W(X���(�B ������uͧ��L����'��M��`����䚕����R Ey[�ƢÓ�ec�Q8�`�jy�Rn���Ϳ����17Z.�b_2�ܨ�+�/-��Q	/���2׶Uk~S��i��ʛ���$�\P�ݩ�U����ۮ�جN�sKz�y��j��ځD�U���&��+aݲ0��g(�i�?��e���������f5(�@P����Z_LO�����<�+��VE<����NP���a�����2Œ��^�)ˆ�bnq+3r��z�K�;r�ρ�1O�DI�Ü��ܓ}�O;rB�n�e���qw��`���g�o��XC"���e�U�Ջ��;P!����k�A H�����9-�h�B��@х��Փ3>W
����?�:�kx����>�$E�Rp��k�iE�T�9#�O0���o�N�"G�dN?Q�{g-(y~��O�ΌB���KL
ϴ�\>nqFqx�18ج��Rn�� J<`Y[k!�-m餺.Z�=n\�M�]��F�F��n�dvyW۳��P:ʛ���ad��u=�Q�
��;��ѻjC��UZn��r�I�m�  .3k�۹��"N��c1�oT�R�sz�*�$��McMVBK����Id?��������_� ���FK��b_��9]a4S��E�U�c��!�Dtrt���y d�5�n��f����縋����%��;�6!x����.��یu ��G�E�����C��˄�����'��da���]�n,@��q�^X:-v�]��
(B��Z �d>�PE���HD�R2	&�2��{E����3}�,}�����|e(K�<)�d5!E>���X���;3	���Yx\�.�My8I��#�V��L����`�CP�+��H�K�5�Dب2u���.��¬������.sq;�ҏ-Y���?�U��}��\�v��y(*�>a��U�~'3��ѳ�>��OCj�9V# {��'8�l�|��H��ց�گ�eD��4�JS=�g ,�w��TF�1q'ď*T���7%c8���1�� L@��s1��,0��&-��Q�6����K���w�Tt�HW�	�|�X[.]����psA��WmEFוP�s�4>o&�����H��/k�|������ࡀ~�r����_�z&�a��C�e����g�u��.6;�����*�46�&=!��Y�����������#?����1�[�}kO�� Jئ%>�I�gKׁ�s(�j*n�n���k��ѕ��@��(+OjV���ha��+�h���B|U�n���?�h�q#������{�14�4nXtF����9&!fQ�t�L�J��Q΄W�6��*�~�@��Rҁ��3�(���q�"�`�����x;ti�l�u? 
�(��n[����\���#+(�	[(����7,ֵ��	%�r�D� 2���]5s�Y��%�+s\�g��@|�N��vW7Z���C��G����R�E�V[࿉ 2��`�(�/�}���3Q��C�^33"�.eV����3���ui+��%q�F�w��|�%xP�!o,T�G�-vhD�O�;�'?�24�+ʦH��f�@ʄ�����%�q���j�	K�� ��������w �ʳ&lev%�ݹ�\���"�Qx�&������*խk�?�Uy{w�����ֈ}��\ŤX�ߋ�j��ZE
�5�$��ѪEN�P���=y�ʳ([^)�`��4�}�����C�r�֞�̅���	�B2�n�b�e�9�M�\OTjo@��>;�G9&�^�ξ������(��M,#U�Ĳd'9��NW����E��h�k��� �����H1G\uN��\�}~�U֢�J�xI�V0�Tw�6~@J9=WZ�s�"*��Y�^@;:���7��j�~�V�+x��{D����Q�Pq�rE�\�%w��(�v<��C��H�s7i�������]{\�b1�Z�X���P�:.�[�X��(^5��2lƞM��H[I]�����X2͈ �9+��s`M�X_����Pu9iq;i��$���;1S�NF͛�޵��b96�*��j�$�EU&�_ޝ����{���ꛈ���wYg��woR�Ak<c
��|hf3Z����Kx�g�9� �����"������(P���0�pZ\� �Y�?��0�x�1�g��0��p�+���i&Q�:a�����:Z5J���8)waqGSWm^��OWL�C+�"���Y� ������T��|9A^���m�U���3��1sŠ��vZX���Tu�>��ѷl�1�>�#�	"�HiI��	��9���q���2�Jٯ�j�h��{���a�Y=a�/�J�����CC�:��!�N
p�D>��Ҋi�.��v�j�Y�9�)���0��3�@]jLO5Z�v��,��8oz�2�g�"V�E�K���l���CJl׀�n����L�8/��\Фp��FH9��MiTnu��р~54��UJ��[�bq�9@4��z)~0O�5K�SK�=kE������#&�����6rZ�%9l����#�F�U(�;ȲL���6q<�$]�����Mhk7`ͨ�2W{�@�?���M�S�{�ެ���|MK(G{�jjR��Q�j$��~s���
���-��O<���)�k1݉���F �M�5q_���kz��$$�%��z��u�[�΃k�����=�L㪠yU�c�\�M��
�Њ���U�nʞ[P\�k����ȴ"+aBl����Re)]�����5A���L�UY17�ڎ������J�	��cI�E{�zGg�i�L�r�rN��X+2"��ꞓ1�.�O�ˣ��9��N��\���ʖ�T��Vu�_d��jT��@���꫄V$AA-��1���vG�[���MGõl(UFl���!���m�^�{�DT��M$9E �/�^7WX�ǔ�������a����ʛo%!\4�va8ڷ}���D{N�U���+�U�߫"��w�r�|m� ��zpFw�jP��6D��~���5v��?K!y�G!��cD��S{l(�6��XT��,�smc���ԙ�u�P��3��Sy�A���M��T�]�{@e]��n/������_O�^rN�c�Ԡ��6x����;^).���d�� M�D7�S�9��aj�(�b��Ca`4y�^$�1~���4�W��#�(��RQ��3���Qj5�<��n�����c�>����4t��7���6�e �R�	� !Jn��d:-m����1��}f/Ap�<���M���H`|[j����,H��;/���z9����s�~Rz&κR�72���K�5?���r!���=ad���C���������W{���w�
Yu�zI	WQ�+ȴ砽a���$�J<RWۍ�_�zg������KC㛛�l�y���$�W2l���w�� �K'gnN�uҚ�D�<c����=�"�AE�����3<��I���:ۊ;�9r��י�43�ǫ�-�����
�n�Q��Ga����x+���kC�ַ�.|e�к�����kĜ��r����ƽKb����@gHm��u.�ϩ��5�~���(��sҲ,"������9��f���[�ЦT�����(��.j�yF>�n�������iF;���,���y�̇v؊�u�0�����DR��������=��"0���%�ɰ�L����d�qX�!��:�5
��iv{M��1�(��-涸YϤ2+N�!'V�I�EG}דg1�����ҋ��uρ][�%���F���)�/�����	dVbJ`��
�����3i���ǆ�
�r`�ʢ���.��W��v��r��2����=�-���L�[��������)KE�G�1�I�!j<��*�hl��7B�^ы���j*3��pQhe}�e�B@YF!�C�Q)�`'���WvC�'E)��P0T�&`��fT�H�V�d�Ğ5<�e����c�i���¶��eNMܸ�(9B�=`�����k�<����ʡ��,k�[+?]�;;\i;͒��1���˸���i?t����G���^����Q�ۂƦ�x���)��_7����F���ƨ��Hk{��x����Yk]��}|c^0��!#�o90o�LK�`�17�h��X��3�o�.�]���}O�'�2�Y>�V������S���K�7t�D��uas��a�8����5�& ����L��칺B��9ж�G +����ga��͋ik�;]�ua鴺�|����Cj	U����(LN�k7M��������Y;ZjM(��P������.�a�i�EZF-�x9#��S9� �DX�˫�[5�m�v�1����I��=��ѐl�!�t?*�� e}�4���o�w�w��Ce��m�(���j�h��U�E��ISX�e��GIxk����\���� ɳ�^��~��?��G>>'�RpOE�A�$�lz�ˏ���#ž�H�v����`�kP���,���JI��K�҇�k��o�F���Tq�j�TI������kKck��B��aR��$��<cM.�=�+�GFόL�餯�����/�U��|K��hfӫ����R���`=��üA���U��I��ȹΘ������|�_�VW���*G��}S�赏�m�kUg�k2��:k����k��{�6aݲ�;ѡ*9 �e}ßHm��t���������{s	˝�.�Y�?fyq� ���A��+�K�Jfu��:@��������뤹��G�T�8�FnXp���[�w����$�>��7a�k��j{�l�Cd2d��-�����&A�w�[s'�^XAc���}�������F�����Ȱ& �N��d1t���$�	��@�I_�Ddn���jlW���Ӏ��#���/\�W�p�x�Rwi�����n,�����8A�h�g�]`d3�&���f1�1²|}&s�m�}��B���(W�p1ā�������	26i"GuD�j�n(��ؾ��6����Iy
`��0%qf�-����u���r�ߌ�G��Q� �+�`qh��fY�ؓ��m��?�4���2�a
��Nj���Y����o��J�~�D��O�7�J�@;�gEF��	�X�S�0	,�A���K`���.�0�|�_a���]�����B�u�)eؙ;��7���ҏ������ag���w&��s@��C/���gc�v��G���2�T��t����tx��3�(t����M�B�k���5at*DN`Щ��)�LS���\&Dv���w���۷�y* H��ju�bΐ��j)���*a]g�B.fNr�x%B�ta��l�,,��%�-l^����1:� ��#ɾ���V�L��#�uѻGX[#�����ze�g�"�9d�![D7R���5C�-�m�܌[�$��S��f �ǽo2D�Tlno�.h��w4]�+/y��a T�[2L�5�P�ɋ�"���ܔ�@�6VA�g���k�P�%�#�Y��ڒ��@�����@����?������) �@Ê�.:�<��<�轡h�G�.2FP�T��VP�RZ�%���wg�Ɉ�Taw	P�\@�l�i�H7�t�Z�	t�*�O��3cP{���0�E��~��Q��!Β�Q�����X���w��5]�����s���֝��q������ qU���v�t�{#�{!<���N	%;A�:G�r�[�Z�=�m8�������#��\q�7k�9����`��MCU�ߚ�Jʘ��d����c&�UT���X��yd4��(�c�����w�&���U�
�Dg�{���8��%�b�Y}>��c�p�0��`(5�T�c�U��C'���ڠ�F�jg�|�ȧ#P��]Ǩ$t�)[8��9����Q3C}��d��|���͌��O�!�m��:����3��e�]`�Q�!0��2>�kk�1U©�P_!|��7N�~[Xd�Q�V.�W����#���O;t&�2}j�璘�?��"*��<N��g���c�U�5W��z@��x2�Q���
���/j�}��"��7Lda��i3vb�1�p�ն�2�s3��X �ȶr+Oc(ҁ�
#�������
˽P���y�A��e���F-�\rv���a���Y9q7@qq�S��p��wo/�XI�P�iR�D��g�o��]�3�)L�(��,�<=ƃØ;*QJ�w���O��4��;ز?�TD��;x0�d�e�;���SvҪU5Α�k�0��$�坵Wė��p���@a3}��{9ʉ��'h��ޛWs�����[���J�Al�P��6��r�����h���R�,"�ŭo�g�~���^q�w���ԊO<K%�	��(�E�#���:���̴����l�%[�> ���Q������o[�`(�-<��vo'&梦&�qsO�JXv'1���G[/�:T2Σ{]��g�DyD���mۢ>3z���l��Z4�g
�.����sr�T/,��&�1�Hajq���~"�1Q���y���Ǽ�ϐ ���%m�Io��q���kZL �6�r{��UH�l7l�B��|z��uwl����E�3���IQ�M����b��Q�ˎRm��0D�76~[�T�O��q���Q�k�ϵ����K>+0���ٷ4��$�<:xM-4|��X��rq�3�����3Z�,J &��mj����#:��������ubWT�Uuᘨ�MH�Ӷ�Ɛ<�+$�r#<�S#�-|�j���Nu����Y�!������H��.-��V�Q3��=�n2Xe�U�c�cCG�9A:���G�-ʲ�?�F�? ���g�ua+#��%��=���Cӯ,=�����b��C���wC�<$#�,��1�����LQ�����@�Z��nW˛څ#�H��	�x���˒ԉ�9��2�K�ocǗYA�(�	�>vT���'���N��5���N�?����Z5��]�m>]?��%�R�b�؞�>�d�ؙM����ֺs���y��`�7όfθnI��š�#�;7(��XGb���ͨ� 4�#�4"u�ǝä�qv�ꇋW�i���C�nC�fSc��������d��2��Z��:~�YT:hA����Qmɚ����Y��P<�!;5��G࣠���Z�_p{���@���ee�|e:4�M(�t+����5a�)p��M�-
��)m|NtA*��%� �Ys����^���;��_3�*���^2JN�☎]���`*����Z���Y���rl������7}FK:�-�r����M������iE9� ��A�p������y��O���fX/'@_b�<�L~��$/�y�`��ùC���������b�<�}�7Or�HGo�'��:me��%	�c�峈�=�ö�,�a�Ad\	z���#�y{��Ѽ�g��.O���3��6H��;���Ӕʡ:��N�Bs%��r�AiFn�6U����ZűG���!|�'8���Z�S�XN��Z�?��>���6�U��ȭ<|,�&�:��VB4�V
���ЛE��V���n����`������Y?����c�`ֵ����a�D��X~gvpo�iٷ۶�R��{Xf��w1�>JGur�p	�^qda0cӮ��>$�D��t�D�>t�$�@�M�|�yI���Ȣ�.�4��_BG���!�W�mi6,����������=b;	:�'~�Y"4y��tE:^��"@$�Jr���׾ӴyU#L�	t}��ô;�� 8XI=Bv����[)�ß䳱 �����:��#�𜯎ݾ�F(RO�����8|O�����/�Ȉ ��̸\
��z`��%��IA����u��̂5���㋟E�Zs�݁��*��[P����7����|��ʘ"�����x�n����:i}Z�iTt�����̥��X#��h=�n쒍h��sj#ܷ<��P$�!]!6���DmAC��-N�
�z6��8�E��%�"P�FϏ��zRq&��d��Ci-?v�4��N#�yE��G ���{E�%�0��X630�huin� H��ACCmx��K�,y��I5������w$�,���QbK�J�$_��U��9bx���k9�vS�2LW6�~�|��`{g���)�Q���#�ϋ���t���)���J&Y<�v�����|�zy v���?�9��r�F�}0�AK8�z��)'N;���j��O �YL�/�I�_�hA-늠�2if݂�Y1�÷DTu��W�(y9�Y�L70-^���Ua��<�����߭GW�
��f`�.}�rܟ��4#��j���'_C����'�^�|K���%g����?;2L?�Wː�GKe� �z�r����:!@��oC�JB���?��;0��h[ߋ��vf}ura���.9,n�N�Ï�4(��Y��ZZ�:�L�[�!���W"�����[F-Y����T�}����z���j6�?�����bT+��:K¦�>��%���PP��$2Z���넁�#,�@��
��9�#��W��HV��n�մ`�׷#�
��90�Z�ŧ�T<��3��z��*9��+�t���!�ezb��AG.X�� a�yX��8�k%i�ki��q���Vn>O>6V�I��T��o*y�5]���8�� DK��&�G�ANUe��}�w��!"�#��&g}'�{+n`�WG%�8*��P�ж 臷���|�<���� Q�� �=aܨ�]	�n�T�(���, %\�x^��#�b̝���O�@�q'.�(���L)��˥���Gy�Vk������7yw�~[8��+�>�32�]-@a�K�� I!e��hg���j�rpz�G��xB�J)�J;��!{�N�Ϝ~�3��_�Þ�=�x��^�Y�q�9��ݳiXh��g�^O��-;����N�=��g#�`}��/U����.��.- ������11�Q�Z�cx�َ��m?�s����!�K�qx+��H�z�q+��Y���<!.��\�#$t|������7Z�Wx��&��'z\�t�!�c
���+"�fO���I�]3� �+>��|��uͣ#~��M�$�5�DK�M�jzƁ����+�T�v-@<��l�2����ߐ��V{;v�HV�p�(@3:�NŰ�#�-��Reh�z�����7�����e�ws����19�Gqi��̈́��F�Hq)��a���:�����to
�ij!����I����'��(W��m}�ܩ�<Kb��$Tr�D�5��M��\��-4,����ƩLF4
�Xt?@kyVaG'�D�cqtB��H�ݯx���Rh� �{�@<�D�����/m���ɤ��nZ�Uton�����~������$�q�Ҝ���@�F1�SOR��;+"Ⱥ|1+�t�E�S�j"Т��7�{�m�QH4���8#��,9~��H�	������E>�3�4L�����UP��*�[-�U�{��M���m�HA/���Uc`�j@V����9.բ�Br~���m\��lAԪN�Q�q�L)'�56�Z�����	b�q�_?r�Ǥѓr�3῟�p�ޛ��9���Yl{{)���彉��P�w��Ax�F2lϽ'����B����/T�08��k�(����Lr� �v����^W�s�$�
&�EM�} �FЙ�;c?"�.��+�t]	@P���w/��oQy�:ds�Z�gl*2� �;B�t��vʧ<\�C�к��f�}��h�an�H45�/���X��L+-�_kb��(�.������/��wF�=TKz�/:>IH{>|���Q���q���1^}A���C蜎Wo����ݺ`����ePj,u�@5Ϩ(�gf�3y��:�p����^P�@�����:�+�B�dݻ��o�{�7^?F?�U�	($�ZD�@p��K�"�(���[y�\��T����ܑڵ��;ܚ�6$�����n�yBOP<&J�R��|tg�}������nҳ�jx�.�಄vg�'p�iJ~�C|]i�#%���I���ʵ.:��0�n�\c���qa�~�R�%M1��]q�/�u��ߢ����p��P'h�ұ�|O0�YI�%��j3��o����D���3�O[�ɳ���]>e��;�y�8&;HYq��_����N�&�7D������Goh3�l�����[ ���X�mֈa��1�፷l"�D[D�Z�#1�Tf�կ�JUFv[U��?F݋6�����¸in��W��4�@���+�@{~��)��z��ea���[���b=O|}M=�K��@D�\R�ߤs:�.��?d�dm<p)R�,�����'#���rԨZ��p!�P,Å��
��m�;_X;��'S��x�.w{ꭖ�~u^\��b`R�ImP��s�^���'{�$��,9k}�9�&R\����[���u4�1E;`����hxfɭl�w�<�;�kǊ�c�w�$4C�kp�Z1���M����}Ą�M�7�7\�5��t)���]� (9މ�+<4V�,�5�-��6n�k���%�q�}4��
S�]H�(�Fz)��ަOG�*w����$jw��b]�1.H0���ç&�W�"&�U!JbP'G���#� ]��u"G��+��"��C8��RET��
��?@�A��EVCA,�je�'E�A�~�z�KѸlh�����+�b�dm�Ai!��F���[�援��� ��{-�:��cS3��"~���<]g����yâk�����Y6[_+�h�0Н#H>IE��
kEN�UW�/׺�t�� 
�xi��<-�{!�j`Bm_'<. ���ͱ
�o�C92	���I9�#9���Ǫ�X "kY��4svN�l���J��<��lv��0\��6�|�c�V�����q���^�����InY��;�Q��>���7E݂�֡��������^�y"�c���dA�ꟀFK�-�ٿ��Y��<��	�������i���+�G`�\E�T���g�r{Z������ދ7�����yV�	�Y�Y&5�����J7ni��0��I�ڤi��@������-�
�#�:z�`��{՚4����fXˆ��K�� �LI-�Iah+Mu�ӛ�xV��k��Zv�ѭ��]�o���v9�3�R�X���קo�������IL�i">-�l(E��rxE�4u˱�1�˨��0���NΎ�qT�,�|�Aݖ�e�����FJ�?_'�������M�o�at��`���Z���8�X�ռ[qj~{̥��->�K��7;�Q�]H��`Z3O�ϗ�o��������<�ɷ�{$LU*�|tƕ�{Q(ٰ����IYd�fW&$y��k
X��M%D(���3m;V~Ѷ������LR���;>Av��%�s3�2�p$TJ��8�Y�C�������ga��x\h��~�a_�2��[�rP��:1{��%2��g-!��	T��\5G2Α}|ps�B��X����P��s��9$�w"C��#װ�1H�쪧�3���ڍ�:�@��Ez-��ǚ�H�٢�G ,6��f���}$p�(3Z�*�=��)�~6��e�CD�B:[7n��e�s���@\�A�� �rJ�C�﵍u]�W�K�`�4i�=����%�f�9a{�L�-��6q�|�f�Q�:�~ص�K�۵�v#XE��b>,U��vn�a�0�32&�ac��)��_�u`]� �>Ro���k�!��C�#ot<l��A����@�O�'H��0ug�S�KL�����(EU̥�-h���;����C�=�C�P�s�*ì^�8ݝWU2����1T��%9$;���	e����A��o��ܧ�������1y\D��iX�K�������Q͘eϲb�n��}�^EƧ�6^���u�)u�'ʱaB������~Y��%^+ �'���hbd/��c�降�����x�Q@m(�T����G#
�Z�1H>� $�t�v��_�.vzA��8"� �8Y���Y��7bP��I�<"}�:}�@Q��3�v�(�Oz@M:]��N���+n؛���+����K�ZY�����c�zs�hg,���H�,ë�E��p+���/P��}���&x��Z�:̸}��'�	����67�JC����)��8M{�A�ݾ��0�x��|�#�MMob�V���N�vv)�ox ���k��c@�������]�0J���i"u,mLT<��pxi��vb68q��5��Yg�`8�xt�I��� ��8X�����M�Eh�	-��+9��lC�h���%�%*���n�Tr۩%ׯ���4z;H�Y�����`L
O$_�h���VWa�-�*�>,���w��bp��y�&�w ����MC�A���$��,i�Bצ:�W&�_ֺ���w+5t}OOZgd��L�����C*���B�k��>�_�v(���qێޜ�.�TIt�=S��A���b �K,!��ЛJ�`ϼ�[�d\��t��!�8!����<r��߄��� ����I#�+/��=���=����4k?H�>����d�q'��0��s�`b��1l��'I������[�,A�Қ��HܨƗ���������lͮ+Ը�F:2Y����CId�ވ�0vF�9�qtZ35�US��	�6���#8��:�k���e���<�xc�f��Z����h3���upv��O�U���Fgѧ�nᴋ����S+dx��b��&�6Ig���`}E�]�� :����V-z]��O!���d��B�Pl6���P��Al�l�I8٘�&!�=X��9˭�{)�',|_嵹 ��9w�>�����q�?����hf)��xw��i��#;
}Y���i��E&�|+#�W�vB��3��@�c�~Q���f��� �9���C�y}w��l3�Z�9TƇɋ�ˋpK�P��Mߞ�6�a���d�	�`����7�3`~K_�<�.��)�����$0�j�x�z�A"h�wէ���` ߵ�����2j�j�%��g������~)�ѻ�{�oqd�މ���%6�r�/p�Bc���3=�u�)KI0Y�d���B��׊��!I��i���8���W�@�,Q z�5�G���n2N�^(�r�Y���� !LT����x��0:��9�H���_D��'qk&�D��?O�߁�9&FxXdS3g/���sLB����R��H�Bmq����nBС�s�����z,�'<��c����G��mTt����)c�1k-���6�ME��=>���Li�0���IA��C�eƽ��j���BX����=�D�\:����ߋU��m//��S���p��A���^>��iU%�I)�=���>T��sW���sx������_��G�1Tl~���9~���,o����e�Q�;���*tVj3n�Fȩ����>��F�URk�=^
���kS�^�D�D�~�gm�_�e�� y]e�x�,�[�B�_��	���^��S�U#/ڌ>��)��~��(�R߶^�$�nJ�8� ����u4O�)���h��k�nEæ���
|O�G`���M�Lv�یo�zkr����#�D��\��@���-oCE�{�ؿ�k������)10(�c{�
��xֻ씬�6LI']�N����H�ܞJ�E����ml���l�<)�X�L!����+I��0}Ԑ�B�9��@Yo;�TRI|#�z�g�"���Pdѽ��}(��F�A=�u��|����
��*T�m�N�ܮ��o1:BlI,w�J7hA��虳�ϦV�K��{�YW����f�3R_��̃Iު3�r7`��@���25��m>I��'z���(�s��U�c��,�7���p�,ڲ���?=���������Ե�.��7G+�jR�7��g�>}'�ԢK�����?���2f������w-��y^����q���!����vv{K��hgOWD*�}�y�������D?!���FT��n��Gp�f!�i��p�R��ۡ`�+Z�Q[��TcH�������M`#MA#��clJ�x��Y#�oFt�A�E+H��Z��gD���5`hM�$?UЁ�� �W�Z���w�}�>����f��c�p�es���vT!�R�oP(GR�c0�K���{���|��P&7F$�6~�����Rd�I�6r;+���@��w׹BE:��TT����g$I�:ZP���T3�A-�f�m4Y�o�l1IY�2d�<�-�T����6��)�Ǵ������8��,h����6�7��.2"kvoTP��w�W%}�3���'��R��n�4Ҟ�N�x=���?�U̺���T��Z��X�C�0��A�!A�D	�=1������$8�M�q]Lӟw
�M�s\@�̓B��� ��!�?��t�lߧ������.ҭS)@T��e�x�T׮xlцC(�.2x���Vf
L�טp��#=s�-��?}�j	?=*C��3�U]l���Y�����м	���@H����],r��޴}��N�	P��&�,&o&V�+���ր=sy�8�gp��"�kk���d�n�[J�PYj�F���锬�m=؏`x����A�$獠S�p�X�":me��1�y�0��o"�v�R�1�d0��3͗��5(�.5S=ݡ��������3{ �5S}���&/���:e�����ZcCb,뷑�/8~L�!qe��Ƌ2Bw-���r�k*^���n\m�_ޢ�rme,�%�[�A�JjՉS6T�=���8B�XKl�WSt�a��d���ov�b�5g)l1�� \:dHIK8��=�m���N�y�߆�
�D��#��	R����xL�p�6jj�8N��.��>�cl��@$��)�R!�о��l�Y�ן�E�<��G5b��������{�lA�<��@(V_�t��%b �eA!K���\�;�R�{-��U�u�$a$C�!�;QtҨ�P�#���=+�Y'7ZC?�D�u�"�p|����uD�pJ5HDgf���c��KG4R�^��&�q-��א�Y�L2V�o���Lyz����=��f�3�q"��kE�HO�RL��LR����XI܇����ԦeQ��}���~�1�@l�s]b��4��_��B�NP\q�80U�|������y�<-�{�9i[��b�Wʠ��i
�g�)G�BJ�,͟~�`0���%��Tec��´k+�~��P����b*d?E������qew��<^bzd������j��׮�X�HB��c{[�%겙Ϋ��&�s]�ad���PB�P�)/&S�
�7 Dm����bjݫU9�qx��d�7v��HT \^������.�.��L���9.�|j��c�'.��R�����	p:�w("��B	��Bl�y��[��V�s�71��ã�[\�� �B1�Y��;��o��%&Z|�j��S��;���}/���݌$Ly�G�<� U+s�6��$(�W3��K[�+�f��B!^C��V	A2����I�VJ,ĪTq��Ť-vAqw��e��������B��%����<$�x�^S�	� #�&�6H�O�� 4�h�9̬��c�2����6��6�4�}30qI�D%5k��`3�#��%��᱒?����j3�B�斈4�yY)�4����~���ѐCӠ�%���`.J��\6��m�~�"�q��Z��^c/A�c���H:�H"x
+GjwB�o��B�R�����{	ϲC ������ �W�5�}[�\�Q� �b�q�iҩ<���-�����6�ёsM��Tͦ週u�߈���w��/0�v�.]�)��B_�4TՇJ��m�xLGz���}mK�Dh����郲K�Z苌.�Jh]�|d���H�vU�Wi������mQ�+x�el�5r�������JMHٓH�m��)�?u�!��aʾV�r3,b������|���C�k�;̊�R�܄��^Z���Q\$j�'ؓb��X]XAv	>�0P;��X�`ꅂW�qM2�/�DR3i
����>G���
TÐ��i<Cr͠��Q����,�fLHV��W'�_3�2��P^��o����_�I�!�9�;~�A�S�¶7;������B��W�?T1n�^`� ��vWI�=p��$�ffw�q�b{%)�;ki���	�i�E!�!�Gx{��yֻ?����.�}����0N�^�@
䂴�l�WB3���0���
�}��R�{�ɍ\�<ri�4x.�f��)
�g$m��u�+�Rӡ���/�噺}���z@�1"wΏ�]G�H:���,�������;f��7��u
�R�kGw�����^A_OQ�D��GsQ��f�5 ���c�ݧ_��B��]���f����D���C&f���~����c�z�9|�S�ۼ=l.���'<�A?�o{Ubn�Nv�w��Dʪ��1u_���n��+:q¼�Uʾ`�KŻ�|��+9�����Sh[��t�N�eo`������4���X;=o����,��m��Z��ש�k�:�'Uq%_{~��c�ZہL+#��-�a���'!c���I�q��E=c;DY5qi�l�CjU�+=٢v��@�U���7ި�V� �+����m���y�{��3?	��}f*��y=��
�m5W�Hg&\�h����	P]t9��\�U�_�GhП�|������o�Krd�s�7h�����y�V��Ћ���G�`����8��5V6^cY��ب_�˗eki��'Z=��q^%�s¸�o�k�tjSO�,3Nc�;!+5�,yq��n)q.�õ`No!�����S c�ڳ�,w3],�v|������Gm|�t7���`/�3Ǭ� 7����p4�I�I2��ZaűH �#�	^�Z<S]�����X�ZP�h�,�ׄ�Ek*@���z�[�N��x�/+�b������R�1d���y���ni�ᤐ���$c쫒"͜N��<!J����3"��@�(]���9Ը��n�3�pI~D�t�k�ؽ�`�4��������?�&����)�	���]<Ȥ� 2T6j!��7a�,����{\)�ȌeM�Geh�/\�.i3��`0�����R�+�����z��\\�N�&��Gm��uR/`y�i��:wl�5�ua��)�n�m�1$G0����5���.���2]�T
���mi"]P]JCq]M�o�u����Fng��C.v�OF�~��ݞI7ɹ����Q� �?���}�s�;�e��V�*3-�� ��([�jЈ�����V�~�ZP8�ǩ�io���_�8���oV��:��:�K���aOؖ;\9��Y���の6�b���!��z�hAQ��Oۀ�+����P[�n��6�Nˏ�e��Ae�|<~a	����L&�Ҋ�_~�.�kp��W&u���-v٫�>�
�"�}���y^�����H���D��. E��V�A�On���	Tg�ul�Qz��6X�<����{��.z;��R�˚@�|但�NB���8�S���mR��ɏ�N��tpǜ�+;D�4����O�Zkl_l�-�LS[fu�:�W���y�P��=�zZ꛶�ӣP��~2���ȂS�}����a������fL�Y�!��Q�+|�a�G�;C��v'F�"�m8��)4�BK��%R�X;����]a�P<���B"L\�
�&n/zs9��<�6���s��O�j��z�=ew�Ƴb���	r�A��WG�eG�v�|���r!�*͝��RZW&`}���X��#�ƽ��H�Nhj�Q{����y��i�^?�	�:�N8����) *����.ў��E���9]�)S!@���N4�Zh�|�ί�m9s�z��n�ǜ��Y�s8,� �_��0�!�p�������<�u�:AT����0���Da�Ib��ҐL2"��c(� yr�b���2�������	 �LY�V��x�O,G'�q�K���+M�!�K_P4>f���	�Q�[S��>ܑ��1���z�ĵ�P�;|�7ES�� P�ש�����D�Lt�9�&�S��<+�CㅛS4����u����5�o��g�*��w~��^��nʁz�`��:i�d���"_t�p��ہV!C��<R�{څϪ�A��O�=�������g�� ��-�kV3ITPn|�2`�s�;f0�Yw�?��@�^��&<�c6�󘱸йp||�I��13���m�|G�X���-�L3t�(�۞iB�ރ��~��Ҏ���_5+����s]��C���j�u��������鐢3�.E�����2�A�D'!3�6���Dtd\j�M`='`���Ahik$*(PzG�����\46T^�3�t.SA�W/��!��b��:a4w�~�ՌE�х���P�ɝdnKj$�<�jտ�~�-�MVşcx�߰Q�+�S2Z�����:�0�a���&5����$1�t$2�BK9ھ4t?"�o�cҁ-7���z�>��9��뙯�5v�{2��	6���@$7�=u�`�v7(���|<2-��n���%YOm��uBzU5!���@����
�\dO�p:3	�%pQ��<p1%5��]���ͷG��m�dc��NU���3h`����ÿ.�ҧ����4Dq����h������V���M����e�e��a�ٜ[6�1v-�N
r��$�oUp��~n�]�+�����6����m��]���h����+u�z���9-[��c;V�8�Ԣ{�g-��i;�]�̢h�J�8#s��,N�$���{�;�1]Ȟ(�|,����g4`qMC.�����$�5�qgr�;�H�M֌�y(��|?�pa�	�Y�����չ��dVZ��%Tݟ�����t{�Ż?p�W ڠ��
}�
�Ef#9� �9����<2=ƎQ��/*��	�,�*ly8NI�X����t���xd�/��c#��k=�R8J-�9Q�jr�ް�F˓L6� �<�2�S�׌��p!+��<U25��YG���O6/�Ήӧ�|x㪋��G���pd�t��2�s*�I�o��ی���I4_���ZB9YrRC�q0M��Y��V���N;��ܤU��4 ����G�Pr��9����*
�8a���Y��0��҄�p�gj*nc�?yѶM��0�+�Q���j,�]vC��h�s�Q��q1ܽ�!�Ҥ��p�'Ǖ���0���̶���&Uk7GE/'w��d���]��\���AI:J�
���a2Mk����fՓ�9z^LE�S�<�[����^�>�҇�1jfȳ�u�}_�a	�B�����ģ�;���Y�$�1�v���EƱ�sƀ�P��Q�I>�TO�����s�-��K2�{2"ʩ�֪Af�R��nm��}�'��	�t��Ϡ"�'8w��Y�"�>��M��,��!^�h�w�U�MY9n�<�yiI�'��]<�bέ�X������sirdPz�XQ5�"�JV�]��S�/X3��`�;��6� ��j$˘��ٛ�9���1������_0�Sg�j�i)��� �#/�@�iev�ŧ1�<��)5���"��ô3SV%�+�if\����{���H���)�PzɧC����N����p���O��{#B��x�K+�^	��]Bk��V�j{�1Y/b��	*��,ӆT�̽O�� �fp��S�Q�)m#���)���8]�뀳�!��9:�+�}�ʤ�z��Y����i���TV��塚�'*�t�H�j$󶕧��������M����/�;G˾?���ch��E�f'���;��.�g$�O�⥹�B�V���߆���NFZ����niM�+�8�ԟ�h��i��vWL��m%)�������i����n]#���GT�@Nb	�����»����G��q��%��I;�����q��)13;�J�e�X~�&3�+�2kچ���"�ѷ��w������� P,(4Z��=��-���50� ���+�i?P�C�'TƜs��.�F+��NPsi̎�-����m讦�a锸�sb�T�)T������G�7��tKg�.��.�أ�������-f�6m��Ȃb(�n�S���
����ÿз��ք,x^y�� �x���>I����	�G�8�I�T}Ԑ�1 6Iag�H>��+6���A����� ��cu�P�f�U9��lR��c%��2(�˦|��9�y�X�)�D��.IR6�&�䉟+���f�6�m���ˆ$;!nQ���o����d�X5H#Yn���Ӟs@�1|����T��u����
Ƞ�Mk�4w}�RiI��pZ#W
ՙ�s���Aθ®T�AG�O��S�5��� � ��ޠ��6w9qX������aҕ��w�s`1dqҷ��r�u;h6��`�5;���hi �z߳����X�7.*��~�~��n9fλ�0�$�5��Z7%R��q�Q �j2�\�_���k#k��
�C)N3��Q~��O�e��]��g��5�k���/حx�* �ֻ����v�Hf��	�����i������{���Rɰ��i����ҳ|�yxI��c�l'�!G�x&`�.�%s��iD�t�Pw�K􍠧(�c��&�璅�^�P4��ڞ�6ţ�#�zؐЧ$ou����nSl(�Y���Xs��d�5�&n��a���i����&;�0��ok�]�	���":�>x}���V����NZ��]]e�n�b� �U+�+�a�����o6�yf�����6	%���$�/S�"�j���Sݲ�;��vC���C��1c��8W�Z�?��Im�xv�1���ٛ����\6��� �R|��W���@�Q���<�xv�ME�z[�s��܁���0JZ��^��g��ç�5��B[���Ռ�PV*U���8�g�Cc��H/�~��D��B-�J��c�=N�B}�_��O�Fl�,��*BV��P�g�X/���i�M&+���i0��9u��x��:��>����nƞ�����N���4e�HH1KV�� C�'��5�jl�����yG����A��a|�Z�hh��L�6��\l��K�%`s��� ~�s$��S�Ψ��T���+�^Qb�5�;���c39!(b��*�v��:J0N�����.�t�3;ȗ~
+�S�P��G�9�7�����}�t��	*N���q���j�oT%?�G��j�X�Ƿr��<�gt����Z'����IωZ2i�Y���O	������E+*Z�E&��)���x7�������	4{����[D�&�&멥�-Vg�`SiW8��V�rÑ����{��2��m�RE��B�Xq,��Mry�?�5}9�?���^�LS�h� ����Zj'�j{ T����jZ���T����-b�n*VU3��V����k6��l e+��,B{l!��N��U[�I��P�J�p?K��횩È^ک�+�~��}p�����RĚY.��2FuG�h�%�5�R�?���/���L�;���ӧ�'��Q�m�H,@���H
��,����u�P�V���%�T��� �[�&���|��~�(}�]��w�@�Al��+�Ր���#�djF�3
D:7�E3��iKKJ��G�!7�˝l��)�9�*�41�[1�c�:IM�
�`g�[����6����O�|}�rñ�i��B T�*S�e�(	���M'CZ��������u��E%���g�&GG�+�������C��Dć��I�&H�'78)o[�M���T����}�lț��
g�ɍ��]A��C҇����r�vIEII�!�o�ȃ!Y�rz�O����R���UY�x�NN�l��UB��-���Rέ���y�1	\sH���v�)��1#~�v����K�4ѿ��Ҩh~=��/��w�Ϟ��6A�օ4)��u��ZLڲ,�J�Hv2�Z��YH۪�JIA���XV~�����F�r�D��q�fab�XN�2x|�`�)%��q8�a+ȶ[��:>*!Tq�ʠOu�b\�*�M_��b�ALcM^���Qc�å���b-ϑ��	�D�uQ0*�͗&Y|� ���2ZUT��Mp�n6���s�1�GA��;#:y�d�܀����)o���w���F������8J���ߒ}OF�?�u�	��][�y��3��҇��Ow/L3$�h#�C)�rqr~�5H�v����&4�*ˣ��T��"/�:�"	Ms��Pz(�����@�;	rc���ȩR���h��(fc�u��2@���/������GQyF#\��-A���3K��u�W����,
@���|�O��Y]��� �+c�����x��9���삼�����B���Xje֠X�q�dqB���EVd�����)8r�i��}�b��B��N½	",����d)�8<4�"q3�=�Ƞ�s�.� m<�MjY���c��B�AE<�TeS�s��_/����+�Û�y�FH<|�n��Ro��[����h�<>.T����a`�4[x��?@Gʚc��v��t�0�̹G�팠1�B2�^�`�Д!ɱ��������-x'K�ȶ�f#[�_aX�;�����/��j��cL���ٱ�j��3,��#<�,��mF,�PÉ5M(����܋�����v��եJb�5D�N�;C�?���~x����]��}.>�e�KM���ń@���b��(<���~�y�k]G�� `"4U�iL��,��ï�E�%ip~(��$}�]�6C���_��%��g�Wץ�6}�Gd\�+p=L�d4�#�`�Kg}f]BbV2-�:��U%Ta�FkP֬_9��Z��(�3�O�)��Z�eVW���/ky�	��B�ޫ�����l��*�f��=x�������S_K�,"�c��-�<x,ri��W�b���
4������i[8��=>�����w�Z~���OuK懀������싪�7������S��i�nQ]��M��0]@�E��Ѻ/i�n�GJE1��Ҫ9��y"�>So��JZ���O����}Կ�[��#��'��㝙���B5���b�"�q��D�x˾	
�_��q��r/}x�i��Z��Α'tǃ�%�^�� ^؉pJ[\蚕9>��n��pu1�tZo�K�����]�Ѭ�E=���>epH�x�!n�rc&��=/!�v~��-�T׺�Z�̺�Ow��B����dh�6�'ج<`dh/ ����*@��.u9�L�I�B�u�e0�)��oj/���T�E*4
�d��m�(:U����,_��]��g�hF%k3$�k�a;�>N���?NsLP4�.������G�8I!���^PR�rɄ�:
0����d��G�2�]��;�B�-B
؍�:��c9�&UIlDÕ���P�B8���9ċP��ng�ϳ�,���{�67ˤ]R�ÒIm�����6%:�rXx
��FL��^�p~�W���@P�&}	Sj��y�Vx���;�|��gV���:B�y��iԠ��h�mK��-I��P�f�p�o
�nA�=-c;sXq�tw�E�]�ۨ��iB7�.��)-��Ȇ��,��۩��Q����W�'��c�!��U��H� '��Ʒ3�Ϻzr�:s6 9AV �2� U��m��
2l�68��u'n��C�/w���^�(5� �#~%Vx�{��U��|��e�A]�(cՄ�g��琏6���E%���L�_b~~����A[;8;��u'3t��0o��33?��g���f�h�`]kl�L�&���Q~)����+�� �䩟AK;�Uǹ����0�u�!.s+�� ��ωC�ƽ9���z�*��~�Ju[�24U�*.t�7��ď� �T�EE@%F�mˎ�d�J�)��a�
�諮��3�qoc0\����u�ea;��R[��q�n�� |b���ocm?�kv�*[e�﬷�яZֆ�P'��
�[qQ쓾
@c��x�������rRE�����V=d	���jC'���H3�#�Bm�X?�:�6C�z3��[�ic�2�<��@�Y�#-G�&U>� �f�D�[w����z���u��3�/�#
۾��\tASF-�4-R�ЁB��ll'L_[vy�p��z���%���is-�V+E�x:>���<EO����P��9Z��S�`�$.��3z��YJ���+�c"4�ߵ��曼��OvU�o㤑m�1{�[k���
��iEaP�F/�'�4fR`�H*#^�ܪb���'��G�P��Q��-�_�z�����]�r�\S�5Oag���΅��{!��{���E�����*|��O��CmHJ�6rH��o�;�����Wv�uqѪuR;�v�a!V��1%���	/�]^S(�"~-F��$4����q�9��ڽ͆�M��m��G�����/�~�Hb���Æ�xt���i��Bn�d fWYbȨZ���I�z��h�YiSw q��C�صi���eY$���ܺg��zګk�{�����{�'�pp�7
JH0��t�P��<h�0?t�G�E|ȧ��c���7�.lT���ɖ�� �I����Д[o��8����@Y����wl����q�@�a�w��'ja�&��۸RHo�I{�V��8��<7��`�7#"��C�����
��Gz�(�L@���&�6���ޖu�}���˳��eݯ��b
/�']ɱ�-}+�zJ�Zs�YU��KW(7D*���R{8k���O����I�mR�QU|�6��F�b��U���z)���̨�Kf��&����BYr;����3\��d��(҉��O+���g����x�ˇ |J �x�y,��J�siԅ=Ң��[r��ƫ���lt���Ȱ�+�b�"z�{>%�mi�J9`eȍ�*g������s��g�W��hj�ԉ�4n4����@S��-+��f��k�;��6��qn��]�46�y�|5�K���bWݱ�Ht��\���^/��̾�]��,i��A����"��:��BB�@Y�B��~�Ԑ��ml���'g�7*{��/?��d�Mt��-��U��;�N���ad8�_ܑto�l�y��x�f��������=^t>�К�O��4��ϱ@c��\.���+o��S��|P�c�R��Q.Y	�(���I��!E҇��r���=���8m�ӧx}`j��z��(��Ƞ�<��k�"
ֲ!d�+��,��P]:����B�/�`���a��|g�ƨ@�<g��O��P�� ��R�d��LR�+*)���\�#��{}1G[Kr���B8�ʥ��5�Mu�祫VJ�� �p�D3򾮯b�R~�ف(��Ǹ2��w��l#�:J�PJ���f{�x�
�&B0Ya���U��f�B}�5������&���^�j����e[��?�������~<\ 戶�4�O�<��^�8Z7+ِ�:���;�HdV�0�:J.t��f�蹄����������9gmë��=l����,�-g��;<��2�[Q=�������e�!�����lK:��4��M�KZ�.1Cj��tL��?p0"��G�79g�A�^W���˘Erw�]��l�~��c;����j@u��5�'ȏ��.RӃP�Y�'��erѨ��k�f�Bf0,�+s=&��7��C��ul:R(����)6�N`����|_��;N/�|��#�g
rh^p���#�d�>�'$?��zڍ��[cM���j��"�PJk���Q�sJ>ŽTʄ@.�dԤYvZ\��jT�2b��<�K!K�P��v��=�2h�1(J
�#�^�b�+���'q����|�p#G������M�c%��fn����ǉ���|@`�V ��;����}�b���_�z��$+�s�p��[)|&��Tm�1�^uh��`H [���4k�[����P��w$�U���?E�T�o���,V90�݆���,Y߶ǫ��_^a�=�T���iz�^rŅY�{���h��������_86/���G��.���.|\d�*
�o6|g�!V �֝R��D�>�NkXm�oG�ΖOM/MZ X$�Z],�܎c��KF���_��b]&s��,����^۴b�qq�g��Ib+�j����f�4��jщ��̐s����w)����
\����%'�֐����%i흃��� R�f��<���cH�Ek]R�t����azJ
��7%ۡ� ��N����-�HO�G�6�[ݣ}�[��+�y8��Zh��"=�bX!Mg����)�ӜK��+"�eq��rz�����S����=}6��Z�H���k�H�%��+Ny���
Z Q�$	@5.�,�cC1�D\9xz�V�H��o�u��D�G_��o.@�n4���b���̢)�D��JI~!�b5J�����b����0���8�|�&�)<�61հ$���B�"#~#��6 r(�˹>��v��;���Yv��D�h)��p���T`��p0�����	[4GO�Ƀ�Q���Xݳ�S��9EXJ���LP�_�,(�F�G�	����A��7k���ż������4��	��g8凟�`m˘�[�S�n9�y"8z�|�$q�s5+��|�z�nV�ܣ������H�p���yhQ�� u��A$©!�/>d&t\����!��������E|��˷S�;TtC�T_��	 ��C�i��hS��eG�*ϙ�O�E�� ��#�n��5s��xy(��>�X���ޛJ��	U`n�>��v6K�}���x��?��C����9'H͇w�o+y���
�O9�S����MZ��S���UHGp���܇ͩ��bŜ�R�?���l�A��SR����Z��@�Ȝ�,}���`�����_��5�Ct��%Dd��02-���5��E�d$u�ۃe2�4�L���ߔ��b��6����Xg0��1]���c����\H�R`���0y�z͞ �*�����b6�y.�wt#�v�
��&��]��C.��H@�W{a��՗�ѰD�C�} �q��"�
׸0 +	�t/��[}�!�;�G�z��x�e�{|�ܟ�1�|u�c�^�Bb�� <��U��l<��?�E���̕pƆ�� W��6��TY�y���<z�	*'�_��YH�;���~�
v<!�S�V2�1��Gc���n�
c'%�+@��tp�9T�y��k��p�,�N�?-��d`����S��4�b���C�)ip�;q ������oҧ`(��W7mΑ��;I��B�	�
�DL��f)}o��	lj��Ӧ�UN��^Ź�Wt��\S<���l�L�f.��!O�)װ	�B�H$��,P龬*5N�ZQ�vmד ����9�M��! �AlÈ�p�@b����xS��kW�cLV����Mz�\���s�2��!���u��O�*�|��^�o����:��������4�T�pl~��@��~�
� (������cN���Y(5��9^[Qy���	<�f�ZG�}�t��v�f~�(��t��P4*-��ls剰�V��ov@�'���B!p!�^��F[��;�Ë ��P� �Q�BO�Hq������_pzm�]9���gH��p8�Q�����&(���|���EZ��E�l[��U���(��f�)�џ*\W"���z&=+��b��?��2
������J��Y:�s�Rc�X���v�W�y�X6�Rm��P� ��]����d,��n��y��-��˻Du���Ԕ��	�nR�-��Y�|� 1�U��A�|��ny!�X�;��yI�5�Zb�0{$ᅂMkiY���S�!�	���{V�_H!�iV���j5�.(^�4p)&��݀8���G���?b���j_�����
��3C�2�T�DJ��,�[��@�����U��z�j<��7-A�n���w0���	�5C�h���?C48�/�o�:߇,?_,j�1FF���%�Z��w�������x-�<�:J �wI�x�M���v���J$E�u:B�x^/�|£k;v`�m���Mh�K,��k8�6t��.�0~��Kw�l��`��/����P2�h.jٰ2��S���<�%��2�о�2V�&�tL �<�㥊��������;��{�Ԯf0g�U�˵x��̗��!���;��l���xr���ɮG?WֵA��]�=}y���㘣�=���nI
s��
L�'���r��| 
H�p�|� M8�?�ƚh7�+��dbeqP�)����� �H ��F��� ]O�n��:�w�9"3p��!�p)�R�W��{@��F�;i�W�iDdA�����Zڙ�iay�8�+F;3|���bK�� �^������P��L��2F/���,&�]4�l�����Nqٗ2!v�쾘�f]m;�9(�G{�����&�BD�Rg_����"�^��
$�zA��/Dm_5��h�f}�C�u�6,�iO�"�&	��_����% *��䘢����܄��`�x�M.ifO�[���͏���A��6�ǥ����@��/N��D�+[�)�7TNJe�0{�kD�9څ�25Y������c���D�Ҷ�0�̏4�\�4e�n륒��w�GS*���$$L�d �~�4��C�9L�CP�.�L,ì1J-��p!|�^�C���k��\���=>p<���Z_�L�ĕ$!��c£dU�;,�H�΢�`M#�!#2cr���r���`�[����CL����gKm'���7.�io��l61��zm%�ܴ]��٤G�Z���Ռ#�Θ����R3	7{��xo"�e_�d�a,�g]���yl0�����!�����ܟ$5�{��߱H0K٪3�Ȗ��{�i�AU԰�6��a���ô#���\����Q����%I��7,t����D�۰N��{z��o�ʾ��R�?���c%^?9ň I�90�*��윙����e��ú|���~z����mG빘�Wl�s�*8v� �;�
�q�BR%�j�gٸ�lxvv��a�-;�[v���&I!Ѻ�$
���hO�{F�zj�8NR�4y��?h��׺n�?B�����N��=, �����@��/����uo:��m:a��'r�Q��֊��r�.�,���
4�b7���R�0qq�xg0̷
�b�Pi���mg��4��\o�,�g�n��I����ä���>s�c���F�9N{�}��Q�]�t��9�����O��NS���ikn���V�+�V�Sݷ���
��pl^7�{�:��Ph��(z�f HX���Qrl��yGV�ܟ��iAK,�<}9U����������Z8�T�6�&cZ�Ǽ~���>*�u���f,]CY���<H�I��m�{�G��_�Dɔ�ȍw��4�?W�-2Z��!?t�zB��GR�+s��G"�L�}"]��<�"O�o�щ�/�����/MB�U�糖�}�8v9��u���b�.u��T�;�r��|�|h�Y�:��g�wt44�z�� ���7UVs����|���h>^ԋj\2k��8������c� ���,�u�Ց�7�4[�#�����3�|5�i*e!�������
J�j/�Ğ)"ܛާ���ӷ�R68�)�a]$��1u;z�@���#�I���} 5*K��l4w���8G8jbM=��t�r�q-�61dRZ(����P!Jzu�~d�i����y��9|:��t�O����	����VCw��Bܼ)9��m��y��㰮i}N��cc�-�@�\	�gk�ʉpZ�S1п����N�k�0=�	���nV(V�XN-��f�T�.�X{�]`� ���ސQ�d|N=q>�h���O��F��(x�po1O��{��e7�h���b�X��c���e�"�ȶ{�DU̺�A��'8�\��	�0\d�#�����W�m�����s�{<h��a��}�-q�:Am����th���䙅�#�U�kƕ]���B?��w����60 ���~7]�l"�����2(mA0ې�@�ҭ:ӳ���E<�(��U�R`=G������"�0l��P��(=��^#��~x`�����)R����Q��2w���l���g� +�ۧ%^WV ؊Y�<�P��^[�N`�����ƹ�Ro3p_Z���:]
��L����}E���u+��N+MF�� {�|M�n�`�LǑ�Ӓ*Sc�\y���s"��3��Daz���4������k3|�� ��n���$�~���?)/ �/(&X2e/;��C7�d�sa%7��cRB�X}�bI�(��2럗 ��~@�}:�\�1�8��Y�a�3P�7�ޅnL�3���i[�ʦ��n��^�F��e^�<�"}��稙� ~��5�I�n�g�%����k ��@��m���RTE=���	�"��Y|u��"K<���1 G��0��d!���@s�E"1�;߾��-�ý��� �<_���qaf$+|ׅU�_��?NQQy.�o���I�����6d&*��"�<Vq�>���>`ݷʍ؍����o>}~�XA����:��٦�mz�"�����\��3�{���^��`���c�]~�T̷��i�>Q� ���C%R��(�`��	���iS���e�����GW���* �[�i
L�:%�g�j��"2[�c�����։����t.��ң��<�"�VT�Tk\Z+�z����|�>�%޾T�Z�y��������|զ#ٸ���>m��;{��e�$G=�l����{jl�p\b��!U6'���zÏv�o}�Ң�o1͓��APvR�w�^@ޕw�%��|�q�`������ڂ!,R6����UU���� �*ivD D��7�%��]�a���A�j��ZuFͺ����\�u]�1�u,��仛�k`��e�~��HuU�;�'���hm:��b+�l~J3�t���RI��Vǋ�:<�*��7�k �z�s���Qd%��ث��yM쥠y�L%��
�?�o3��fN��n����,Ϊ1�|;�eV�Ux�i�$�.�+�#�s������Y���+�!D��ܽ �|<���q�����l�l��{T\N�g�!���MG�'�TA��o�4�5�Iz �
�Г��"��"��y7�!@�'&
�3�`���i���X���]��1wXȽ�G6P��#*i��_��\�V/Me��˵=����vX�K��O'�I"�G֭Fă�z]�+D9�:p,��e �/��No �i�1%�# 0�G�� Gh��^W�3�&�:0�S5������:����(���bTDҟ>��� OPu*�Hl=�a�q뜯��)�Bl���$S�.[#1K�Ɂ���q�v=�#m �@���s�DTR*�ɔ�f�6Q����UK�_
��g���N;�d\2���2:���������f���w��T�C�xI�T���뼜�;E9���RVK
gf�=�݌���:L�i�����.�ա�/�Cfi�?=�.5�?��n�*��9'�poC9]f��IZ-̿�W�G�U�c^�����cD@��ּ���v9���
�꜎s�z1�hr����.9 �yh�aȠHY���3�Kd:��l`�w��P:���g�	�Z� ^\�P/���dn�à%�.R�e3�9U�4�ǧ�^E�h`|���ˬ��"���&�]:>���	�d[��u��̷4Xh�
��eh�BcA��7c��{�NM�9|hk&����n�e-7��R,pe~�h�l�Nu�*��RD��&�NFH6��=M�����$8e���`��~�O���tP����泏�d�EL㗪R�t��fA�����p,�P���pBEt������BQY�c�ZA:�,��_ގ�D�Ѓ%brJ��Q�rm�!`�=d�`QƵ`ݧ��b�ה������$,�)�+�&����i�������C�]�M�Sΐ�f�"x�?��g������#5xG&}�cۯW�}���j<�"Y��d��ʔ���� ���Nイ{�%R�HR�Ǭ�e��_���YʙxN���N�2���R�I_5�X��y0�N(g�Ÿ`��QA䡭�����3��c��Bp|w��m y��t������ݖ��~y�9�y���RJ�Rb�N�C����N��[�X�BV�=S�k$8�����<�1�'����a������V���?�����/���)�Dd@�&�/��P���y�����k�r�!Z�z��ì����lޱ�¡��� ��ey�p�yT���H��X���)[��{<�rr�3`�a!�o¦����uT�xB�2�����9X�g :��d�f<˷�.u�Y����ɫ�|�i�(8<
�&����{tʏ�!�7��N#n��`��,��7[�kb>�L�3�U?��1�Q�������?�)��z=6�J����Lnc���0	e�͊=�n^q��$�C	���������5S�z�D���H1�?�@Eru|�u�3��~l2�*��	���Ωh6e��T���!��mg?T'W@w?ן�٨P��N܎��-�7���YO�Q��O���ߗ]���!M.�t�pT>֏���$>�rM�=�E�3u�Ŵ�[C(3�eb��<T���"�T��Ad�rp�$*7J�R��j�
4;��(��'��2�SZ+β����fq��n���n(l����H7(����m� �5:U�{�o����q6  y0z J~ہ3��1Ϲ��r)?�_��	�C�̅�-c�+�Rd�n<�_�峎�<�����<x,��_�oz7M'ثYUɤ�oa��JO@ۃ�I� Q6Ե�q}��2p�4���E`��ˍ7 �s�WX��Zz����SE���ija^l��z�W���M�Y#�X�rl��G��m��<�P��D�\�ީ���wI� 2��_�F� ��0 M����3�Hˉ�o���4@�_��-<0�c�ԲIv�`WI7j��T�m��r83ȡ��3e�E��؋��mߒKݢy���V��щ��r[X)��4�`)&O�Ąǝ@��e�|���94�����Y� �ͱ�D68��*��4�z��n��Ee�&�ti��k���ie����14��`g�6����u��=�R���*r�~t���U���)�Lz8��0�����iP��3�� `]��L�H��Rk+�b���W���q��]_T<J��}/�t%�|{{[-t����~^��}S2zM���~f�Svz�@?r��<�i�oũ^~��sQ�f��:�ګ��Z��jP��d��ߟL�ڠ+k|7��OUA{�8����	��)�J�(u���S\��]�c�ľW��{x\U�xt�G���'1:�m={��_Ngܒ^�ڱ�������%�f��i�IK!������x�{��SR�!f��nq��{��9F��J��j�Ùm(t.��c����Y�C6u�A��aE�1G'��B�
���2�t؀xm#�L]9�l�R�LB
NB�M�E��-	�2>7�f���e���̙�k��&�%�������]��s�s띈;f�:#EA1��v�ޚ@�nN�@�ȁ����a@gY���]��A��ߕ8�5W
ۙvGW2b�W��yR{*w�����c�#����
���8�G�w�k~!	Pm�4�J�g`('�]I"C-[�q5�.1>:�J��F�_�Rë�ҚlN�֬�F�Q�N7��\��������ʺ�����I��*�1xj�x��ϛ��N�������:�I�]���3+2�O�LǞW��A�Ү
�Xw�eKE��yO4h�R��-x�Jt'�J�?�/<�c`�-~)�'bj���c7��&!tO�tr��#\gX�)�Gҧ��'�'���w�j7�������6�c��L�}h���;���$!�ΒM��M�z����y>	h�z��$��]���ǌ�c�N3��L��BU���?�Td�����a7� �;(zsB�x��Κ��QO��a��#���8g�>�Mކ���K.�{g$.��*u��uUR�d(������֓���J:b�b��������'�����]!	)�cu pw1�		��B|���n�>��\���T8��]_�b?�c�E�i��O:!A\W�8�v��-�q�W�X։�ݥ����<2�~�����IT��{��E����*�W�/�h���L��E�zy�颏A�aOrF��%24��;6�q�O�ט�ʥ�?U9��fn淎I����p����w�����[�4Il��z�m�C�q	�y��j�]x��� �uT�V�y7�.Y�$ШK_N����Y�!�#�O;�uJ9W�V����$�OIaŖ=A-�v�`�Ea]7Ӆ��F�#+�kM;��Rl�_��unVy�`��i)�g� ޏ�	�R&��&J\�Z��4�vg���v�e`I��E��:��{�w�UlJ��D]M�'����S�42����h�>+H������z��Ƈ����|�����Bq����+�W]�ВX�4��WF�"A,W��ߞ:���^0��w쮌�*�d7� 	�������h��pT���Wm���X�9�Ӆy�WvL�L�$�-7 �	��
p���J~�-����9�^��d� �U�͚�ɋ��KRE3�f���kȶu����]�e"ڿӦE��f��2����ㇰ)`�ΐL�\�g<D���"8�:'�D����mT�*\a�q���+�9���f����&b��8������u����|���$�t!�����~��nX�e�ѓQ�4�\و�	��\�녻�fY"~�e�~�����U R���_����J�?̄�/s��J����MV'�%��K"�N~�K�F��^�{���r�R���@ނZZi���C){"xץ4ȫ�b�3���;̷lp��{'�OŹ��U7:E����ޑ�O7(�V�͟����X�6�L��S�QWOJ�}�mw�����SW�xo/�j�B-<�-�`���WU�p�4T�K�_���syh��e��R�9+�r�k'z���,rX,�Y��ڛ�]Hj�.q���|Ӛ���%��@O��Xf�?G�J������5ym�VY�������	�uE$kk0m:�.����k-�J�C2����*��B�s/���D`jm<%T�f�#Q���v��_R�	ʡ���@�g3�i���B�GƠ�D<�^��%����[8���������19H24�ѳ�4C��^�?^�����r22�Rz���b� �{�Bz��BG%��C�|�Z�#W_d��X�B��P!�?B��/�Զ�ގ_>Of��c�4�7�9.�H�m�8FH)���&ՆF��g��` L�Zz�IB�����.�c+����j���*�u�����v�pH�A<:�a	ړ3W�� Fx�POľu
��K/@�6�U���G~B��Qb�=�Zd���I���̇n}�~M������V��N�^��"2Y>�tc��+�h��lp�/��'zR�9�lp�3����7S���JU'����Yn�Hh�r?)kx�)�S��Q�4C�:�L:��X�ױQ�^+&}�˷tH�ϲ�@�#�آ�j��,x����m�c6�1�"-�J��$�#-������m���K�~9ŎBVU_���*J5�B�5��V$���⣰��s����1�A��jy6p��h��BkH=��Iy�I��x¥n,�;�dal�@O��w��Ơ�T|��\����e����O=�A6���9O��.p�1a�1q̧���ː���
��q�|K�����r`<��Vg��E������n J\��0-��?�u���np9%�xq:�=�NS֟C�޼{	({K@�8�,�r�G���R~�Q#F��Qv�S��EC �[�H���������kln�+��$� ����UF�q�u/]{��	�g�}�!x��Y�)Yį@��1�y�&�P�:�����ܺ���v&��/��t1���.%�8�q�(�EGfո��)��}��}���oy������^���� ����nx;?�ҳ���|S@�NQ���v���RW� ����.Ȯ�,s�s�@�}v���/y%��x��Rvɢ�V�93��g!l2,�315�q�`,F[����ڹ��d��BH���[7���$�Tw��uNU�g�$��S�\PI(�8��V��o�Nvxɛs.���Z��ʸi+:��i�<k)Qjm�z��ݾ�17p�b��zz�y�����)�x~�V�Sw���>MVFH�B;2T1i"��5��� f�E0kI �>����V��I��7�ۊ9	��Z�Wc��b��Q��#k���1��[xh�F��cs�ou��&����m�.����(�
}�J�D$ֽ��[�Q���z}�I�yQ�&Md)O�Օ�� vV5�¢YT^(A9�Jf�8��ǝ�l�_�r�Os8���5�e�N`�����!v���
��=�p��?�]�Am��1�CĜ��<��n�6�B�oR��/���PN�ü!�,����E�ur��G���������ے
���j��(:��iB�ho�Fm�_���v�������R��O�W��Y�T�����3 	�S��Y�JGf��#�����,�_� ��E��'�x�Ht��{锜��d:����Yf�޸}覊#ي lV��}��Yr�!^$dg$�˯�N��*�H��� C�^�Q�(w�/Y�^�טj�R�#tv�)�=C��o�C�os	���70�:�x���Ms��:�e�>Q�si���nSLR��#��ƞ����A���c|��r��/8�t]l��U�_��̹}la���bc�3=�N�U��IYu��Y���5����&�w7��!򃐒)�ye���	1���p�c�/�7�����v���1a%<��ស��\;̓v��g,��'@�M$=��M􈄿�����o��o��"\.N͑2p�7X���,\����`�aHX)�Z$��OBI08�������#ݝowL����#u~3�hu�k\2N��;^��;�����"�S"���yRe?��N<^$}��b��xi��k{Lw��s+_�5�`y $��Y��C����x��>a�~Z��4h@TGe��u^����@%wB��f���\]�
�Ђm���(���Q?���ްD�Q�^NP����J	��{zn��%�R�3�yKH=�D������~f�¨�e��m	$)[�����@Z���eb�W��uڶ�O����}|�0�Ӆ(��e�M���(�������I�*�y��w�d��r����Ϝ~�)�f~���[�S�H��؁y��>�x��/_�0^"��݃v�Ll���ʞ���x�4��/;�#I��Y;��a3G����� ؝BV�����^���B�_�^[�pm�u��wlotvt�Sy"���k5_Ҋ�0NV�����G�\���}����O5N�Ɨ��TeE�\�;I�� }��Cཛ,|�P��	����0Ȟ����`�W�#
�	
_��*��ΟٳG�9�lE�1���n���L��&��/�W�B�����F�:�?IyH]n�F�O���o�p�*�a%���PO��.�c����a
���t@Ь�y�|�?FjR�綁��tq|��TG��"֪Y��{���(�{5}�#@H�3�t�8�'ٰ$4IF��A �������/pptW�aj�t:y��F�f�gK+�Es:-�C^�dlvZ��џ���M�37
aa���5��T(?y7
�� 8���,�{ߍ��n�V�	�J^����+qY�{�8�n��kF��p$C��rMp��ת@�y�3_�#n ��sG9Ī`���C2P�U��t��ҫ��$_` ��W���`��HCCqK=�a��U�b��U�PxuQ�5U��"�U;�#�0*w��b���Owa+����== H=?���y������M��і5U|�ϗ�XYg���Q���&����m�E+�D���"_"��m#w�����_R�Y����N2�lZ��ʍ�	U�'�F��$�,	!�겁�f �0е�����䴺7�����j�A�vB��/���,l?{N�"#�]O�:�����zƀ<�?v3��Ѓ��LE��6�$j�k�J����^	]���?e/"U*>[І� �+�<�g�)D�,����� Պ9��k��g����}�dŪ&(3*g)~��=k��D��mDҁ[�c����|,BIi�;:/ڗ��R�J�7�:�ܨy�<��הE�W�d��F�rN�	2-cz|9��F'�tO�����3m�?��M�r��}���Ⱦ@i�vޖ���d���F��ה�B7.����n{���thm?> �V�
:,��0��'���k*tc�|�§�d�F�n����є
i*WBm����oҤ��g~��)�E�,>�睳/
�ĝo��}r����#�T��N,o��f�Gy�0���L��S��b�F�ѹ�2�X�� `+?.���������M�m���,���|,x�x9����ܔ���5$x��4��Y��v�ê��t߯Vw$L�P�.w�B� {C�*�+����$ט��+���Q��	$��탥'� ǀ?����-��u=�"��%0�|�b��ػ���ZK>9zF��ܚ����<��1$�M_�h64 �x`��W%���N�1�D���Y@7}�����`!��壜�H1h�j��̱ܮ,� �mM��䛟�����+l��o�!�r2h��z�?�Yc5��KZ��&��Mf-��X'\�^��/9��>l�W2R^�>����șX��i%'���*c�%9��0Ս��,�ߍ��fkH-�ST�u�1��f�οo̦� S���d���3@����)�O�K�'�3��q:�j�	[Ȼ,|q�Z�"/W�oK�(Vr����ͱt΁('���0-:��.��yA%�'��)�ZHh*�K|��-��J�����y�S�)iĊf�x'pi�%0֙SoesN@�I}��%�b��Z4'�ɱ�6����u�M���_��LJ���W��7.���R����.�ʜ�� ��� ��
�7 h4fh�2��2Pf9�I��]YӺ��-���t���hV:�Ʈ�v���0*u
v.w���h�����p�>	�����Ry�Sq�������,%𹊼K��5 #��`��*C$�TG���Ym�.�&~�;YT�;nOpIBY�E�=��a��(�۷�bYbBw[��P�B���=����@rg��Ĺ&��qg��/�����şΡ�~t��3͑��=׮1ԑA�0Q��׊��B�~!�z�:p��R������Y��f�/}f��s�i^�(���ր&�l��| �~�� ��S�	�	o��4&�C��"܀���_��Dj�7|��!e��J�e4L2��:���W)�l�u�jM���Q��5{O�<"e��������B�<�ofZ�u��*$�S�'?�D���A<��ZY��_k	�hϵU����o�Fu�h1�t�!�$��7;�K�ր%'��-��7��O��B�M�5��T)�j��C��t7pP�����7_}L`D�-���63�lK&8�J�gt�PƙmٴH���m��՞"���;=�_z���iOy
��gu=����^�P���D�+�X}�)
ŋ�T贸�>�0�=A&\Ur�fVt��P?��F�|�O�d���G���3�l�3EE�Q�MKp)��H�}1����D��JT�R�\��k�gi:�
3��%��h�w�qx���V�n��w/���C�pޥ�e�� ����b�fUW��ų79��/�+%��m+"g0�z~�>��SB�$4��I�}����W����c�"�c���h�>��5������G� �Pk٘���'5�J�΄��1{��R�0۞��k�y28a��;�˶��Ȥѡ=�@���#9�%�{RR͝�a�΄�;Ff(��d?FT��Վ�j�N��O��߁�C����߀�3��oT<̦_2HI9�#5�f���M͊�Oa	�Z�p:VT"v'�"�+�ꚣx�5v��N���*K�6�]T;V Vx�-G�ھ�C�ﳿ[N;��'��~�vI�⡕kJ��Ca��;��{�ꌹNC�� ��	�Ϣ�*q���h����PB��~���^>�E��K��4<c�>|"aG��q6�,*�}��"�v�0���z4)2���A���c�Á%a�N�,��%�:��$-y��|zX���Q*�5�$?���h���Σb
7{g�7�)��:a�Ԁe���������.C���+gh�G5��3#r-���Y�kI{�r?��$Y�5��U��D���:?+9�E.	�7����X�$_�ԛ��/O��g������2����ƘG��h�}��q��Z��3�ds矇�s%�[^�~�����Ki��o����RODP��$ٛ눌����k�ɜv�)9�tV�^����9�l�iW�I�d)?!4u�͛ͣ�0x���P�^`b/)�Mx���KgpS��zc0�EL�3�Զ�b�-��m�SGG���Ċ���埵�ZK9�4S��;/�O;!ε�$-����4����Jv���З��F�����Z��	R�� -0tۦ�3~��^���2���o�m+P��	��X�9�:��L���Xo��56��uV{���(���T�ލ#&�[_�.h�B��[���B-��d6���m�S��x�Cea9~Yiu�A����~�g�6�����`Μ{K���ǰ;_R�8�QA����:�+x&���2 ��;�oH=m�58M&����TVz��m�|�:��T��S��喻���H��oD�#�C)� �	4ᲦK �*�u���
ҵO�<�f70�"�3s��e�Nm�9l(��s7��rʪ�-0�4���v�z�#5���*�;P:��`�dXPd5LS�&vߺ��x��4&ыm=�%�Q���%��|��O=>l�ENe>�H9C���`;���Y!�ƁS���Q�P׵�9c�/O׉N�x���.�[��#SJ�5����Y�x��E!X�3�3���K@UE�SGW��i0��
1W�AqOXhX>g�]dW�vݬ�F)' ��$�%�Z �*�e(�N��.�S��r��kD6D���'`�ڠ<L���I��Ǹ��Eɷ�w���ArC�����L��,�sA��*?ri��_6$r�B÷͙:�_�ţ���e]ד�i,�NK5���L�
.�|H��*!Zǹ��ꙁ/����K���4�e�V�6�>�ܼ�q��fH��锪�$����V|P첸	�[�[˟c%�r(�3�$&� ����+x#��)i9/�ϼ��m������;m,��� NM��"N�s��u�T5����4��C�I�ZN�V���ç���N�M� �h�fL8�4�i��dht���a�_�K��"���e��uE��~ ��%E1S�}�gV�\��*�2Q�K���}��)f\���'�������������}�W����"�o��[YT����{�O%��������Eg�Ժ _lU��T��r�K��V���*p:���)�1�zB�](^pY	�ڄyn4����Cp<�� �0o��'\R[(�B�	�L��7��1���]��i����6%������e����K�������.��=���V(�ScAf�����0���!{���ě1�9~mXO�,5g��:��`��"�<7���$8�ѵgF��](r�3ޡu`��	Kh|�l�{V��m`^pM��,�e�٘*|�.�BB�z�2�W���JQ�;�26g�z���D�K-���oFy��K �e-b	�������^Olp\g����u�4�?�HR
mt l=���G��G���⡐v�p�6��<Lا�8���h'�78m*�g���h�%���M�{�Vz`�nP���K�F�j�W����dd�ףOu�b��x2%Z���3������8�龍E�0.����5��`U�j�J�լ�.�Y��!��(�Ð ��Z{��u��8���/�E\^ӛ���e�5-��K5�m7�*�*e�OQFfǱ⢄�~!%�C�D$)O�}�ܼ��#ݦx�Ԉ �V�E�^]��=U�3��j1t���a����>!��^�(���ޖ?���Q���|<|�,�)�D��R�Mw&Ixw�X�������q�4��`�#dQ�����$zeB'��^\f^k~�$~���M����O���9�%62@���:*���79~�X��LK\�ۚVRt^����qYXH�NBa�P�~�߷J'���ʤMO:`T>��H0�D���/_@S# ��X6�oїe������m9v)��Ϩ�1?�[��x�{M�b.�Ⱦ�=�,��P�Yс��1�+ۧ\lCƆv$4E��^��f�S�j�9�T�@t2+]:����(	�:�4�\�{��T��]�fp0�21ӷez7c����}}!�l�s\���Z�����
��V��l���u_��7q��uc$��s�k��p��,�qrP$��lt��B�Q�%�o<�ľ;���'����HWZ�[���{���>��]��j�J1"ȶTT~d,뺲�[y�$�⌇@�#����J�|ѩ�H��5W�6��%�Ҿ�˛4$|�9���{����^�� ��|\Q��L��ףgf���{�e�y�]	�o��K�d�g�� =,c
f�'p�!)�i���u\|Z'���TO�u�m|��H;&�7s�`�g�&��Mx�₿�!Q�St&y9`�nظ����9S��fZ�*�1��$n^C�B9����U���rG�z�"��(�	9���o%��w0@�<��ϝ)⮇�D��$y,4{\���Ҧ�.��S>J�4O]���}�)	�g�@
����#y��W�Uu��9�ZE��0�0	�q�,�vs���m��\�_�-�5��(V������9��a��Q��n��8���9I��ˋ��{�w�{��O<<�}駟4�]�Q�C2�d3����ġ����npO�<oEI�^p3k�00�m|�uhtٔ猕��&�����I)�(mZ��|3m=v�+�ȟ����x���,�n��t�W����tϽ󚌿�:}@�B}�Y�#@p�G�5�p�Y�<[
-�c��@��>]�ʋ�l�l����І=bXD�*om%r1��i86��d����� >ug4e���Zd��lȅ���,�0Kɨ
D�	CZ�p)g#���t	UR���>i�ʘ�� I-��o�\Yo�I?�j� g^��Ы�xJ���-�R�+5�˳�r����ݿ8vt�l�/��u=�~�/,����w�VL|ࡐ �R9] �HS_d���jl@�Җ_臒��/�vK,1�h/֡(���г����3J �b�!���Z,3ͭ���t���iJ��w$���<�3�Y����ŀTJ�sf��Й��?��#�Gg�������j�iotk�K�'h�%  �yeJ��|���V����K��fЉuC9ū�ʇ�u$e� Z�^��zigʎ���A��tL���t�Μ��9~/s5�[\|=5��}$�F^!����X�r�F�ź���R�?G�������i��};/����MQ���޸N�^ -��4�
�-H}����!�a`
5H���rK��5mW���t tp��fv[LI	`���`�;�f���G�gB�S@|t3/��!E$'��e7*��A�"ˠ��y�ňiJb��eo��.o�r�P�=��ox%ݧ~��7Mw��=^�q��X�����J�}&�l�6��S���8Eh,m���zZ��U&�l%_�)��� �����huڽz�`R�q���ქ��5jZ1��~��R���QAV������{�Gc��ӴQ  ̝�5e$����n�h�m==$��@��V�n(����PFԫ&�����Z�uI�l�Q"��������WY<⼂ԯJ�8���j4F@��%�����Z��Q�5ld�2д՞�m�h����'U�m�Oybys����ٮ,�(�������D>��'�n>�´��A�>L��azZU~l��Z�lGe[�9�MHzd�D�2�F��B-kn���՚�`�ׂ��h��MUM�����.h���>���� .�Onא�ߤ���`����a��e����[�$&}���(�+Cc���`��O�uQ`�B*k�?��ߚ�$��>Ю�4�}PD-���sJv�j���'U�!fw���p���.^���E� �8U��I` ��E-y�Tڿ+�a�viB#՘�x�^�Y�#J�p�i��X"~�Ǚ���n�� #���O^���(���KGQ�>��t���1���@��%��24y��xѳ:
��,6�8
۹��tő�J��Y9�x$f����@/���o8Q��G*��<o.D��X��a0F�%�_�>�Q ���].EO��ٰ4/�Y-�Ui3�f��L��ϓM�Ca��rf�"0��Y5ป0s	x�D;��	j\����S M:nix����.E!�I/�@Q�3��h���hl8��X?��'�ri4��b�d�l���k�|��3Z�ȽC��u0��}�[��q��x���J��S5���x�s������-�,9�z��<���w���Hǰ�S������1�p�kj�Z<݃�5jG���drY�ߺ�Ż�i�TT�7M����!��W�bt��v5�����}
7�@�8w)�w��-�A��G�9J;�/Sܾ�V�3��x�q?��
q��F�\(�]��\_5��ư9��ִ,%ema�'�n��������6�~Q#�Vʢ��H�Q���2������VEQ��+�0���~WKe�h����4�c�/T�%�a�?��*�D�������b�%4�k�
v��w�j��\�<�%
����Mh'�H�#7�㝽������<�y�7��Ew�YOM�z�5�ԩhv(���BA,E9��V�.��g�6|"`/�~5<~:��Ո� h�>Թ�B��]��8Ԍ�:��+��cEeg*[�qd�!�!�!�X��b��J�{�J=�l��"T>%���x�\ܼvt5F��r�r�~����]��;2Z�k��V�'�$k7`)��x3�d�R˼���t5�%��p�	��r�˓@oz`.��isl���[ ��Ǔ�!��/�{��tKƭ�F�;��`��)�x�m��d�4/4�$A��R���rM@��Ȯ�O��&�&:H�7�%�נg�OF5S�~^����������(d��(T�E|2�b��U��[������y�U]j3���k���X:O���wX�8D�X��uɐ��8��%o��X�tub�^N��$O��>}�=� �i	U��J�J#?lˡV�������2�MA��d�]��\�l4c��7QK0<R�Y���xU��7(��&y	���UA���J�>���ß��=�+�| 5t�l:�k�LŲ�r$�����1�*t�<�]� tN��7����_M��:���j�Ӭ?�E�̗0�t���޹6�XL�U,�~6b�8 S�N9D$�O&���rp����_i�ua�#�����t�HӞNN�MGP���m2�.�d�|���	�������$�.����bV�P���m1qmI���/YL0�!�==,bv�m�\�]��_$�������Bz!���_nU���^
��0��?�E���4��&w�
}�^�����A`J��������[ぬS�vx��^���X�H�st��1��	�hJ�?��˒�}�+WG��og��I��OyT��2�aē�(WS������9z9��%�%�ϸ���=3N�HX�{����v�s־��I+ ѯG��}���y��,�-5�� ,�}5	,0�+Ę1��^P�2�t}�^l�G���˷|�YCa�a{S��aȐӏ��G"�`�`��\����}4U �#��&�dS��%�\dF�g0�H��S�}(��� �L�m��;�{������)|���L�D����������Q`�7ԕ[���Qa�SU�s�	�M�>k���1�%� ��K�4�LJ\|��z4���P���9�~�h�T�Ǿe{�.�	xA�e.%�AS�=�n;�gx�'�����y:����eJ|�U�)	B���p7f��I��l(w�h�p��״�W��M;���"����ty���<�
����'K�qSU�N��7�%y���/1l� ,E4�!.<����io�#&v�^X��f�pNL=s$�����L�akщ�`|��῰A��,���)���턪g���%�s��køXp ����9;ْ�ȥ�a	�$�)Eࡉ��لy� پr��JS6䯾�B51�f~�@vR�fIq&#�<�n&k�O��\w�y�7��Ws�9 �	��~�\�#ތb�S�˛�/&�x�Sj{w�� ��'R%�V�A�`�脌RrƩ��p��=/�ȿ3VP�Xr~��� �G���d�a��9�A�4i{�l�/Kh�elJ}�4#!���hk���+�<Ra]�R���n��љKq��:�XZVhC&����2=��+��%���l(���,�W��tO�Sx������K�?��ڦ�j�N����g��e}Gh!6��)m��V藮� >)BZeq��?u/7�%��.A�}�;���Կ� '�.uOӅJ�@�`t�{L �ȡS�������C=��M��]���B�)b`+q>z�?|d4�j�!�2�{��,L�}�:}�]��]#�!X��:��U6�w[T�o�/��h���4�T�x��/������=����L���X� /N����Ro�Jy��p�qi���	���5Xu�Y��1
�4��b��l圕��H�X���~'ÝeW��b���t�rE��F�1����H�oC
:
2]ŵ{ ��X�AM����EE���݄z�d��M���̼]����	�^�:㹛��vE���[* �F��m�|�dl�+���B���v��O8:]F�Iey�1`�q@� mu�E�����W�+}s��#�G �ĵ_��i�$�p�L��V+��H�c�oX�F����"퉊q��B�K:^�.�!߀5cK�r3�鹘�l�cy�p�Z5�H҆�à}�T!{�o����^���]�Xwq8R��4�vд���>4�� �?K*53]�Y�$O���t�Ƞ'�y�TU��\�V��1��������%8���+�e�~,]1q����Ⱦ��ֱֲWD��^o���O��#�����1��/������ɴ��<���u�`��-@_W�x�����w���Gb���i����*/r����um
Ї�z�$���G'�\` >Gx8�^�_pY�5���3�]SN��V)��U*�$��}��P�.*ym�P��7YA,Ӛ!��v�1��`�v-�l����:����V�&ը���Q�?|��aoYs��������6���]kk��١xX'������@��^���K�$~�\��������3Ml���=J�=�(��vD��_�����j-Q���d�����;�$�1b驆B{D���H���u���FQ/s��(Y�n��?�yh�I��.����{
�{�	�R��xjWT9]l@��9��b7����L�a�:Ҏ�� j��#0�v�w^&��2��/�N=1~^��-`*��<	A�����
�4��t@��p�:�*oW	�a0Yiu���5�}
�R���߄�r�zR|�3��o�5��(-��v��N�!L��U	�r-���UQ�"jv���jS@�����7'iW�6�^�"֗8&M6������M�1�bha%�;�Y(��FQ���yxW
�� ��p�����7qG3�����,��*���.��b�&a���@&1t��`�a�	�P�ٟ�+tr�n��Q�xґF���_ǈלcn޶������gvTu�e���c�T�u=`�0�����+�v�����g����aԪ&r�B]
G�C��?�-�.�4�nȖ܂>G�Y�k~�?T��������������.��;��:�ZF�yj������~���^�&ϸgiZj�ŵr�[���Q=�]���l�79B���Ǥ��;U������I�!K'(�Q«��)�A.f#�'��SfH%�}���!�+݅�Sk�r/F�@ubO�1hv�๶z=�it��N+���ZA��P�	6�MTN=�4U�D���_9@_�⦑o)���cYTmK� ~�0�B�H��Ä�,�6�tnn=Ј9��)�,�!���OM�6�83N�O�|�`K/�_�S���T��li�߉'0�~uH�Q�`s�a_�&rQ]�ۻ���4i�E�����}/d�<a��[�v�#^�y�Iv�i7w�nͰ��Y���Z�
O��y �(�$��9EVUfa�/�l�eC;�)M/���U�I��0�=�o��N��!���xې�����Ð�0��?�Au�H�8���ԁ�]\��� �َ�ܽ�~�}����\����c�<����X�q1e\�fi�up�Dg��(�}��lCC1���ܵ����lZ_7W�tP93g��uo�b���N368��,W�Ҳԡ����S�i�+
��qZ8P�3F\�w�v��.F֋��[`K8�A(�!F��6��4CI�o�>���u��G����;Rv��x&�(lvLI�Q�:�.�\Y�;IkJ�/�c5\/  �X��V�Eɳ���i1���տ�	
hd�i���������8��&PO+���C�\R(� �V -"���|��4�;�x�ezdV�� ��m�M��{��J������[k�J�ٶcBp��?ixY�+�\�5s��ǉ�xbWYk���������f>(��xpz	d����iu�A�}݃���H�P���eF�Z|�	��b�V�ZKK�ċ2c��_)D�>6�-~��R(��g�/����~:(��1���"�g�:J����}��^:Hv[�^C�#�B��8v|:4{����X8	�9�y˃�1r>Y�\k^䫵�f�W��Z~J��:�H-���,���h�!�θ�uS�LS���x�9�a�p�U ��a�vP��ǘo����w<=C�c���ڪ����%)�O��\3V)^k�u�V���e�=�����Z��<�k<���(e��w���a�M�^wQ$l7\EYaN83}m0E��z�����<o3NR�P�D��|��c��fWI��s}��/oۊ\E$Z��o�ܸO6!�&��%������H�C#�������,EG��������nȂ/!W�SjR{�o�=p�AŁ������I�𷶏AQLS���B��f���E�C	���6O�pjeC�H=|�}	u��Y��3{�w���q:Q��#�`�f��C��E^�Ʀ*�=ȷIQ^�]����hʤ����8f%�$���#Ay��z1�^��R���v�*ǻ�_�����u�'���hxt�` ��F����=�C����f��x���rN�B_��V���gb�'AO�1��d9�WE���X��j�j��*{\i�?~����F,������Ȉ�W����!f��?E�UV#��s�;�9�d��O��.:�d<0��Nn����saE����'�i�u�%[����4�����pR#�c���/�b)����?�ƚ�q 2GZSj���M�=���{�T��^�>�n�p�1w̸����(x�8�^2�&�b�9w�qW ��!�������4���e"�m��0+1-'�9�)S���G��A�Q}�3f'� ��e���!��㸧^:l�!��8n�B�u��3r�r�Xі/��
丹Puℙ���/�8j�
��H)!$F��{:ᒸ�������'�ʓY��p����	��q���Тƻ�~�dړ��l�ڲ�ҵ�rz�"�rFx�i�!�ץ�����w��.���"�0 *.O�P���
	������ױ)��!
n�ap�N��-<%A-b�#B![������3_8��2I��� 5��:q�D##ח�U ��D��~w��!�p$�����Rd��8�s�Q��})������^G�IHᠻ��I]��
��5��r��z�����Fg���O-�큰ˇ��m����jtN5�a���&�H���VRnők�N?�/�fk��9�>)�k�yŗU����A�OCK�H�7���;!���<���F�b��D�N[F9�<����a$z���kJ��X�R�|ּu��|�wDm���:�D`���ҕ.�JE��i�M�Wb�bh��q�7�p��Jn�Y�e@���X�;�XB�i;�P!��x�[��+����@=?�6��S��P0-����
8�h(�"Cn5O��֗��k�4b�+ 帲��3\TB�3,T\�䙫x1����p5N�ZUk( a�$i'+^���`���@��p*�����S&^Sc]���>s���a�o�3��z?�Yd`�-��ڰ�P* �hGp1{æ��c��!��u��;Zxy¢I��Y��Ľ���;<��G���N�r��K�x�ڜ=�=�����P�i��D��UC���7�%9F�*�sUS��n�ݞ[<�d}�KVŠ95zuD��u����e~�i�'�	�ĳ�ȁ`A�^Ԝ����b6y`�:�mrË���G�������x>U{9�(�x����)z��B	�.6V���)�'�r ��}����{�@�!�#�k��p!+���8��~S����rP���)���.��dhBJ�<c�������U��J�4s:���+���+�x�&`�򺉞8W]�j���9��R��6��,%IY��%�N����$�QK�D�ȼ�c���L�)���F&k|��YZL���M���@bB�=��8n��+*�}���m�Rpf	J@�d��h<�=����^X}�H��<Ȝz�]+��/�u.By,8݆҇r^��3NYuA�Hx�RGg��ߌ�&��
s�~fq�Rr����KS$WM��́2!��S$H���7��jp0R���Y&��B�!EB��´茨���磬�R�e��Qq��T,�ӠS#O(�Óp�������Y��s]���"�x:��d�c�O5����p
�%9	(�d8�<�� dJN-K��}�����|��W�>�魕ug�s�m���G���*UZ����>g�*+\��[�7$ֿ��\���t�#�ϩ�����f�k�S�(&8�����!˺���r�cq���l�y��KU��0�&9n9��8�("��+�_dwG��-ۧZ��ҝ^��հ?�9B�E�!�>N�a�X(e�Xe5R�/�@ɀ	>�.��Dcؙ����KU"��
�e���V�6��L$ !����!�m��pH�z��f��ָ+������^9�x�����x�n�-�G5�)�&�C��ѿs�M[U��n�-+��|��B��S^���r�o�/�r��\���ϔ�c�b�69#�q}=�Jџl��� ��Z�y���f�+E��~������զI����]����3�GvB�Q&�p�(���Ku�k�s(�ގ�	��	����t�W�5[���K���V�yt>��RB
��c`) ��
Nr��t��f���@�Z-��(f|�^�T���^n��a�l#�;4��Ov)N�&���3eh��D=!
�$���,�+��-� {:x��li�כ费H���Pصͥ����S�+w���(Wte��4*���2@Aɐ�)%ӱ�]�VoL�co���J+�G�+�~a�6�L�mC��t����ɌyV8����lx�>�U����������=G'�8':�-�R�N��w�#"+�{�H���v��J+��a�����0�L�<�6)��|�?��jׯ0g�	��>Ν�+�/�܄�ȯ�mM��Ҕ�Ϊ� ����Tu�����[l>��v�j�@.���gTKg�q�r�=���/�'��l�C�m����7.h���K���1zb�Mh���ݼi!��m��������nN[�ʁ�~�$�J�B����f�v�ǣέH�w����yf���51Xߓ�?j��J)�x+T6�g���!gUoj��.s����<��V+�����m���V�LA�T.uD�|��
�V/)1�iw����\r��J&q/�䵙X���'nQ)@H�NpR�.Yƾ��:n�9+Ќ����y��iZ���]^(�}_l�#_�Ҹ�Bg�`��W�ri+9�v`x�h����Z���S� �����%���k]���)��8�tk�J\.+� ������{b3#ZŪ�m�	6HK��
�#��}�2w!�����B���Y�����j�ˈ���a>��>�W���ٯ���3c�!E�C�^���'p5�|�p{H'cؽ�&�v׷�d��2�H�RD��Yo$d��3iX��s�U���������)4� �ʞ�hؔ�J�K�"�'�V8����8-�͘2E�B�Jd,AyDމD�W#�n�z���H��ң�K"6A��J�$��O������hUR���2���\qdVt9�2~G)L����sXY�7G��̦�u��"����y�G�#��e�N���6�`1�f����6+��;ťk���`?�S]���o�}�Q����`}/O2h�5slOdb3��H�:'N�P���N&�$�X��J��Mj.��Œ!���$����t�����r�ɭ�8��|p�_M��C��)YY���$�˖���T�6QJ�&�B��٤���u��}:LX;����^�"�ʔ��$�c�N=;�Lk����QW�Zj�*��a�gZh��	D(��഍��p�g�j�W�E3�+;�D�K}�co�Y�Ң;Y����8�f=���.t�g��L�y�?۳�'XL����%�l���|Wǟ��M���ݩo�t˝�*�j�> ���t�*	���,�C�s���o&I��`�DzJ�$����33�0��<�7�q;��:2��g����]H��A�C�*R��g� �aM�;
��^`��������6*��A��G�0�8@=���Ӂ���d(\�������
5��q��9�>vJ#]j���5�����l���a��)d�m�y�Wl��J�P�we�R���줯ʉk]��Z��摺���P,���`hV�Nm����^�‖�ݍ�w�T�=�ʔ���nb5c̣-~���p�,0��q��hNc�O��'���[�zV�>����c�n�'��FG���� �2T%�V��T�F�,F%u����(*(�Q�:hO��}d�H ��K�,���xf�]������$=o0�F]����}��&�=��<8��J���"VȘ�O�Z�2}~���=�t{"\Z1�Q�̟�c�Aa'����ng�OM�#�ֿ���p��է�'0�.6[��'t�=e�`I�Ż��)�(���0Zf赢x�li޺���q��5R"�����<�l����K*�4�9=��iL!���	�x��m� �x���W.�3�K�^�|�BW����i��WٲyNk^�س�3�>�w@��1���<=R�=.�����Eu�c&�c�Gv��hfs��	�K���u���o[-�)-w��H�ʚcT&��-��7��1?��$������|:̽R�_]�֟1�K~�X�e|0<ع+`�kl�R8�6M<�����O���U�'l���*D��2�21b�
&OuT�sh�q^E���r�K��n4LjbR���M����g�>�C1��"W4���'k7�;�Kjh����|EA)��[Z�M��vω�� �{"/yރ�Ę�W����)y��^Rf�I�獋\/jLd�}`Qe�D�(r/��
?�3�$�%��V�E`w�� �\��v���'峿��e�����OogK���#Z�1K�S�NT��೼$b܋�,J�1�����=�~���`e\����˅���`+�=�i��������4Wٹ����6K��r4�L�0��X%M�6	�~��%��}錐*\*�lځ�_�I�]ZO���Σ;L�j�'wJb��i�r�M٘"t]K�'Č|@g��k�@Y�|(��'r~�k���.�D���[-6��jeD=�MK���8M�R}_�:�*���V��Q�Y%B� ��o$���q�@�a����9�4WU��u+;�(� �����
S���t������wK^nV���:X?#�|R��),}r!��ï�zϪ,&�]�9��&J!|4VDS�Z�)��NҘ�=�Ɣ$��5���a��$�5{�t\m�)nbPu-�y>>�#_C�����f�����k<� F]&�A���Q��ʙ��������Ď���h`��ju�Hv@��������OS�2�U����WM��]�P-���7��%I�ϖ��c�n�c��B�� O'֗�@u"��(u~#���U4���4b�6��`���X�u���J�6FxoQ���4&�%��X��mgU�獒��DV˚��mH�I�;�2���+�0�W�gPs��z@ghq�ѕ�7��1��q5�!*7��D[���{�����JF�NK3]�%�1�_�ڙ�ܾ.��tr�ohj�{�P����F�
��
�XS�/q7C�#�(� ��]���xN�: �ͫ�	u�ݺ���;C��'���G�3�Y��-��T�$�p��16�_�O�gBa��� 9]��h���KW<����R��k`>�L�X�6pM_�>yK�qn;�5�ǖ5�%;�{���]��/��YL�]?�{bm���m+�ܐ�wb>C��5�a%E-Hѱ��§pu/J��/Eæh���L�/���̳��DNQT+v��]ksC��P�Tm�T�V�Z�.i�W5LRx��̡�'Ǝ!��O]u��%qs��`iw�e�ɨ����=cʚ��G��(�kB��i�U4�<G�v��*�P�PD����Q�k��ᑒ6t�6�T�T��e<�ۭ�-g�/�pڢ���|\�i�O�
�_}zp�eЦ�L���80�1��j�{»�.� J�R[X���ߋXV++�z[̋��T��7}�m�!�$G�ۀW,U�vg]OqBp�r���2���oX��4�^]�=:��9N��V���%�2�L7�.����À{���ã�s�r(	aV��d���ؕ�y%b%��[#n��Ӑn�'���l��z�3Ǵ��`�}w-R(����^?� 9\�)G�ǰPn�P C$�ӷ�iGR7�Mb�_ۑ�� B�j1�n8�%�H�9+u�L����Ŏ�K�\~���K�M��5[����<S�[Ѻf
ԩ5P6	�g�VmB�KϠ��	�4=�2f��c��n�gW�2�c�	��?r��	O
�8J&����:�PlC�Q�Z�1��=!�j����^^L����"@ž�/#�������1a����"��{9�ږY����M�_�`���t-�t%G�����J}P�f����_xh�b�xN �ݕ��(�ˀ*�ni%�0�3� RM_��)�f�����a�/:�Z�4̨�b�9Դ*n, �nWWH{�Fo��J���*ԅ~z�� 9�nX�*�z�J����gsj���0h��&,��c�|P��$Ν���ꊡ�5Tr.��f�u���;�p��F�E���q�|��mǽ�C�8����-o�����H|f�/�9o~uqX��ロ����Yk�3,Mʙ-�v���{w�W���H�"{�i�_���lFh�?�j��R��6U�2��=��_�Մ�	��F�op'xiP� z<�`~�z�O�	�_��uC��>�R:K@/�K�>�!f����t��&������R%���@��Ymo�- ���X$v�=�1E���L�����-���e��B9��d��%9t�N���� 9�Z�bGM��?;Y�P��Km;����_�ͣ��^~��_!:�t��z�,�J�DY�y.�`G���|�w�ݒ��ir�)�!n+7f$�}D譑QX��۶��lG�W�����Ƒ`����7§T�ݸ�-��GD �����tmS���
�9I�(]���] �M�
��Ժ]�3K�h�a�e'��J����L�BY��Z�ˊV��,���:���Re�U
�i*D�L��b�IN��������G(����B�F^�J��^����'╶
B�I`�wBx�+2�,�é;�ᪧ�b��?�Eo7��#�~N����7W	Ǘ��D�ZR�3gxȢ=�e�h��,���iM��o�$:�QS�&e��2�h�/{U.�ᯞ��*���_�;<�|S�2�9� X���*�}D��+��3��Y�VMPm4-�h�F���/�H��ݭ�coP �\İ �@��@��P�[�<�N+p\��B�4��cA�ٳ,�����O7���T�2E�DQl��y�v�ɡ�ǿq�A��0ә�Þ|�FE�T1��j���Ҡ�(]���0�?������g���k�
#�gM�����^[���K�;���l��V�ia)7T�%�}��0xk�~�t�c�y������)��3�S7����M3;��!�?�\^a��k��,@Ͼ��'_�gg�\b�U'��c�R��{�:����m�	��X(�k;c���[�����e3ג��Q�$#�s2(��	���X��fȫ�ݍ�I���H��F:��F> ]�򜵚ci���i�w�z��uox�C�O��m&����V|�um�;��믶Dx�gM�t+���GXv̼�o{��u��HіS`ڕC��p&�%�^��L��U�#��.��i5�f�����$��i�����#p�Wk1�̈́�v2��8�a��4����kf E��<�kx'(��5,�?��4ɽ�"�ϐ� "Sߧ��EqLOk��M���w-Ϧ��!��L�*�n{�NQ�m�R��^D���4��J���nGvT���F���`�����"�o�w�K�k-J|{�%_��DU´��-y��QYG�#@�%��E�]�$)��$u���/�Z���k�w��+�j�����0{�*�5�g���B�wŇ�3'7G��j��['6���H����'�~�٥М����P7���8ai?�J�-�'�����Je�s�Z�$�*�W�WQ쥍��5Fl��a��F��p�	��a��BW3�j����X�Ry0'[A`�rR�2f�E�������\[/��=U~�x?�n2��sgO[ԉ��g�k*S-ƌy� ���k���4�4���	i�}-V�v/�_R��7�O��u�m�����9�pr�����y�O
֍�y�B�Y�fm�&�E�4���C[؆23�!Vj�����_/�z��� �M
c�o9�����<��)��G�]'EV�s@	1FO�и[��ʼM��i]���	, �*H־��H&��N���{۲��SD���J�s�3$'Uo�6�Ňj��v�:uֆ�\�J��n����Bi7z�nO+.��ך��s�#�����lM�GZ}hьf���X(��/��$}��i1fx!H�Y�`����G����M.��_�&|�f^���ݔ�Z�x:gx]�hAE�SC�R(D��F��׿v:�i�+J�Ɍ�)��O��%)�?�-�^m��A���n�>q�wŜ�w�F�2WŪ��g���� B8p�0utĒ��'"�;TT��N/ �Vy�L���o�.��-C��-�}��|V�Ks�\��?B�}�PPl�N����%��ӂ�z�EP��ji��2��J0�%gK1׿����Hs�r�wT���$�r3��=��՟5��ڢy��we��[�d6*	0��xƁ�ǒ�MO�d��a��*+}}�+j�_��*G��掭��y�>�9 ��+��a�i���D�m��7T�#��׀��)���9�;,��o}�]D�6�ܳ�9Y�Ox;�Ľ�3f��y�������;�u���8�
�y]N�U�Lb ��J�=���޲h\݊&7�I��ߏ���I��s�y����.H��?K�i�)c��M80�����K����6������Ae�A� z�T<��g)�I��=�����T�6����^�.���h�l�/�d���*���4��k�__�ѐ�F^�t��
k�h<�%�Ľ5�L|D��������%��t� �9���Z
�B�u�e�ϒy-���Z|�<YER`��$�zZ�s*7���I����_[��+�����V�M6XR������j�"�Ϲ+~ƍU�ղ�ɩ 9�����6?�x�6��	�+ʶ�%zB��Wzq��K�eE'Z"�4�BP\'%H!�y�I�gt����:����2�Є�/c�@��c���Z��g�\Y�((��"�t����A<�ش��f�����O���P�ms��<.��:���&V��H���m��x��Lvʃ�CJ����9)���(�B�K��_��y��z�J����d{y8�S�)"!��/=uD `>�)a����u���POʗ�A��EaIxS�W������הՂ4<��bk��h�XaK��a�û������.�y�Z�:5c�2�����
�fiOĕ�쾟�F7�*{|~PB��K���g�<WeE���������M�Ж���R�]��-���2G���*�h�h`����Eh� ����sM���oD��G]��cF��24��עK�~�O������}�G�Od�����c������챳$��*`�/-:�JW��l�q\�*���u��]®T4��՛��(.��D\c��(��Sv�,�;;|?����D�����۔�2v:����
��3 [��9$�8
7M6�T�Gi@0ȑ��o�ag8aTvc���fnxK^����BZ,h�x�`J���(���8���i�4� �%��6��ҸU?�G������<��d��3�b������;;,�1
��YC�H��-,��z5�rE	ֱ&����Tr��%1Hs\zDk��I�؞>&�����>����K
eXĞ��T����}������y֑ӪPQs�yY�`��\)m���h>����S��;6�+���7?��Y���b6�vu�_3F��?�({��H�lKĵ��uk�I'�#U��1�X�D���y���K�$�cY��f$�#�_��£|��Y��
)"��x��zYa�R���>[��������V+r���S� �/I՛z]kV�X�US%5e�0�c~�)G�#��|`�h�-��Ai�Y{��G��1�-��<y>J�F�d�0��	����=,'��fGדvh|(0ҞVHطE�s�������#n�Y���3���Q�G�������vЇ%�	 ��L5$���2�-��P:�ʢǮ �h=�`�*��Rs�77&n��Z����p��NNfJd������V/@d����|9����V�Dh��1x���\S_)"��b�B��x'S�!G �	�b{`�l�#�^�q����EH�v��q�eϙ%l��7Hh��5 �N"|v�w䠕���;���>w�(��t���5]��X�̵9�5d���
��G�83	5��ի��7(�'������g��nw����,��I$,��tݑ3�U��U�ef]|��ǀ�&q_r�m��8�>f��q�p�]vA���zPm߮�L��7��s�L�\�B��G��]��AI���i�֓����J;sͫ�)H�S��Dk�6[^�J�p5�BL>Y�!�P�f//r(��t��;*�wOW���/;�� ���d�נoE2�*�*���7�83F�	$���p���m��E����08gl6�1慱v��k�Đ}��H��S�e��g<}�N6�H(|��P_j��b�L�%~+h�T�g�,��d�挻�ޣ���@3�ִ���������X���wqUtjr���Z5���Vt^��;�����'Έ>�w�k�ج�$mY��yrHv�Ѫ5���I�.��lJ��ŵ��XϹ������]��B��:��a�H�gē�YvyRʞA�BS�sA�RL۝,vTcw/�l�3�̆<�H�8#Ǣd��5�e�E�fG�6�p��Dk�@�Dg4�LeqU:��Ͳ�.��Y��۝_ȵ��9"0��~��%�c˰���~�t+��<���Q"����4*�l��T][3�l�7�\�K�+N�d�Z;�+t>&�wu�7S��V��T�[cQ���H5bc\p3��vz��N��rc���9�sSk�M	w��P���"p��Gk�02k�d�����]j��z��ϗsM�!mEwB&���= ^�Q�B��\�o�1^��z�~����zs�k����E �y{C��� ���M]�U�����Q3��N�����{�*�Z��	A/�`#,E��*
��s�X{}n���%tܣ��c�KYŔ�Am,rlf¢�wܒwy}��=�P7D�����:�< ��&�M��JTQ5�I<���#HAd��L.^����jȾ�;Q]Г�X���ۇ+��4��W֫�e������%���*�G�n\9�r^ڮ�Ω��Q����}!��-���_%8c� ˁJcDۤ0���QSf��P����?�/��J	ʲ� ��%o�z[�|�<����B5��A�,lV5~��sG����̼��4\�����{�g����2�p�*�S�&����=-;{Y��D9(�Q�P���Ԟ�j�u���9����>��Pŋg�|��9��]|p�va�@�� G��\��qj��X�
���(��C�@�H�[EC��Th�$�z4�S��<�c�9���f�s�i_�5� c�q�fv͖kuͻ�P��J��a��r_��3'�iOh��#�v�4�\��mP�>�Mf�&4�?���b����!��\�-Ώ�5 �*C��py���͉f�	�oJU�<�U�[S����d�k���fc�,�U��oN��KQZ7�~�oj�5^�6��+���MM�Z\� ޱ)�m���`�9�L�^���
��V�$H���m�m�Ot>v
���ݺ���{@Er�*D2ݬ�NCb�eZ�6
C��=z�qk^��r�뷊�9�W�g:�	-�۠�D�)�� #�66Ue��]��X	xi��JԙQA���R�᭚���Vu�h6!�?�x4lڬemvFϞ|.
�&p�3����e��P�d�ͤ��W
�qC����T��6t��F�I��XG4�:?{�sT�5�s�_孍g}̗��Z3�����f��#|u<$��xش� 1wg��|��&8rXT����oANx��@���jj��}�+�7�[x:Kq�(�j�:@��P��@�{-�h�~)�����`��ٞa�:vn��ߋ �뱏ϸ��I�㯜�8ǄvQ���`�޾Y�~N���TDȽ����,�@\�(���~ʠA�7��sv��['�K�ە��!�pDp�b.�Y$�~${V�a��>P.�{��-�<���z1����WQ�=oP���g�����z4�c=����L����l���Fj����0V�y��T�<Xk'���7�(Xq8���]W���{�X+�יGň�&%��Լ��n�i\)�,���5�Ɋ=���b�S;�:e� �]i������&�N����ƏZҟ$Ԩ�����t�y �vdnU�F�4��ױ��g���G��x����s�x&�ޛ�u����SV�;�wp�N�*$���~"x�σ�2�G��f�B�N���yu��=���h�*�������E��� ��b�:\�CP>��+W'��J-��9�^�Ѫ�۫ՉNק]Z�p��uK<�1����^��5k(G63TaE܊�E��� +��&�ϓ����g�[C;ծ��)��V��8D�ыM�('/w`p<���#�&*�Ï.�*
�j�k��X���]3������TD�?�1z�g�� ���i�:S��w��cE�-��2�HU��`Ʌ&��Z�O��}��qjȑ�C8���ހ�h�e)m�%�v��E�e�J.�������.�.&�yS"+|{
��Q_����a�҃w�I�
����#�,�&PD]�bp]iS�) c1�y�x�|~B�~��Q&M�Cá@=�pi<Q���l�|��rD��V��js"wu��U��YHް�{s(H�
,��fy�}�닲�*����<�̃NO�s�W����+��ʶ�aF�U��\�]��p[Ճ9�1���a[�7^��7*��)���Q;�Y�)[�	����P����n�t��ѻ�4,�Ǩ���D������ȗ�|�>�汀"�I����P7�ސF9KJ�!#R�0J�KC�k�zM�"���g*�Z&���mUC����i��C9ʩ����/"�&����.q+��ک�:S�x��pV���4pE�^� ����uY�i�Sa�� JUK%�`0��}*��r��'1� �rE߰��_��K'l�Q�7��2��GH�Z�:�u]7X�ӰG7d� D�7G�J��	��C�x���d���j>����b��ny�nd㸜L��(�l���:��-m�dݧ}�����^3S�:2����~�<�3y�`P]���Q:�+.Ng	<�sw��V/_{�l

�P�
�Dޙ�  �C3�z�le�s��Ω�+$�����%�e?E��p����%Oܬ��)�섵���$��,"���Ĝ)&+�ő$Ǿ�\x���O6`]��E5�y(m#�g���A'���������a7���xh�� ?^z�y	��UU����q�x���#���L^]����&sg��q5>Ӛ%U���BTBr�^����"��X�K�ws|�L2�Ŝ��$k����>P��%=eT) � �jH���b$?�Q��&\kr�k �,f<f���W+L�F����Ŵ*@b*�W����E�AD�B�	rM��E�Q!AY��m�0-,45�f���;$V"����J��p0X�28�'��lm�KU��hS������{�m�oD�JU��[on�S�<�LN�u\وO$�j	t*���-��4��e��>����6��Jִ!��O}G���(�<S%�{J0r��k+7\J~�}���R��[�	Y_�Ϛ����p��ƀ�$���?t��n@t���giN�Ų�G�%Pf��L!��#�~|��B��J��3�,	�x ��a�3a��	{?�	u�������'k�{I��o��a���Z_��-PU�� 4��y���ɭS�`K˼*�Ʊ�R�
ȕ�S6P�Y�l�]�@&4�Y��#$�*����Ѡe
L�j�N�޷R~ћcL�-��0�S��P���Vc��h�:��n�4P���e�G��@p�z��o��1Y��� �v���/��O���v_��ͧ�L,b��Y�C��/����U�@�������R�g��$�FFJb���ާm�p��@X�"�U�ƫ��o���A�����(��kԶН�p����Uc �֐��Ň`�*8�zn�Gk�;ѣ��j$ڎ���
E�v���m}sC[:�-ɦ�����ꌴZ;�����os{��1���5[Fjv�gIC����P�w�y�Z�nc(��E��l�*��rh�`u�.�#6�5]y8�1��w�C䭢!%$�@+��@���h�r�ˈ��l���aQ�U5v(��X`B���EEɫ�cx�x�D^�@��<
�g��'r~!���?�U S�/O^���SX���EΊ%-���i@��aܣJ[���wH�P�B�K��Jﾀ�_�y��8����JtY��j�{���t�gd�bQq�D��wa�n�Yz�ڎGK����X"��������U�Ll^����rZyE����
�����N���G�R����J-��{�7L@>��2�#=n��Ɯ]�$.�Z�dl�5��X6˒��t��(�]B����u��E]3fw��9��7r�]�@;�PKC͆VC�<GRP�2�T�!a�i?:�
/�y��H۷SL�ߑg��Q�i��hk��l_%A�й�睩q��]0^���!�sYZ�������X��P�6�D{�u3�;`_�����Rz{��*7�TUskF�Bј8xt����Ri��+?tW|'�bV@��^��(���g6A��+Ϯ�i$6^�$) �1xC~q�DE�ɓ�;fX������ޠ
����0j-�O4��!{�1/4sx㶄}؈�#q6�@��Ђg�4*.�2Q@����Àۀ���bkQ{�����&PLr�)6[v���l,�� )�gT%���.��V��H�B�ə�!�\�#Y���<��+����<��&e3G���<f+���#��E�K�B���A))!�%���[kn��7�/{M��R�vƅD�&4�z�|��3�����<WH闼����eJ���C͐�)��Ν�w����*��t/
fuf.bO�a4v�o�\��M���j3�駾	�(�`*��!z;��$?l"�7W����|a>\6���7���s�>��Z�@q)�>z�*���{��Y���u~h�c��H܉�6�m�����O���ϓ�n��~j{IwOt"�Dg,a��öܬ����%?"����!���@��V�ģ�q3�����h���-硂 �6��^X^�5��W�׎-6u`V�#H����5H�*3��1^�a��"���/��x	e�D�)�񐠊~���^�R���V3hF��Yt��FǗZ_��9A�/J7���i���v�<�9`��ܴ8�H��&-|M!$��ZJQ�k;lk0�a��� ����ݭ娨c`�Ōk+��=9x(�������D!k�64jj����-ZD�����%�è����o���v�pr싋��#�)9��l3�pl�5��h��(����a��%3ۺ>�2W��ϳB1���
qp��2����o4ђ0g741���r_p>�5sW�s���ڏf���Pa�$��j$�Ӊ���::�Ϡ�%����s���[B"o�����������և�Hxf�;�2���S�&�8X�+.#�R[��C؍a�#�n`�O��!eޓ�=����Z*w��ȕ�%o�dg���|�L�Iۻpcj�k69�G.�F��� r���j��˓�5mh��N�us�m{��V�Re�=���q�@cD���|S�+�=�OZ��������#J�����&|�~zD[��[�BS5�A؍^&�5�g�ĪF�e��N��.)#��-T���qdr�t�o:\��v�|qY7����h��gH��@���)�q�f_/ ?���g�7J�&����0/� �#[�����u�N���V���XN4���¹DO�VF�FY�}�F
�IPMS�)ah�
�1�9����[Z��x���RwOR�~��T�7	=��@T�g�.%�t&�a��@|�7�H�����b���0(�)`�3#Z%�}�Ƕ��ugR�ف�j�9�565�Iݮu�a�L�ϺP/��3k��N�[1���Y�r�030��[���oʃK�Le���Fƨz�)�L�:�>z��^����gKseg-b���}M�����V7�<�A��l{S��H8��Y!���À�56��G�9^d������sŀ/Cd���I�q*��9�`�:��з�V�7vb1���a`���`.D�k�w�+x�P�;�R�s�b
*սǐ3ܘVb/�t�P�J��n�B��A�x|���VKeN�@�f_�� 
'B,,,��R��0�����H]��x`�k��#�B��c"@	4
�y��~xq������0e*vQ�K Β��%S����)�Kk�a]���a��0P9WJ]�P���Ȧ��[Oc�.-a��&�:�Bf=)"���-����Pxtb�kΚ7XȆ�h�2�˨�3'��w�������r���ݓ���=<l�<��!7�6�,����phd�<�'�ў�N~�� �ؗ۷<��1�� ��`��t�V����Z���x�h�N�ÑU|�ܞ�ťcx�)��������^ ���kč^�&��s
y����P�hv%��$��^�"�bye�׃�����yٺ�s��/-A�y�ݱ�a���H$���\����'ȋ���=���t��n�{㓹zx w{g�dh�`����E���y�����E���Q����Z��O:�
�r�A�M��(�$e���	�#��wO2�rȼ��E�	�'���G�%�Zt�nx��J��y�����%�.e8/��"ѥ��+!��N'R-��!,��XH���PcXw����l�̭���.�`쾢z�)��z�I��-+����Y��1;�w�@���E�m$���H��M�4W-��� ��ɪ�q����d#>1��9�F�����s�U���=D�h���W�\� ��N4��1/������"���[�	����'~���]n�y�q��60םv�>�pm�;G]-�J����m�@|�(����G��ޕ}�ux�������J
�F��8��ۃc]�b5qo�y=S��l���
�Z����iZˆa�ؒ���
�d �i7
+0j���n�U*�IG�m�^�ɡq���c��(<�Ž�V%�K�gmU�_	��kˠ�Ƒ�V&��%��49z"Z�K�=gBX~/�	�h�6�˘��(ۓ8V��M��|j���9g���'�R#��YbN��@�#�L��]8>���`�W8+nS7� �8����0���z��Ur�ct����"�x����c!<�J�H.������k��+='�Zx��$�����eA�֦�(4�V9u�����e^� �RwqyRh��ǅT��U�Y ��y�(P�B���)���-�q��1@i
&5 (7i���hR��]#����Vӂ6����q*:�^j�x�"��a��
��g8����la������x��i�%*��P���%'��8$�bϒ��%ÞH!��>D!Π�1��6=�.L�gH;��XQ)����Jd��Vɘj�3�Um� ��:osr&�K������$�:*��"|,�Q�j�K�&v�$Q��b����F���r}��5o�O�������!�U�@������u��Y@0�f�ɲl���:�����]�懯�`�,5�
�%���H,t�M�
��4EgG��GD��|g3��]��\-R����>��P��q�D�~�C��HuAK	ǹ)�>\^G��(З����}2	M�GF�RL���0�ά�kJV)��-��pt(�1�Ŗ��:ܽ����l���7{��2�Q{��q����
Q
b{���pN1�M0�-�,W��f��K8W�-'s�@|~;��	�ΌE���V���o꬞�	�9)g?�S�������Y&e����l���8�2��%�����4v��t�C�Vy��b�omJ6�(?�%�k2��W�#� )9l�R�r[�@�X�pT0]P׵�V7���2�|�B^K����R%!/�=��7�6�C�D�>�M�;&At�%�d��ڍF�+�lB�4%�O�
���}�La����c��s�	u�fi;��Es�|�&�z�-#�LCLJ��zǺA>Y���O	1���CY 
���`�.ܖ�RS�s�<��P_*b�l6�Gԫ�����@�bU.��>���a������I�U~ե�b��~(T� k��uN���$�A�fO�&���V�f��3��Nd �Y����N&E�A$��Pn�f�1��~����iH�s6~~NߧFZ���i=�8厩�ė]B�ב�y�R89a=k�;iTx8#{@����lE��XA�M��qHX b�t}4` 
p�d�8醿��ԅ-�kɰmض
��|nt�7˻��b�#�T�u� n9�GV��#f0mY4�
ӭ.|��_ËM�さ'lI<��'��) ��4���*�J#'���~,��L�mS�̵w��=��eD<t_i�2yr��V�(�.�����=�!)�!�ٰ�>B�`���|�'�l�&{�%�zћ����<՛�Bé~�cۇJ�'��4V7Me�c���:��@�S��(2�~�J?�i�	��I�%����LT65 ��>e�0�(�����7�ˮqvE�oTOJ��$3�L�Ч���97eb;� �PC�R��{�����bX�@_��g�� �Z~D��j�ل����e�F���>��m�a'׺d��w9�EQ�"�I������ ���ݑ;Z⠽���P�L�ݖ^��M�:�O�(���j�c�7EvLֿ�ȧ%��5D9�z`})�u�޽l�
W��D��n���&�枯�v)���;|�J���[���7N�� �AQ������H��qKT���)��V ��O�Z�ہіjC�g���
ٰ���P��8�!�ײ6L��3��Ӥ�|"q@ev ����8�CҢ%�Uc�Ws6%>6�����,w��U�	�,c������eaV<�am���0�������96�b9ʖ��Lw-�
��M��2<+�FORH��k��f/0煦`�V�h ��K�6oα9��A�+-D�����'�,fM��.���MВ���.�1א��5}
u��w��M<��34��2kP����56��n\�φ�d��#���q���1~��?gئG�'P�s� <�a��F��˯f�sf����Znc�ݪn�~
��v�zqG0�n��^e���BLjj� _������΂,�;ǚKt% ������rx�6'0�TU��$�O�6(�Xȇ!�>�u�I顚�dV��3���|G����@I�\��� ;��*lLzI>r������w��� �z���T�mພ}wNs6p�p��+w���pڌ�;C��O��4H�0x��J�vj���+նl�g�����w- v��Lm�������.�E�#y�:��wF4����E?8m�j�Ǡ}n�:��^��]<��Ǝ��z9�IXI.�i��<ŞA��¡f�Oӵ��f��ɴ���U!��_z���ݭO��y�g��
����7V�RP���Wv��HDtŭ%'��+�A�׃��d�8��6�f�L0�<�)C,<����͂l����g���,���r}�4爺5�Z�u�~��=-=״���%����,�f;���^�>1��V�o��?��2�}]׳%�����R���s�>PK�%�H�l2�>n�D�r̹�z�#q��M���bƙ�[��:Q�Wӑ5Nլ�n��3���|?a�P�K���_s_������哩p�Z�,�Uh�r�J֢ggR�4w/OS��zdڛ��c�ΙD���ҥZ�f'C����d&n����0t�i���1�wP��ޱ�D��·T1�Y���6N�����I/W��;$?UN��{��a��-f����M�bj�,�N�����QUxIZ����e��o��j��!P�AG�; �(ъ�$�?-��!Pq�i%/�&^d��g6,�o�e+fw��u��x�2�&�y����l�~%C���+ƣ�9F�J(��`A�z�R�z�"b$y�+\%2i�5�CV#��r�J���y �>�/��:�T�AW1�v��XDYW�x��oukXV�p4H���n�j,�<�z���㵧�٘�x2��7-F�*�&Jcw�5쳼)��=N��:�g��� ��h:����Z5�"b<^�ݜĴB��2Z���ߕ���}{2��̯��x����U��h��x=J=�-�M��E3���\��\j\%&�{#�c<3�$�m6��&�k���{б��)6��	�u��N������;�0V�0U�j��+�i��s|��a��a�F	���B#.��Iږ��@�ɽ�b{��J1��YG�T�BD��\����4=��8"�IC���Ή�`����S�MWӴ�?�,��6�h������	�7��mӑ��M��0�D}"�0�F;��YgR�H��1��ʭ�}���C�'�}�e�xդ�l\b)6���v+�߄�����k�Ҳ9��wu��������ÑJ@�͛�)%�������88r|��_͉5K�M �iAp�u� 6P��T�Z�-c��.0�x�K�J�ӷyS	��i֗GI��˩�t�	i��~%@P-���jb�]?qf�Ɨ��<�/ҽ�OԈ�)͈�f� �I�]�Bg�U�;���c�͛��Sϝ�rIʧ(U��nG����# 2��D��A���{�#�x@����Y��jI{�I�G����I~�y�ÿ��TT[��@�"��c,�e�a�ޭV,�aAAGγ�.�r���g��:��&s�NA�8�PH�.��R�eߢv�����7CT2_5��Që�Ѱ�G���{8|�������E�4��s%�ۼ����1�g���ּ��W�'T<����JO#�-iwp�5jo��&��z���ba��ܼ��, iP��xPK��yѮa�	���Z��r���,ς��;V,�:M�\�R��` %m��N��YÜ�0�L?,��RoZV^�M����I=^b:B�ϐ��S���zzm2o���;��W��&�����Ͱ���#�$�Cx�6�����h���pAI�����?��k����w�#���,0U� ���׊`���ǈ� ��5�>*FlR��]�"�x�i�=`u/t��E+��K(LՖ��EY���T�gb��:jS�J�O5L�&"�NQ?�4E�`Fa�]KeEbm����\� �]�I�2�0���7�j6E����u%x.mqp�DM;5�\
ͭ���'�l��~�0��f�cu�i�HL\����8Ӂ�h��h��R�k�昼9/�'�]D��g�/�+R�e���ip?15�!�q��I2D�dh9��}��$�LǗۦ�����ʴ��H+��(���Q���+ME@G������Uجܲ�e��X�p?�+���7m���KnŤ���8u;^��r�F�m���9���F",i�"�k�7Is����L�{ȝdd�$Z%���.�tl��0�H�=]=�XS�����$����F�:�OP�Lz�8�.�-r^w��Tu�'i�w	��� ���Nx�ÑdV\�	�E����u2T�)1���ڔ�>yj��
���>�D&��Wa���pVʐ���T�DE׈�!��hc��|B��hHB�h���� *u�⤬.�;j���A�fV��[ 9M6���,�4���g=��V��D��E�:Pv&X�N�vƹ���Kr�;=�#[$h���A8c�����i�2���b�|� 8>���J��;g:L��l�4ISƑ%`�:��l�T��re����U'#��IC�����)�!�IaDc�Yd�@��Z�r1�S�눴;�o�W1�{�&�/ q�şɻ,:�	�Q?D�2�
���)�����o��Z�۳����'�ߊ��F\^Ua���CW�fX����7͖Shz����1i����!^�w�X=��*��w/�KBԁ�Rc*[Ex���0c�q�Q�36�W��b-ѕo�3���9�H,�@�c}'�R�{�A�i#����YUo���� ?Tql�i<����cxDw�K�֌Ӭt�H�of)�U�/��4J�[i�B{�4Y�c�"������-�f�h���O��1�XF��r?K������5[(:�߂{�F'>Hh ��M[n/�vf[�̝i����|�q�q������0���A!>\o��G���XA'͗�Bf����X��	�\��$�eF�̈��M�$5>LB�:D�LX�����3 jA4��?f��oR���0�=��Y���z>��"�����)֪��j�����9�2C9ęgP���r�rJ�t/2��9#�n4b�x����³�m3*�|Y.Bp��[�v����@?�~��7vO�s����Jz�;=�#����k��H���m.6�y[��b�R��W��Lx��$�! �.��S�"Q��M�G"���=M�x�bg��d�%P���9���x�c�6�#���=�q&��$�`z.�G���z�l�2E���Sy5���d,K��E����ͫXZ!��خr����ОuQwc�HM���֡��)�-�����V+���8o�y�;Ĝ2��>�>�vi�N�3jA��
����֑�	j����l���Bi�l���H= �+�LJ�b[�d��x�kP�Y��4n;N�~E���)AH�s�h���I��
���U���*����D�c�\�tP�.})P� �"�"{_��	Z����WH@���Ń��ΐׇLpY�m�T@ Pu��S��NL�t<����X)���)X�7��:b�T���T�!K���&�w�:���z4KH'� �W����g޾��,%����Zб,�Q3k�omP)�*�����M�
D)���l�0g�#k�}�?��� ^��� `�:���Z�h<��哺�+��y��c��R�fS�D�{n���VWh�������Zz/,� a��ƾ�u�{`ئ�Dv�����XGm�����v�ܮ���J�5��wЗ	�c?<N$�y�?��7�0H������m��T�+�G�ɤJ��9��s�&f/�G� S�� �y��D����;@�H���CJ��H�Ӹ�s�e�KQ���`���Bf�!� ��7m}�ӽ�ܵ_Mh4$@$� q�2W%�C{��h]>��B�X��fAǭ���*
�)�ܣ��||���jj���&��s�Ep��B�L:�Z�z�,<^���6c[��e?"�ہ�'�F��b�/OclX�2�S׏�G�[ƙR�,���}B*eD=��Wʿ�Sl�,���s��-��;�3 jJC<b�#���b{��"�*�"\��,�t:�Q=
|�;Wl��e�8�,�c��T_(!��CV�ꩆ~�~�qbOa�#�"��
�X���~����D�f6F�*����ڛ���rk���'�_���#�6��Ǣ�����
gUBJ��kȂ03����#�^,S�,_r��`�#
����R��ee�cz6���zf	k	�ܣ��Xg�t^�y��d�$��e����=^%���H��x���U���Lz��ń84$��q!<ƙ>��D��Ĩ�F`��w|�ohM�KN�-7-yhU�5u��������1��ܰ�|ނo���N �v���Ɂ�o]ۛƦ%f����Ja
j��Hc4�h�;'��mk����b|���Al�7�ݥ��MW���v����S��K�jGJ���U'd��})z!&��]c�iH��]V��2�|�t����x%i���ڻO�j�H~�fg�'>��Z�Zû}&z���9ސ$cܾÈi�\�;{��3j8mg������c�`��g�V�Ff�6ua���f9�)�%	��6��cǁ�eN\6����� �e+J��������?�MODP�=��ښf�%��m�Uŕ�Q��iZ���N�7�$�J#�X>*u	��b2/�:t o>���l����fe�3oW�l�b	*��c&W����� M���*b<���*�L�,P2�����<	a?e+E_��6\�\�%��IL���L)%2��*��Nyq�ˌ�H:�����GL���(<����ǳ�/��U�v
�<7�׷}oV�>��z���EΨN�R׾��!bj�Da�7$Pو���"!<-�/'7����p���)���\��s��u�7��=��!1�5���«yC-^�=���3l���S�0��zL�x�i��?}�%sbv���F�Eos'a�On�0�^��� �C@��L�p�XN����%�վz{1Y��]�w�Ӌ5�"�s=��;k�Q��W��C3[�F/#0h�Y�e���z|S�|Ri�qḥ�Uh��r%������d�����p�ܸ�c�6�����5�t��\2J���G�Է������9��%��J���	��l��R&��}Dʏ���-�}�M�zB�xʀR�B�	toY,��ob�L>hT����#a��bh��n�`2Y#�pp�,�9I!�,\Ǔ�_װ��rzp��v��}�������6q�����d��d�����%����<�sn��A:�	1R�������9._�i;>�R���^���lM�̡)n�+n[D��f@�����t�0�Q�YS$c2_�etp[ 67��#��F���SY�W��#n)E{�%�Oż����O��#a6�/O�c���qX���CQQe� ����r���qR�H1����1}O� ߿����-ò2'��^�gT}c'I�fjA�f��Y��afu��[d{�3��ݓ?S��0wj�z62�
`�C������Hl���90�v�Fי^�iנ��Ef�O�t��2�I��z�e?�G��ݟ��宿׾1n=U�c4�b1Пo��nZx�?�<�InЙ���F�2�E�J#p[t����]��A�~H���i@/ޱB��/�O�Z<��5�&��y�f/5e��Q�mԙ�ɲc�;�ų�S]�鸨mt�jCy�����x;�䶯%��Ny��v?RO��f*�,�l1�ת�Kx�V�|�v*ٴ�iw�X��@�QM�Ӧ��.|�B�x�j�2߽<f���Ϩ]��H�e��O��c��w�O���|�J3b��^V�s��?[��y��P�qq� �/�Uo��(�n9B��0�,�eOϺ�ֶ��msx�K��iT8�H�i�s���e��C7�ʥd����c�c_+F
;9����U�9܁+_<Qy��x�t@�SB�#�2�(c���|	�)�&�R:H�
��y�%d2?��J�!A�H5��	52�w����;7lEOBSbٙ��]�K[FYȍ�e���^��R��g��x.m�ڀ�7���Q[b��O9����:<�3�@y�='U=�S�cF|{�]@�~貞����X�~��^�Ɨ1�·�2�^�r;?id�FDA=s��B ��#����S�1"L;�@�L ��&�Ԥ�M3���H���;� �9SE$[������zV���T�n
k˼�.
�� �"�+��krIo���FpN��~�����$�xE\�q�M�>�X�~��1ˌ�,�^��!y::��o[q��o�QN��,Oݫe[�띀NLM�d���ڂ��"�|F�f�/�?mt���޹@�|���O��Y'���f���
�^�i�=u%d)P)��=pN���w721��i��$�=�aYDTE��>��d�}SAT9�Sk��y�;�C���q(�b+��7�}��iT���C	�%k^�x��	�,�RG7	���^�@�f�a�8�)f* `"�E8��ב>��KPa��8!���?���o�Wt!u�,����Sd8U���l^R�m���%��x�F��o���
�_]��Lo؊�R�HY+��C���FM3&ULQEԲ�5{R�X������֎ۀ�G�/���09ִ0�i�nqY/���JM�8m܆���-.l�����}6J����@@X�>S�>m�	��R㾧J�3���7�lZctw�{X+����x\��'uys��l��#�堆4�D��kD�c�0x���X��bm)���V%�����J�8�����#\�Q�M ��V�>{���*ū�j�V���'�jn:��C<�tw�>`A�=vf|��K�r�

�����7[OP�w�*�G��r�������ԅ����S�(r��FUc}���W(,?��~%H!բi�lt�Q�M̌$�����=N4_ۇ�oL�K��j�x�L>o3qR��j��R�\�ʮ]���7���IQ\d��7�WG�!����?T.za�&�������ˌ�m>C�q�d6z�#�Hs&k+���iga�z��LV`��u��� ��71���
����w�JB&�O���t5���M��"�#�.:	 آQ��r��!�[�Pu�I�\��!�����]��Vsa�Ÿ�A��e�V�R0>� �D�W�n��ձ]{�TzV\lg�g��KR,�#�C>��Z�NeVꟿ/HZ����HԴ��A��w��\(m���P�w� ٤�r?�dR�V��n���j�Inȏ~���ٲ��5�_a�#��O��dP�Ţ@�~ZB7=����@v���r�؟�I�虫�ؾ��Ko��q�b����������#'�nzC���{��_�5��l��W��x"�豎�26LN�m`�3����W���WO�7y�(� ��)��"�B�G&C[{a��j�����W����S�ͥ��?{��so�#�hB�B:b����|������S���P��� @��)c��:���0!q�_��3=����C�.���s֑�������������;MT�35�C����Q�f���Pk�_�ڸ�&d��	g`��	�5�/�!�nj�Ѱ>�8u瑱��0��6&���ǎ��<bn��W�h�v�j�о1&���9�����@�J%����(�Iԫci��;]�