��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��E����$nz p�D�mM� n��eR�7u�w�֕���>�s!���C�@�!������id�_Yd8��)DIl�
7�+J�)�[�;�Դ4;3t	m����E���mp<�:��9��]�L8��g�[�x͗��cr�5�~�c�t�3�mr���W��B�pb�m���[����GC$�������Ɯ+�Cu${#��I�v.&�{L��
$ƚ�q)�\���xz2_����J�-p����h����^�?��+��C*�r*2t$h�����m��zM���\��0B^z�!�7?���4>�
QH����ωw��leo���a���C�8t9:��Z�`��Ԥ�=X-w�h�ޱdU�k*�>��W��A@��DS�{�#�]�d����HMb�8�d�~�9���)b1"#w!��ք̫�8�k��@x(�ʧA7e\��Sf6}p������W�
���](o�z�B�놲^Kƕ��~��KPM�*�������tD�sU��N`
>OHzF]o���N0z��ɚ� /p�TTy�6}�-5h�~��v!�[4 �?^ �WO/�2�7Jd�F��`��/�/x���A��&�@�[����|[~5d,<���8��kt�@����%���^����R���/?:B�z�6��q�4��GN.H�:��qj ]V�~�`J��?9�������c�\v�*c�y��{�b��LX���� ����F��p�C��ĭktQ�'�X�2�/%�ݹrJ��$�����Zu�M)�P���wACJ"�G�l�ΐJ=���~Z�ѶdО�;Z�X��ߗ��$h�Ԇ�ֵm�`�����K�L����'"WXW�X��ƴ��7�P�o��m�����!��l�M
��~͇T�����$q$]�������j��+�* 	<h�G5�U+p=�}n4Bo]��
]�2AZ�!My��f_���≾�ٶP���[�i��0Ԑ^XB:�X.�@��&��ިȇ=|��=�dC���p{�@��O����Y��p4�K���S��C ��*�Ј�¬��7�	Z9�Jۚ�`�}ǩ`nW�xH��TMr��� ��#A���͆s?��jB-NNcmØ�[���w�̼u-MZE>f}?�}�_��4��Z����M�a�Sg!x�_�J%���v��=����^+yg��,�$?H{�O$k�w�_#Va?��m�m�`{��O�e�B�7�C��h�����KH$�0̚�\:�9lq<sF���S�%�q��N�����L?������X��S���:l�0�Ld�j�-���|A\,J��2���i0B�8џ3��#�)����X������贷}E�z�$��HEALƈ.5�,�a0���:�LdK�ɷG4#u��X�56����t񬍔y����Q��]Y��˂� �3�('˸��zD\�3}>L�|�۽��Q,�����/x/m&sK��W�.yPdH�C�_��
�<��r}��Ҝ��V� �h{.O�L^$���Y∠x�д�����/��G���lH���	��1����͎�$��lj��d@��~��I+�j5�oGh��z�Ռ*��d$Ԋ��J!�С�{��h@�?��;b)�:�����FPk�F����2 ���I�H���'<ُf^����G-��!�s�.��A�^��
YD��Z���X��S�"��A��
�=���m��G���3�{�:�
���\�>2�!�.����c��<���u]�M*t3ZG�GǏ�B��~�B�z�ڸھ�Mn4;������J����)�����5^��=,\�n��,I���5��7h�mڅt�.�Z����5Ya��h��&���x���f��8��.b��҃��zw;�qg5����1l�*�h[����]��V�T����bB���?�
�?~�܈��i��9��V����J�V�B�b7�c�hy`����Dw5�+՘�����Q?�	�bx����L��;�K�º~�"r)x�M��j����D�[V�w���"�������ґ��oӖ; ��2	�u��\�=�r���c��䆔��W���:��	�t롡������h��@'�񄨛>x�#���L��J�듫��RL��l�f��C�V�4�϶X�
:o�t n�Ym.oޔ1rO�k;��i2��:��6�M)T�K�=�����&�ۮF<�zJ��wG϶J}n�KBOCI�&�a;�Q�	Y �!U���R����4ak.b�'���1���lx�����������X1!����!��`P��T��V���L�UM�uEd�+_D L��k�?������%���N��}E������D�mV(�X�F�cI�D�Y�����x?"sz���|2!�`�=�@t���+�^wE
�c��|���N�d��9�(�"~@��+Dq%�`"<�������[N������Ե�����]\i�p���0N4r���%WRSBDD��v�����<�Q�GîV��tO٠���bZaV�Pcp�X^ƿ
z"kk��J �IO:_����ɝ�},*���HMn�kΙ^��T[xW�xQ&se�O���Z�I�б�>�Ԯ�t�!@��r/��g�h�[�K�z��hJt�����t	M�E�a��"�᧽i�IM�Wz���གྷS���u�#񕞧D���ż��cZ��汯�̞��6�Q�z*��,�����r�	d��0���E�lO{]ȁ[�5��Zﯼ4? �_�K.;6�����=<8_��sh�!�7`r3e����vOB�J�$U�UV�T��� ��f�%�Z���+���r�!c����i1��V�=�b����X�_�~���� ��>P)�JSZ)�	Lq�����"�$9�^��I
���5�Ҽ�4�C���7;�l�JEB;K�U"�v�qR���)vC�B�a���¡9�t������SsN��V�Xݿ��ߠ�:���\>R�`�S�-�����k���K6t
�;���-��'wJVx���g�h�~W���?s��(o����k.L����ed�,h��#�A�J�<̩d)L�r�{�0NA��eҬ�{+�JD�����S8EӜ�E*��C߄W�l��(7����}gG�m	֦C�ړT�Q��f~�n��={��8�E�&D&�y���1�˼ȇtփ�#k�Ì
/��h�&���-6�O����:C�9��wHO���mJ��c��s�aDH� �q#Hj^S:}r�D�r&ItO��P`��1���_(�#h�=_�z���%J��o"ty���U��Ї��d�zw���N� ҏ�j-�PP���/�Z�H�XyG�o���F�r&�,�'�I�)#M,�b*c��:e�FD�
�;ĵ$!?4��qAVŤz��>{����p�|�4���5��ӌ5+��>�1���s�/�PxWs}�˿���	�6�_K�����`阰��6����&fja���;�yjQ�6R͈���s�f��b���O��e���j¦-h��i���o�������.i�=T ����N�zbh�:Q�ʽ}-�{u���=�78�����C�$�\��D�����qlĻ�s�Q�2�4�'�Ŕ�����4z@�MY��"R�YN��L�o�e�HvR�I�6�Ϻ�`>�<v8���Vm���`Fv�������y��V�<#���q&�J��x��	JO"�B��g�w;�N�d��:|Þ4��>"��{Ir��&�� L���E>���"(Nj�;ԡm�e�$��׃��T��]\�W6k`��C��>,ܒ"�9��G_��D�ڮ{�WU��k��]�Fi�����{�Jݱq�^=/��)d>�R����-Cn�fG�a��^5_����C7�Ew�S9$���Qs�o|�s����"���bёvޛXM >b��/��q�5���JQb�#8�<g���g}�Kp4�p���'��k��'���j��4�v��)�Nؘ�.4���SH����?���J��u��rƻ�eQ I��͂�D��dB�2��l1�=�{��F��	�=��_���cB�8��MѰ���W� E|��0� |���^B�i��W��:ϸ�n{���Q8$>3��o�}x�w���>#6��u�9���T�]�^�.�&�[���rɳ�y௏�g�g�^:y*��<����+.:G���Ԣ릌.����(�6.���u'�f2���t�ϥ흉P	7Нm/�@�'��&��.Q0�_GY����f��IO��v�T!�1�)�����)�U���8Hg��A_���oW�U�
�f�I@�q�ɥ��M�SX����nY��D� :L����ϽE�\̹�ԹT�h�r��{a	&&�D�m�oL{v�F�^�IE毡'ť�_lƭ�<���,�$1��h����D_����8Sv!q��9���x��`�W�����_�xvϮ��|�0��J�ٻ0��h��;��vBX��g��T�_��p�� l��<̔�[ ��$����8���8
���i�r��:Q*��D>��u�㴌���j��W�s�wxK�W����\~r*M4-O]l��~-�c���aL�G��諭z��l���C����p���1��Ro_��b�6�Ww\����������tt����R(��u�3����������E��+'@�ا�I�,�m��5n���{֜I^IA�$` ~>�')���0F���=
�L��O�X`����]����iMm�v�h;C��`�c�u��r�����0�����kC�ﮈ�0h��$�s�
�2d���`��r����|Un�`v�Pz�!`��4���F�N�_�_��Ǫ�hM`2`�̪:��<�~�`S�_�\ f�;��桫=��/ɉCՀ���&f���|[�-�K����x�"ߋ�2y.�h}��G�m����t^Ҭ�/$��y��j�x�k�����5��M"ݠ	��w���C��	ZB��y"��u Эⲕ�Ry����O�����������Ծ�j��L�3���l@Y��໌�5.6�	��^�;�bn����ND�|c������ݤO�v��Z�`\�eERt:����g=���ՔC�f�3L�Y|Cz^�
T�hL�uh�ڇ�V��6'S��'A��w��N!xm51�H6^J�><�e��˹��㴂)�:G��J�����rz���``�!���t�7'�n����ԭ]��*ԜW,��(���UAN��D{22IbX�ȗ�ax�e��)����0V�@鑻;�A���ߋn����6�G� h>B�	�����_���|&�M���6�r�t�H�L@���A��p���#�7lw��Bқ~�zR�Ќ�B��S����/��-h���0.���eK��l��;`�5�{�\���"h�M��l�hM��eJ&qƟ�E�Yn���7�.�WU>����=�{qca�C���!��mwO����+����H6'6�hœSu��)�y ���_�7��؜�v\;�l��ǯn�*�d�[��x�����J
O�$��z�狘�5L����I�UsEJc�>ׂ�)U(�e?��9�Qx�G�扶ߴH���AFz�DS�Q$�r��C�(��W���	�؏��ͦ�YB?������bY��^�y�Ց}߸ml��t�6T�f�����k�wz@���JLT�{ /�����N��Zؠ��q���2~��	�ͧ���3d�v����+��T��z~�`�m��fa�)�A�7h[
s��д����9B�����O��uj7��1����s1�]��s��rc�C�6c���Z]z���7�1#��x��0Z6�p��u�V��R�}���2������=��ΐ��u�9�`�v��Uqz��P7jZ>�¤�J�D�H�bݐp��ψ=�r-�Ƥ��	�
/����V��6t��\�=���}q��YzD?c!G�Lyi���t_�d���X�Sε�9	-��UB���_ĉd)u��P�-O�S�D`�]�n7��co�C�y%��	�e�z��GJB���jC�uu���{���e�mw���j<)]~�5��F�^�$3=ed�llUb�p�1�����$�=�i$-Z���)KU������w�L�����K�$Y����� oI�~BC���v�7��"��
,R�p��A��|��y�����yv��Q.t4ގd�GН�O�6�$	�����|�UP��=gӃ�$�㐑��sYg��G0!�'�  ��0Ljy���$�&fe�:�n�(�8����� �]�0�&^�܀�Fr]#�����D�	fg�02��|V[R��ȑ� �I4k~���i�N�X�G>5}�3l
4�z���^쨅�+�i��4�\j���2��/�"�e���(fT�cd�r��(}��C�D�=ȭ�Qq"�+��J���ʿ,3w����V���p�:��w�:Sm M(����Z�ɕ�I�<���%|W=�y(�-�8�k�
�9.vJ\q"��B5�}%S�,:R��	�.9Zm�)�]0��j"	5�D�.���{��!��ˉM��d�ڦ�L(bBo�ƚ� �8����C#;�H�	&^�a������A ��\�8�����
�}�b��|c��]�7 °�h�P/]�ʿn��Q������
F_@%4`-�?������gB+ӛ��'��g��J�<1��B���ּP��jrY��n~�r���}Q8��h�<�bǿ��(�X�cGYJ�P�C�,8�`�?�0�;�2~R�v�!6���|����}�`�?,K�%Y$��l(��7Xw#�Υ�0f�z挖s]���(�5&��3!C$�N�`���Iw����&�t�o<��MI2?���u��P`|�xZ��8!�r5cH���g�L�9~k���KM[菒*v �ė�2$y�=1����bU��j�T�c������e����-r�>e����?8� >��/'�Z��[/�Otx(Y�E�ւ�a�G�̀������Y�+/�׫��M<�4ю�]e�Z��Jf�üR�; \����z��#��aH��TU�(Y��C�#�x3��[�]c�F�Q�L�	�e8��.s�_^���.��0�`�rSN��z�1`�tX��y���$y��^8�g��x Ϙ0��x���֐A5� 2��`���̂:���hҰ: p\cF��>����=)���^,.��伕+̪�UZ�%lFU��&R�1�:*��/����`�x}�I�m���9��' [�EX�K���w��}Q��Ue�n��pw��U�ؗ ��ɻ����7�S+X̧I1�5YaCǋ�=�
KM��=f%��D�#��m��l`r���n*(rj���Q�!�K��~��[U�q��2eC-Y�7�\��F��+j��m<v�j�:��rͷ�h�9*3\Q�j*� �aД~O�-���؈b���(T�;���-Yt0;�:�6������eƤ����n:�����9aN�ym���V�7x�EV�B3��y��Xὑ�:� �9S��&���l�:�A�����/��C7�/^��/�߽m�BS�9ej�0��ژ�؂(��#�{���+4�cW�iT~���@W��4�h�W6�ae:�i�o��e�	 ]�5p���[Mp��;�.�9�"� �A���ǉ!�,c1+�g|�P�(��@ĺyG��|�?���2?�س��y��@�6Q՜�:b��ƶ���%�es0,ؔ�CiZ؄ᶆbX����ъ��%\���4��%�,�`/�y�V[2Ms���umf���? �"��M�(�;��dCTt+:<7o���\���;�[P�xL���Zs��%W��*�:ܾ'(��g��N��j%�����Ԑ�(a��o�%�f��\#w�(Ѵeh�y)���P���6��K�=_���*Ɵ�{� ����Ȱ߾@Y^N=�REv
z��&��m��4���-��D6J��Ut`Vb�>�L��v%3<�kC�}�q�*�.>cڒ���>�lFU_���	QЛq,���U ;=��D4�}M[i�.HVI��O?q�D}av��><u�yO�uN�\#j��f�{&��%�rʣ�ZՎ�cGj�f��*�c�'K�ر��Xܖ铠�{W*�V����@뉞Y�����2j0VZ$:�*�h��"1�Kҫ �P��`�ocڈ�*�4%�<܈�A���� �/�c��������V��Ww��P_+��4 ����t��%cn�i����-��tq�R62���)%�7��cҜ��>�`�D]9$������"W|�Sg�VK���QyW�m:]�4 R9����G}�N����烱�P(#%�=bx�GR@	���3#L���%/
���{>�ؗ��j�Q��j�[=�����o�r"����f?�mVJ��TC�:ۊ򠐟�U�e����<|h��A.KC�(�M_D�X����D�Ѹr>U����˲N�C�����e @�!�X���� t�ɡ^�.v�AGQKT"��!���BI�1�����䐍n�n@� K\��8��9����
�"6�B��ђ�f$��g������q%���->;��̨;�0y��DG���x������B�7��0{*0�,R��&G�a�h��k{L�Lh��nJ��IG��14ؗ"�9=�2�p����T�e��|?�xF��40�Z�s���i��Sj~����^`֭���e(~rK@�fP�(��)ʆnnN�DGf�L�Z�P��@���Ee���W;Ēa������_\�/E΂ۥY������Ļ�5����fF|`=�h2�W̪,~�aY��=ʁ�0�?��f*�ܥ�>?.�T*!����p������ 3��.�9�/��~v�U��>��,W���㔥�Fϐl��R�P��z$���K����*���'��
I����H�}�Ųnw��`���6�����|r^�e�K���9���B��XF��U��������v�(:���>C1��)`��3_n�">Mc�a��AW�P�^�L9/+��>U= �����F)JX�X�H6�TLϥx�k[cgt��?7Z�p_u7ˑ&LDK%��lJ�q�𤝖ϻ�&��Cf���
�8��H�,����~f���>D����jsK5�'�@�����RN|_��4��6'�33�фN������!� O��Ljֹ݆�q��ȋ�!mY��K&V�����%��-ºŋ���ь��@F��Yqe��;�d��=u����(Z HS�,�H�1#���njr�Lʋd��N��%o·:)�Y��"=�t����l��LO�!�������̚p�֯��ҋG�Pa���IЁǍ|Ut����F�����s�����8��6ix\#%G��H�.�萐&u�[��x\?����feU���1��ƥ�Gu��#�z�D����k{���p����	>��Q3������j&^��5�I�^R�:V�G���y�)�g&JM�7ct�������|���ۏ�JKΨ���-a�s���_�m����'�!��T;Ht�S�Qr��Ϟ�Uř{���?vħ�IgO\�C[=�����@���ڂP�Ω쳭^ǱHw�F
��x����2kWߖ\�`SPw9h�C�>��B~�ty��*��}����9e�����A���Xw�͆\��K=75�Y�ݝ�$�L���X�rw92��{�$�X;�R�9��,�މ:3M�w�En ��0X�ٻ��fD�L�bh'��Cs�n���b�e8��yo={�g/�Ŗc�H�����}�JM��F
Nx�O9���RU��� 5M�u<�=���;�G��!���pyh�����p����e!�uX�@��y�X�������W$��4���&�_豝��2���y�"�bq\��I�Mڏ��t��-v�
j=�P�L�����-��G��,�p'����(1h�ģ�b��b��G؞� �'	������)�����ÙK/��	��4�Sx����l��jC�i3$[9���(�����4ԉ% ì���W����ɴ΋˖����),��E���::�� =7�����=�Sa)�y��ܑŁ�[�f,�e2T� ���͋�������UM.:��OЂ�W҃�Ǜx�:(�~�].?x��u4-i���^��u��u-9y�_�HI?�c���z4^y�K ��C������v��=�r�?�]��~���b�?;�"�U�ic��B�t��Ѕ�Ƃ��<F�}����R�&HHI�=z|cD���V"�Ϯ�rF�Q�z����PAh�/�>��h��8��@g a9WMxO�I'������X�O]��2_�f�CA�V�q���-��D�]�N����C��W��t�:�:��p\^݊�I���0fX�iD�S1�Ee���+3Vͳ8��ޱ?9��[)�c�8��9���r��s�M�����#t'M�B[�Rq�ojGê���3����9V�K^^L&'��$ݧ�U�9^Ã�����&ҋFa�0(��k��q�f�	���302��@�)w������~D���0��>�5��u|�ɰ�3��&��H�]�ࢅW�n)톷�1oH������D}��5� ݖ11�%{�����H�iD�M�T*`saD�)_޿6��nP/�[5vf�-�Eq��ʝD�= Jۋi�F��ۀ������>�B[�1-���C&�<<�n�t���Z�cm9ص��myF�~H�T�ںs��E���G��g�%a�T/U}���h"zU��R�������Q�7��ͪ��K��?�7T��=��-wvW�5��ƾ���~n����� =t�{�)+��#�a~͙�D5�y���
�fZB��p��}$�ɰ�1Po|��3������ǒTH�>̀[��2%nL�*�?�3�M�U���#2���NԼ�f��X���4��6�<��=���ΐ�#��B�A��2[06���8͚�Z�I��{����¬�S��d��ݲ�ѝ�H��b/R�\������Ur<#Jt�ܬ6�kl$������_{<C�|]�f���ym�)����4��wk9�[O��X����H�.�T����`3����)�#���^'y�C�@DN�ZHpb& ?�-�Ig��~�Q�+vE�`�|� �j���&�����cr�9�J)��1/��3M&��E�®���ZL+�~��, ?h�*��E�ޘ�:d��PL"�F�E�ʃu��7�7�5�[�h�,���xOX�9&>�ʫ��RZ��A4ZeP�U��h�a |3�3�ڥS�ud��H�h.��"��>�Q�-�����++k�i)��!�Ķ=F����V�qVuθ��,��ozoQ7���'ok���aM�>�y�{�ON����\��ܫ����Z����D� b^�������q��怛���De����BZS�IW�C�v�ji��U���
�޿��nuu��.�,���G�>Y�+#�(j��i.J5��]��L�5��/�8>���MN�Z<��
�s&"��.J�O�j�E��.��N�trz�J�|�'y%�7/��e����o���B�O�8C�u#Z�(���D�t��/B���,g?A{�����c㋄'4�hP�7LvH�]��pI��E��IɋlI[���ɡ���:�(�XeJ�����WKԂ�Mhue�3�_���܊�ƞ����?]�n��4m>d­�������W�^G�N�R�P��>��Ƕ	����0%���+�Սj�܃`�\���ܙ�Zf�'|��]<���76Bh1#�k[�l����^�}]Oi,7�����c�j�&Qz���'��	�����Nz*����Rb�.�s�� �%5��2�Z���^���	�7�?�v�o��}�����9��4ʂagh�2�RƸ!���;D2�[z��3��L8�&&�ʎ�wlӅ��i6r�9�<���?���f�@�7
��c0A������[�x�`��0"4H���,�t/ゥ�Gd�c�]bᦚ����N�)�[�Ѱu���a�ѷ��<�Ö�K��R|�b�{;� �����9�9ʩI��5�!FWk�`��E�=䬶��cAT�l��y�`Ԁ����IZ
�l��������4;��c����5mB6� 9e�%FI��BV�+�������F��ݙ��v�Co�V��y+<N�)�j�n�଩�(W��Ga�7���O��wI	p�v���l!qW�����ۀ�PVԂh���9m�������o��T��C�����z��#��It���ay(�2	�y �Xg�4�@{Y��O�-�hK�v��bc��`x�^L���F��ަ��~J)�ϕǤ?lI���5S!���t�3U�<ҿm%�Ƕ�,�_��&n���U[ZO�.`��f/E��i�h+�s���\�N�1��
�]�,�(��
TI䫳ڧ�2= e9<�8r�b��ޓ�Ӛ�1E�����8ꤣ8r�ǡ�1���o������e����W�k&�%2�Z��Xv�5܌�t�(��V4ؓ���!�ņ�mW�0�4,�yXKI��k��2���|������FAKlŪ�ٿ���)K���n���M9���?��
����mI�}|����Ml����lv�H��v��"7')�G�kJ�,��o��d�+[��/��Iz7F%)Ͻz���q�����!
�.��C�4����=��M'�0*�����%Xu�d#�F�_O��Y�|Ȥ�"��}e�8���z� ��� ���:� ~�^�;�� ��ӬO��G�&��-򍗱�h�j��6��pR��K�#�F���yX��NǼT6y���PV�Ҙ��.��*���q�Y'�y�nO&3L�-���C��K!�%3/е�M���z7q��񻸰Ռ��ZAG�^B;��Q2�9��ѓP�V~�cE���7�'N{k4u�on� >GSGi �9�?��3h�(��yp��a����-B��)g���i\f@RB/�> �6h�m����]�"zT�������ǹ(�䯲Ji�6���E;.Tkr�n$h�������|��3�[y|o��o,�%@����ڀ٘�4�`I��+�/�|�q�TOf魤��#*���7 �0��s��7���:��љE;���Xg����IMFLl�Mr.h�zݟ����Az(1Ys/�̝�I���pq!]KNh���䧕Y;R^hz��,��cA�p���(�@�6Y�@cr��iF�*�����|��TC���X�^��a:B��e?��^��@��p��h�T�bb��,��u�ӚL�RU��:�C��Ɏ��F�? �8Z�Y��Hb��H<� 0��k`��b.' e9R�_�z�~�x��|!�)�A��$����\v�X¨㘈�	���̓S����g�C�������r�fZ�ǯ3	n��GoO8���\�,�܈�q֖��`�Ύ�
nDWF8Qj��nU&+��jm-{�k�~z�U�ДN%���P���`�m�/1�����ƕ�++N�ȋ8�O��3�X��5j��)S_��Ѷ��ORA����8U� �����7ԵZI�K�`��,�޺̸`��J�o���Z������ä�x`�i�i���dD>�m����̌�*�r�>�M����~��֟�"�@��
ĥ֒MI~�;��ߖ{[��2�Zwre��ywu�י�
q��!-�c����x�t�����F+��,ˏ�F{��^�XRy[~W:�)��Ű&u�ј�fN�@��r󧤯b0FRu���K��"M@�`�(� �T_��Xs������u�����Px$R)��ڋ����`���;����sx��dm��(C�$F��V�����p|�
�
[��9�:���\.h��I��O���Z�ڭ������PLS�E�T��y1>�Ey]��"�9�
.e+��y���Ɏ,�j�,�2(\"Fr��5�z؏�����/�a?���B�:Lt��o�u 8�`�)�S����vm*�-�uJ?�},�������j`��j���.%�M/i����`��~�x��������}G���i���P�k��"���vnZ) �@�qB�~N�nm�ל����)[ �f���`ۦ,� �������Bh�١��GH떃v��7`R��)�yw��,K.�������lUwH�[|x�WI0�vz9��dB%ckHI�	���<��b���A���}��b�_��=CVV�Fu��cnh2Q���+o'pF�qD"��c����<?1���4�&&{7�]�f�C�HOm�#Q²�AbQ�wR.S=Y�:���g��%:��	��tp±���?dl�T��#܍���/���;��p �b� �z�Z��Xao�;�gC�ؘ;֣*rKb��g �E���2��v��a�G*����ZE ��^�p����;���2I���,Μ�[N6�$����������!���3����E&��l��ҽ˞h�e9�6�ĎT�����cd�[�o�=V����t'���� jڑ���Sgt�2Yボ�Ԡٍ��u#ˇ��K�'��J�vI_��u��*C|ԩd��JGe�����(�T�a�"a��K��+� �͞�LtS��VQ�X�6�ġ�۬�����h���8ފ1�|j�f��:�zNd��pm�[#`$c���4d|J,|�o���G���fVnӭ�ν���ӗ��O'��	Yʴ�eڢ� 1��"22=���dk�Nd�"F&H@�܄��B� ^��T8-섞,����PB3�FB�����=���y��V�okP	��1wF����ϵ�u!�bp+Q�ͧ��-��GV\�?�_?�Fx;@"�#@���ꙷ*��� n�C�g�0D��#�G� ��w�,�E��r�t�_�p�-~C���W6�v����%��+������<����I�'�j����<3��Vv*ZQ-��o��d��٥=PU���U���O����z�9L���dS(�w��w��XQ��Z�&�z2����!�)��3����ڍgؕ�0�SpE��obR&�c|�#q��z�뚮�� �+����t�dL�FW�%/�l�k�#�L�.��,�6ٖ�3(k��9�xqv94!v:��g]�N���hM�x�D�M^�7�f0�U�DZ�_	FոS��>Z����K`���/�*��*�=���T�!n��R�,�L�(g��b�"Q?�jx��E@{�D��y%;Y��uͅ���	�b���KM�ؖ�6�ƛ����v��a;\�=:Vظq�b�EO�P}V���zc�33n��wHkULl\L��"-�C�'�d��& �@��u.���޺����]�+I���Нt��k���0X$H9�'�|��ǟnȔ)[��,�I���m�כ�v��E�j�1�i�d�7ս�=��
!��q0�0�[�@X{���a�|!�>��m���.%qf�XR��_̨�MZ�}z� �pt���4��Ĵ��_����C-X�aK��92U��@��Jq�N�����P�R�v�IpsQfE�5�ra	����b��r���������pu��ٻ���wJ�� ��������֭ܨ�o]��=g�e��,�8�3�Q+� ]�^)֩1�VI�8��%���������P�?>�tuc��H�C. �<��x{�io2���͇c�X�����^�h�������r���g�v>1Z�&5{*Q�%������;l$~F���Q��-����9�#e�?��>���H�9�<�40\�MHX���}����Ʀo�z�ƀ�n�.:�����%Y�0�zG{fC��o������$��mp*�ϖa�ZMC�1�GfS��+S-�N�#�2�3.�M�q�$uF��S��ch���� ��l��S��Ы)�U��R2�Qc�o�Ѣy����bI�H�-}��^����o�:�`s?���o�P��k��s�Ѧ�>ytו���-	���ձ$���U�W[��~���Q߹�? �f�ܩA���?�H- k��=�0[I����9�m:^������(K�6zSz�CfDb&a�iV ���脶��Q�_WD���Fo@��"�*tٻ�����)�_a�����Ț�jl�ʬy~�o�h�G�D}��k��B�T&�r2EEn��L��Qi[�$ꀮ4���V����T��1����v�n �M;}诹��$� �&`N4����J7]ꯘ�.D$�!��|�d��]�/��)�'Wzt8�Y���9� f�݆�W�\�%�X��a�d���LC�5��G�ҳ�B��L֫_�qQ����.��b�m#i���t�˘[�"5>P0u�:��t�d�=�	�B�e`����cn4&�]z�ק�H�&K��AǇ������Ch�{�z�@�%�6r���`z�S6[aU���|~�h��ր�x�0)��
w��o/j��c���|\�m�E�A"����:fGc-K���M����Y!9��<�Pd��9���K�ߥ&�`H���
l_��F�Q��%5�#[Y�S�^��cI����_�� �'E���� .��3%��	�{�߬�Z�W3���c����G����G��q��zC�9��(V81�o�[B�Fc�"��3 H><ͨl�z�u9x�,���#�P��d��<�)�ӡ�Kd�][ϔ+��H��$�,<��嫉�6l�4�윟�V1N?o�.��|:�H́V�E�(��
^��ìt`�ج�� ��}g��}�:�2 
ϣ'��)��oJ�ر�k;_=�
�`z؛��� ��u떈��Y',۞��.��J�|Q(_�g��]�ȵ��ڄ�� �E>�0:`�f<��|�8I(l�_�f  ��$���9/M�T,⨞�°��^��WQ���nd�@���������{�Ş���@��ޣ~�btO���wۍ�z�Z��!
(�j癯
s�ٷY��=Mg�=h����ѽ96&W�$�.�ߘΘ���WE�ة%8��R0�!L���G��(Ĕgk�w����L\s{ʁmj��;�ط����lP�P�!�.�Z�yLx�h��[y�aW�Ob+z-Y�&0�66q�0D� ��翅��.2�?wŀ�O���1����
�Dy�'��r��
S<P���ew����%�ǿ}�Q�EX �>��|�w�J�R
	ç�t/�Dհ!�|��x#��~�t��%�ܓ::���3f�� U�����	Yo����kNO!w1�"K�Sԥx��l}?&Z�V�W�P�N��@K<�h���g?�\����I�S�\c~Hfe����i��Y�Sp��J���9�6�ćI!�67���ٸ�Ok���9�������iʆ:�J�S��%h*����2X��<7�		K�1
pZZ��1-4�Q�	�^��_� �/�/ua(��>șd��\]�h����a/2��������`�K��7r����4g�	�`^IbJ"<�m�bL �y�!y��~�"l��n9��B�
1��'j��?|�-��Z�ֳ����`��{�����M��m��H�w��M���4��!;�������� ��E@Īg~j�D��;����<���r[�ހY�0  e}��AzY���(����)�q��s���D@�D�fj��рV9߻'^����;�]�A(�_]��P������7
�#�z`ͯ����~Y,�G�L�"J=4w���x^LD����.3���D��x�I8鷍hш�	�B6���զ�45cS29��d��H�Xܚ�G�
C�q[,����\�z��Zb�v�}v=��J���P�8�Ft�V�܉u)�� �4���ж}ڌe.���$�.Q���\�˽�Ŀ�y��;�w	C�f�½�n�1�����nᐡ}��I���
u\�i,e|\��wǝ$����[�����|�f��*����:�&�ns����X�3�������MW_��p�m�R�mtJz	jc����lw��s��-��&�UG*<����!6n�-�Y��ؤ�`X0��.>���8��FVDםA�eeKF���ܚFJ�X�� }���'`6Q��� Yb*ʷ��;/_K��c�����ހ��q
]���=�*(�N_���3p���E[��-��eq�P�q|�S;�hn!�A�_�'�j���-=��OEd�EYq��J���;��)���%�&�e����x� OlB)�*l��>�e3�w�a�=��:��r�>�_΁���zG ��[�n��g98�1�]Sr�Wyj�	3��va�
�*Q�k���[ºSL�a�����9J�|WJ�5yt_.����-R�XT]��K���]�����<z��Cc��A��-�}؆�#�4�ư�֤��8�y�Ѧ��h�z?�VMTSF�tM\�lsA5�զsvL���K��s�:��G��޾�������2���/��;�"��7BN}vx�F������R���`
�,���x2�����
F�x3��w���.�e�d/cX��K0�=�Z(T�����]ia:P|N���6�����_lX�ھ�}�˔C���F�0����� 
�W���6,U�Oɶ�Q�V��X2����:�`�{�Hdp�U�V�,��Q�֊��K�'�5E��YUי��͠��no��!�pq(|=�-?��c���W�l�E��+�w*��r4�,��HDZ����lw�9�~�m��i\pm~�L��Q�8�&��2^Y����e��lKG�0����E5��HS��U�/WjqX=�bh@a('N��O�q�{vL�K"����c�h�*��˿}�p�Y�����5��2L.���N�����D��?�Y$���n���t�C�oŔ3S����-X^�&���#�Ad���ޜ��n�\�x����^��T3h}����6K4ؼ	S��(�)�aҮ0���b�u��%��_ߤ!��� ,bBVm�u��(P�1��A�{@ð|,�t���,�/!'��Ȝ>����o�q�P��O�����Q ����Fo�#g˛�.����姢�+��,��<.Y���\��k('�_gm�������;M&J:7H�_��LYѣd�]6��w �j5<�E-�:� z�;��L_�>��x�p����LD�"YO���Ro�@7_b*�n��(شT�V M�b#,�6����ɤ�rNE�.��5��_�xBrȹf�(gw��\H�i��jo�e|���N�1F��rª�ͨa�9 N��~
d�И�IZ����
-��Q���L�`ˮ��|�y�u����y�Z�$ݶj�@�ܷ�^WSML�6R-s7�W��p��rȃ��E��#�;c~����m���X_G>��#܀
��S��%�l���h���U�&�G�ܠ��QjQ,o!H�%dR�{oP�)j)�����|��Ȩ�d)��FO;k#�C������GV���^]g)(��`s|k�-�w,Mc������X9�Z(U�h���s�,ت�4���lw���P��{��`zk��d�7��0m�CA =�H13��'@q(т:۪�R��&���r�E�gR�u�'ѣd ��8���3<�,�ԋ-x�t�D���G�1'����syݡ!�Vn6���ґ���X�؇��JQ��;���<�	��T�n"�M:�Br 
l9�њ4n�ú��b=$_6Ch����c�t���k:z|�ER,�w�4��߹��p��zC9n6�p�K�s���#(�zM��Qt�̖o��˷�4��O�'�T�W�o���4�]����@Z�ݷ��^
rB�͇��sZ;�>��6�ٱ>`4HF5@ۀ@����(�?0Q�u{�Mh��4��T�y��i�$s5i59tp��6%!EHh�I�'�|-�W�E�˨�6���^Q��=�*(@��0q�Rv���o;
�G�	����3T�cċ��ciކ��� %�T�c��09���
�%9�I��u�V=�y�/S������_��%Z�M����_�-\�pm�ؼ+��d�ƍ�r�"q�l�Y��SY���P2��^�`T	�Jt�E�J�V�J{eW�>f��Q�1�D7�rw �t�4�����^���\�ID0u��ʹo��S�،sXWz]�T�aUf��
�"P6�u����!v��}~�6�L�BޜO�L��N�ޯf����#�!�x�L�n��qx@�"�tzq��PD��EVj�0ǿ��M���`���ČL��G���>�5N�(ť=�0���)��y���^>�Eϰݱ�DV_[<�}g�N����9x�E{�yL�J��#�r�ATjFJ@���]�C� ����Z����=�"�M��r�ٌ�H����mM�A��!���7���8s<s��uϠ�n�zOT,�W��,��>Az����g�	�P�͐�Gtsn:9~��?�st�[����;�F,M��,=�(^��w�n���9�ج.G^����0߶�g��<�0���Y�窒\�D��\���۷��|�}M��0c\�'����w!k'Z[D��z�늻 ib`�@�AB�ݪq|dSA9{�;>g�G��fi�_�e�-X����O�*�-�`E׆�Gk7�`L*���$0��\��v��.G����(;��K4Qfr�XK����@��:�$��J�kt�����⛓�d},Թ��-�u"�!�ឞ�Far�t��coϔ�Z7.��	Λ\=j��%V������ {�t�8-ܶ}8�s��<��'%�߾�C� 9�z����� AJ�S٬���u���P�PH�Kx�s�Yx�@����򾬝ߖ�S�8*#V�QC�ni��3k��s<E��a;U��p��+cc�1�$��U�j�&Qca��.ЏY��rX���� ��U���W7?m�%�~�tnw�������
�}q6p-c����d�>$Ÿl�U�����7��D� ��q;������<O_����Z�)w"Sj
�����1�u�uVAcZ-Q���%��k�Ԯ/`Ӭ�b���ji���P�֭���h,�;��<y?�� �a�勣������W/w1�e��'O�]�j��u_��v�S�¤�:���
U��x+��s|N�ǳo�]��`t�W5�n�۔ƻ573"p掜��NS�\[f�nwb�S��o3���ǜ��x,t�%I���˞G��&+xI|5�ս��H��E �O\D?lѓ���q}r{NX�FF��e��E�~��ʎ+����w8a��VC� Wg7�#6)T���y��C݌�0�7�9��!�'�����<ɼ�r�9��N��Q'6�l�]��dF����Gg���\�d�0T�"����"Ph�K�?�h�=�������ֈͺĜd ��y��_6�5��uc�ʻbL�v8�*k���)�g�RK1a��c��X���1�F˄lNbl~'���Y��#��C����S��KN�������POJe��9:�H˄�\��)��2.�����M�Dt#�O�!�  0��+�\�fJ�#/�^=���8���(i'}l�%xl�M���a6�������������&�\�˸���[̮��PQLA&��n/ej��r���>�H������j�l���/�� /�ٕ�^���H(�Pd>�W��q*DLf�0�-$Xh	�7����{p	�1k�7�G�*H�c�V�~%ܗd��%��v 9�����O&����WR<6��-�d��;ta޲ƪ��j��14���.쫫�n��aꗋ��%��=0�}�w�&ɀ��O��j?��d�%�O3u����W���<�$�����S��0�I:�To�RS���cg�i.-�p��o*�B��_�qdX��j�)I\�&M� �H�������[/�<����t�� `IPi�����i�#ʠ��Y�ʮ����}:��Ժ�䨲�5~�|=����>L
���@�CMk$6~�w��������k�3��l�B�u��Qdi�qK4@�qtp�l �4ݮ�>/g\K���*�KL@���3N>:���e��65���5*�.�����D˽�~�ζҔ��%3��J�*�.n���I��a��Y!�}�Б�1�O��9Q*)��F�i�Ȧ��Q盧;�l�S:�����Cs���q �M�8��F���2x�*��W�d@��xL!��<oL�$c3ܠ�͉Y �v$q��ae��o�T�ǒ<s�,$�/C���o�q�7��6�g܂�Ϲ5�^WQ�!=�7Ղ[�tַ����"�r�<�G��2�Ж��O8K~HZjh���S4\\�,�Ŝ�� �&k���*N��b>��I��K��������e��1�p�mu?7�"S������7r���%^9wu�%e���#V�eR�0��[zQZ�}T������W�h�o��(�M��2\ �=��b	~ _��Z{����7�
�0�N�2�$U���kX�cY�������W�f�>J��`nS�@��4���rl��\���oUI�Җ.�Ql������<���U ��/2N\��g��}�K.[
�9ݱ�<�b;��V@s�N]�q}"(�D!���7�W�˪���m>PP`�(�az$�>Y$iy`d�HyX�&�?���7.�"ܖ�!�8�������H��n�tEMpr��[��	d��D7���h"];���[,ɺBK\L�����)v�Vt�_ �7T���^ˎ矞$���9KDox�Ni$�#�S
��%Q�e��v��d�%���c4�"�Ɇ�,6�*�8G�����y�tWݞm�S�:0I]Y��"#l��S0��q}��@k�;d�8��K|�A�� SW�Z��E��!����I�3j�u�3�8�5W2:i�-���(d~a�iv�Ԗ�I�sb����e�W�H]B[u
��d�jD~��B+�w��"At�;(٫�e��L�,G܉<�8�P�N�A�$�w]�G�4�$k�}Y�mXi�_u�g�m��>̇ն�,? ���(s���~�7��e]cOPm���� F�zc����}m��
c��*���~��*�?ɕo7�>�/�z��̳�0W�W5N���"�����%�b���w��̽m�0���=D#!Ъ�
�7�?=^-���]�Vn��f$��F�|�u����T�iK�M&�n��@��_IG�j�UP\���[Hx+�7�gb�cG$@����n����zk~���uR͵�ݴ�A�\,(b��K��ԣ�8�Q5�e��D)%wj��<�G��ks0��+��(�M£������,fkV�p����J�_8\�t}4��w���o���0�q�l"��h��n�N����`y��\��"��s{?��x�cn���;f���"n�G�[���Y��g���ذ]�,�2� s�_�zW���M��ͥ΢��?ȸ�n�⯉	���ô��$����A�c��:�i�����z��<$�í���J�~��4�	AmEB� �~�~#�k��5����Zc)GKu�׵�A�p��Fo�T���ҪI�`�yW%٠d�~o��ZΌj��փ�r�Iv�R>�aP�+�Xcvv���\�X\{v���M�U��T ��v��.]��l&fIe�X��N��H��[-���&�jn���iF�� ����K�Qȁ�?�][q�H�X2�N�̂�O����������1�k�c4B�äb-.�E�vc�OIQA�鷾'��H��޲ ��S����u�v;�=����):�	j�v� _h�g䑦1yp�]�W���ƥ�6�Y��< 2�.��c�l<� ~)��j�C��wi'+��.�ԯ��7z�`E-m�?��	o��ӭO�ܒʞ�	�����/�A����@���d3h&��o
yP���i�6+;���UM��@�!U��C��hJ������b>�6o���xNL��4���\F���Ty'�l��-0~���y�s���ӡ�/����KJJ2�{�N����jY�T�����D��6D����6C⨳n�v��F�vq<������[?F.\4l�$�(��E�TQ1��6}j��6�Yu2,���KQ�=`7�b�bk�ܮ�7���R��Zk-jҽ�'	��"���|��;�g%8�3s����#�J��1 �5���	Ƕ��`C&K�����]@�*��1A��kWc'�%%4�����YP����FE���>*\�ZG��!j()�p�m0�lW��$��3�!?��|(��߮���ve0�$�
����%�!P�{�����ky~�N��v~���#�Rk0��Ks0ګA��3a���P~|�1� %μҲO~�#g+�9#}�>�B����9(/�@�!<����"	]�5��Rk�y�U�>q����dz��K X�Z�,L�I)N�v�q���mТ:J+p��E�W�W!oR�>��A�e���:�G*_ �'�.��]T��lķ�%�1���&��>i��S����>��S6C$|�;�) d}�zO��4����H��ɹ��ƕ�����v>�u��t�m4�:�,����K��]������T�?�
�*rFW�b�:dn�,2�~�!K�z�1#�mW����̴:��6�_`hĉ��E'�1Na	3c)�Eз�=p�����x�](,��J�g��Ӓ��=|��	+�`��2�a�etrs�׮oQ���1��tؽYH�@d�˹��.�m��y�PD��c�k<��.~����dؠڵ�xWiGj����㹗6���Y��wR����l��(,���n-�ֆ���1���P���«k�z���W��pN��0�L�Ck�q����Qu�2����i;�
�AI0gF,1�$F�ȑ0�� zإ��ˆ�c0nɑ�o�GZ��~t�Wd�Y^�֙�UeK ��\G�C��`��+���u{7���΅_�9�6�k t�B>��#Y�Fɐ ��y��N$]�9y��Op$zg�7�0� #����������� ���#5j�o���D�m3\V���46���΀H�f7 i����#�:�pb���F}��vG�ĸ��1u̾�21�yQ�ɦ��lH9�O�UEN�N޷4��$)\۫�b��Дn[5�4��E"�V�b������誀}3�>ZB�^Ҫ�V՜~��M�5�MI*Km#�S��t|Լ&�? R��S|�`u���o!\<����b�
R��tO$Lț2�t�_�p�BS�͡� ���û���)iJl<�x���[z��T]0s���"�X����a�1��6���.�IC����z��l���	ŕaV�NQ00$�P�W�\lꪌ�[ݝ��'��"���b5�*�WewN�M���䉦�.� V�xD��zIW�`�@{�ڽé1cE
'�� �dJ]�Y}�q�jͥ��b�1�ya7��p�;p�gi��r���ޱ\�����Pe�O�>��|�����9]F����2ī T�%l=�ۍ��˽��Z����v�!����ȃ�bg1a6��A�6����K��C_d�;�#O0�(�n��w�X\y�C�s��^l�
|����5Dm�*�K�$� �S��x��/�8�6��m�;QeY���������*�f4�}�dn�$�Rs���q��u�1�!Lpڸ$˭���>L"��
�S����)���c�����q�Tf�7�?�D���?^& &����z�;x�~�Nԁ��r�!{����~��.a�����C w+^�Y
�-�����e�/]D�V��d���*�	�Gƴv��&D�V%�P��.L\~0=�L1�*�[����nk��9�[a�i�QC���B�/�}�1`�A7������pa휟��5Bc�>Ǻ+��3���tl��X�C���鲗��@�����	�qY��i_�Ŀ�O��b�6ɶT�j�򩊗��B|�0} lWS�F;���B2Gō�7���j�yK����M3� �`ZZ���Ҙ�b������U���P����d\E��f�r�?�v�Ԝ��'���}y�A��t���K�"+�X~�<���!Q>���j�%����z��P�^���wG2�Y�w����!n�gdv�	M�HN7�0jgJBMF3��������t�p/��f'�(k,�[����M'y6���g�.�n�������(�����W�����]]����A��R�J���[T�9�{�*��|�c-�>���H����N$��>��:y�2Y�"�n\��)}
�����C֖�B>�b�}C�B�r��B�ʾ��D�[�JWk�0:�hk{�.��又j�w� ��$X��C�G�/6��"�c>�6&��ERց�E�ы��6���ּ�K밫j���)�v<�&�Zq�)�)DW�t�|0kM�{7.�GC��`S��o���D�.����9���_EV%�G�����3��Y��J���1<n��t=�Rrj-6]^G˄�� ~��)����*\pp�Yv����O� 4Ւ��s�(l[u$]���Qɸ��~g�� �̿W=��n����U3�>"���2w͕�C�gr�/��$!�N�
)��g�-�,á�0���S ���}���K�L�>aW�p��՟��uO�,e&��e�XC�Y�v5R��qB ��@��_/Yوղ�dp@A��#ѝ�fc�%�ׯbH�7�Ԟ�,޻���H���,e��8�md3�tW���2KN��}Tt��)YYȦ�u��.����5�?-�`7���H���j�^��<�C��C�����u��L�h֡.ކ�Y�3	G9�`2�:��{�7A��8���}�l4ux�����aqT`\��u.�2���*'!*M�]Ɂ��T�f:�u�Q�S�,	�-���;LC�{=RH��cZ�y�(��E���%+���]�1	����T�`�y!����F@��:4��o�w<�k����bTtSZ�vf�{v_�{�[���AQ��0nt�V|�CkK�M�V������(S��̤E�ӜΣ�@��S�.�5��Q8)�sV�e\H�H�C���C�,�u�T}3 ��v{��5H�z&�����o�:i�P�W�� ��]:�^/0k<N�N/vᏐ8K:�a�~��h��^O��^�
�2����)ÀM�2���G�j�A"'�F�eutZ>i?��dr� ~����ԙ������ƪ�I/�|�Ùߕ�N�%JfCq�(Yxq��10͒���Ú���[ޔ��
����D�%�F�f�#c�*%*��m�iS�:3�wV��)�Dؒ�������� V�|Wo�]$�V"�|�t�o�L�0m�V;?���*���0��T�?�^���Ņg4*��y^�]��Ǻj��O����ՙH�溜pO��?���1�@G�r��G��\4�޾�U��,�ǂwL=�U-}��6y����1��K'-m,f���C��S�	