��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��TdO���ښ+�j8(�aS���x�YH�O��ʅR��hT�����K��n��o��T�k�E��7�����*��{#&����<9�� {K�C��4˄��Νf�߇ݡ���"�B(��,�W�?�8)na��{�� #��4�!��5�1f 8�>�m�`�LE�d�l��	\����Ӹ�&�:!Z"��w�P_��
�5xMW�~��~�"����n�M�f��B���	)��FÈ�=�����0BE��O9�N�4Ӗl�(�g9����L����\�֐��&�O���o
��#ƣӯߎYPAH)�����K����_��]" &e��
�v�8�H��W��PZ��lJ���WҚ�}��,��O��2����T%S@��A��=�4���0��CAQݴ���%�ʽY[�<�p�N��I2MV�t3�\S�p����"j֙�s� J�n�ft�̞x��청���K���ʱ1�~	y��?o֑t���9�©D��:���v����]i�'����&[�׌�MC6M����j��-b��л�!��g�!t-.�E��)wX?�Sm,*..gn����5��ǵf��e<g�M�^IЫ��h�0���W�3�ٳy��,����� �=WEi��V�|�zӞ����~)Z��������iݪG�y��S��e��f������6�M�I��l`�7�ܭI�=���%_U�L������E�E�U�'�!��\#
�Ԇ�#_�(��n�F��ӵu���]~x�^���R�t���M��
��Bx���>
G����|��5���-K�?��|�
�W� ��	�/�W��a$f!�X;��v�|��0?ݥ��d��.9�O��zX���#�����@��G�Y \+ c
�](��dΊLJ=�
v2
���rAR��y�DD:6xt�hs��wJ�y�©�'K���"e;�)/×��l�<�,�T�H�g~�do�~��ɩ"*ao��d�}5q[�BZ��Ρ*RYjL����Y�1L&�$O��t?KBԾk*���k;�K	���[C%�/���W�Ơ��d7'�ć������m;�
HH8��� ���,Pd!��n��B3�Kq;YM,)�cf�!,@^�H�	�y���d`�R���NE�("H-��Ew��XoE�W�7����B~�\LO�����5�×6L�c�@h��W�J�ۖ�>N�S>�,p��Zfx��XN�=�4P�
�ޤ�I����e�F�A<��^jPǨ���	���\[�L �L,Fr�JaDI*��gI�+��FUy0?: ��o�����Ӭ�͇u�}(P��^xC�]�aT�@��u)��[��/_�#x��np�6�`~��f5���x78�[�Lc���,*�ٗ�Ϊ|.ׯ�l#Z$\����#|��@[a幧��g�V�:�A|�3h�ږ�4���o�*L�R��R!��`�nڑ����_��,�N0���J�T9�
8�}H�'��"D����]ڳlG�I�a� 
����P3��w �L����� ɂq<�U�`�M)��񰀿{�9��\6�[z� O��p����$\���i@L�!6zᖷo�D�TRZ���B؀�2gq,!��z	��(KOX�yBKhl�79�D���>�ԧΩ�A$9_�ɿ�<�0:M���\�/$L�� %a$�W�G���SJ�n��DRַ���Z�Ć��g�B������~��0�~�Em�� ���6b/f�A����޿��i^��Z~E绀��	s�4���Q��Ib\��T�L;<u�+h�u������Q��76��,Q��B�V������ݿ�>���RE�WF�9�;� �d,0R�ۧ����h@T0�6�np��OK��^��;�{S�u"F���� �C
�iB��Ih׋�;ވ/_]s������
���$Q�����9�D�4��b���V�UQ�K9~���xU;d�*j���#1O���k�5ޓ�Ɲ��hO};��#(�3�T�S �}d���'8����CKCWޖ-�լ�����!��2d���nK��8�WT�p�O�w�0g-.u>�xz�]�:�F�lèd_鐔)�c�4�4�q��nd���̈���$\�6�vG8S�6�lU�6����P���������}��o���ț�>�\7�#j�=E�U>F��Rs����vG���S��j=Fެ��Z�ȟ�"�e��'?� �@-����Җe�R�}���v��uA�X՚�j���k($3{�#W+nzO�e~�1W!�)��U�!��< �H೺��R�H!�����ҷ�EU��Cv텯����<�S-�Tl��i�0h8�F�^A�#��Ⱥr	�KO�ghJ����(��3!2'/����şz+�طtӰN��[�'��̧�x�K�M���q�M�(@��X�}�qx�B�`n�'w{����z�K�8b�X�
�-$Ȅ����H+��eL'�}~3H�n]��n�Vk���l���K�ο�Tǫ���@��߰*�(Q5Fm;[�Rm�*X���_�S�e ����_�#����I\9���Q��������"e�������8l���s�Ǌ��|�a��$-����t\�����2���Ru��_�FZ�pUu~F	Va����{���Tt*��ں�5v�W ��b��η���ݛ�LB�4z�}^�" �H<����=UD�T�L#���Ni6���Pef�)#�ص��œ���y\�����Ik�U�#������l\Id�AC�H��x�w��{un��lAh�������������G���?_��K&��� ��"�����~:,�5�d 9�Qp��� �W�7a�D~ft�H�c/(�����^ ��e�Ř�5�cn�\���M"�jw�),�c˰��Z�|ՠ��Nj�tW��WN>�v��w1�DQM���4qhOȠ�����h���t���Q�CGjF�%^6,�sq
;zBG�]<�U�OY5��U�,��c
��yb1 ;r�XCy'�,w�_����Mۖl2Cc��-H�9p�T�]^�������D��ZD���V�$�*�)������l����>�Y��k�NaP��2�e��>Β/7���L�(��L-����&���3� }��ieИ?��J�Ԟ�jh'���L�[^��f��	6��eO���ߢ������3x��h�Rpڷ]~8��F�õѷ=?GFmޫ�J�����Q��c[���-ȸ��M���'�h\���o���	9a�H�Gn�^>3#�T^(uq@a��E�l���Y
�i���ڄ�#��w�-Kq�(�L<+Q��.$8�d�NZ��h	a\O%Y�&�d>>n�����iq�����T������#7Ju�(d�G!�&3��Z����2c
p�,}��qՎ�r3�䮬l��o�����b��NkKo�}�n���]4�[H۷����6���'�#=���"`��+!ڋ�� ,O�J��5!c����H�K��j���օ�1�Q`*A �C�U�8��
��P��G�����3ϓ/Xʶ�&ő���dЯQ��1*�Z��ʤ0|=��`fr=�?S�ར��wd#�~�]V���*��}c�c��&JWs�l}8��v$#�	4� sE�P�Ā�D�U2Pz��=����Z�>q��{�6���C��y�����<k���v�Ñ\����TS��-cY�@��5Ŵ��SK�1��*��=��vajE��+�Q��1a9��Z�o;J�8�%oKmz����ImO�ky:���%�G����⫼ֳ�r�R�U�7���'K���U�"�$�{<%��om�q�;hL�`�?��/ �-���]�'��%Q�Ĳo�Y�yG���0��v��1�H�uzN�s!�7�/�$۳��iG�:��})^��GhҶC��(='<S�U`5~��r�}��v���I�2H��P�+"��w�
P�=�%���ӬaXW����X�������>�+�֠ ����b�|�!��fװ?"�����ͩ����7�ss|���E�)=��:��+n9�\�oT]݊$u��3b��H�Й��,���Wv�f]�f��JI);�Q�5�x�]]U3�8"Ъ���X�_)��@��|����}�T��{w>a���We��J� Th�R���yR�WY ��]���3o���-j���P9	A��!QM��t��Ln��o���� �n�-޿�ƕP9�\kĬ����<%�_����P��b�\H_P|u��Sz��E �:�X�c�gET�9�m��t�C.�����&�]!m���2u�[���8��\�6>��6��8��n:U�l	zzJ�q�Y���"	~�{"�{|w5��c-�o��=��?������,k�'�O^��S}��31kJ�.�����p�ay���C.e��&�d��Ć��{�Pe��w�\	� fM-��'1�s�[�3��.AQ�L5H�x)lL�a�k�p��F+a@q;U�����8���f0g~+��uK�����
��z�mVVx��-IΓ}��Y�����ZTB�P��_��s���$v�=�Z������t�� ��