��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��N��~���#r�p�H�����W5G��� �ƙ{k��U�K��F�����ZE�?��o�d㽈�{�<����%��,8��d��P�7�t�.����u�FqU\\�'3x��Wx���
����h9 �0��Q3�.?!�*M���w�*�(����<U��E�4L�b�3��Pkӏ'�b�����K�^�N/�d�ЪwR!��-��^��J�yiz~��f=ʭG����=^��������~�)�ꁃ����C(�{��Y����	fq��`a�$�]]��Y���:[���h��4Cw�(��+��.bc�a�pz"��]��Ғ��]ț��*�-�A�Ɖ��ҋ��/g�������2�"�^%%��7�c����5v1V�ۓ1uyֽ�D$��}��+��*L�7U��xh[b|���������0��ۯ�濙��\Y�o�7<)�mUBsn�dג㛎�����K��3����׺2W�9:�}�[�{+Eh<OU�7(�?j�T>��y�C�'�fi8�+.f��EA�7.^�;O���h��L~]R=���5}(�?a�	^�aj���Y)��M3�R�2�¯ �u��Z�I�d��F�Oǳ/���eZ.����`p��[k�^�w4�ȃ���L?�X�vK��R!ג��+�\_�`�\�/�E@�g>�d���+��6�w��;�@8���+i�i~Rh�B�u0�;�0�BEc���0�^�uq�Z���˷r�~c�M�_���Y��P%��FA`,%�/�2<�������n1<��iqN; M#�&�#W�8z�,@#�ϟD�]��Š�L�:���8%Ula؅iр`��y�����\h�i?�tu�C��Ο5�z��췡2�r�����[�P/�5 Q�ۃ(eN�i?h����4Θ&>�F-"�:������߸�18Gg��Rf�c({5+��JR�6p"�l������OJ�%���f�3��F�����b�Rq��V�9��1�6�dì�q=I�0O�#�g����yp�[�^ø2��0���$
��
-�yVI.���H��"5Z<��%���g�C5�7�	Ƣ��y�ƻ�|�Wܢ�E ��
��&�'"ґ��׻8�0�` p翠�h-� x�ڟ�I���b��ҍ|�NY-^�s|]��sZ֤�g����\���d�dJ<5I�ؼ�S��?�<��_~i �fh�ʚ^��t@�и�;����J$u�ԳCK=�����oD�K��Td2�63ܱF>�c^D���I���LAV�V+Zj=uN:O,>=��C��z��	����g�ἶ�Dv*<F�Ԍ�9�}�e [�O.��!�m���.γn�{y*	���y�,G�G'�ټ��,T`����1r�@�0S��7��Ԕ���aΘZ��Iǟr�K�;F��vL�����5x���E�o��47λ��:�����)��g�뜷p��e���al���tCB���|�#���%l]?�3�)a��1���:P� �|�gGY�v��O�C4�`zL��=W���q˿�Q�Q<������2i�=S$�2�p\�ҷ�:�c�nTcCǩvjs��ZԗC��C%4������u��:6�[y�p�K�/�l��z}���,(Q&�H*�~���`��Z��{!��F��H��w`Wa�2�s�q��f��}\iv�U3^p���͆����#�'��>�H�ڕ�E�Ħ�l�CT���4x��S�>j�(������`ъ-a	�$�Vn�!��9��y�:-���i��F���l���p�yܑXH�y���*4Y��l��gF'2�F����a�����-���"2���D�Y�\���4�iIہ_�EY��.Sz�se�qw��
S�
�<���u�8V��M�&��G�=%C����6���� 4���?���[�Z�mGz\�ˉ ���0��T'k��ͧ�i	�uC�2�
���j-=�x-�H��vg��vq�"�;�X$�j	����s_�e��H�ѹ{��~+R��+!w����P�ٲ��Č��?	oWW*��H�0ꏘ����}9�f7�e`��NբM��Ƃ�0�R��#�.�.�@��PJ����7��E�f0��N�^=Z��h\_��ԍ�UY���N��ü� ;`=�]��W�nh��@�3�<yQ��>�o�Ǔ9V[LZZI�`��N�'��/J=�N�!��G�h�e@U�����ₔGV����M���A�Q?���mX=A�~[�pF� ?�n�����J�hIYt�9"_`)S]�/�싞J����K�����0#�/�ZY�
��x���[=��a����+�@��B��Q�1�v,2�����V��ž��+߁����ϩ��_�iXᡣtI���1�Of��s�.�Ę���P�2�P��^��=rU�d�&r��U�k� ���;�v٢��]	^�^} ��I�*�TAʙV�u����/�"f���V�7�>��� ��s3]�S�jw8�wpx7�"%9,m� s���d0F��h*Oz	U�����T1"��������!���UPsǽ�R��xF`6�~�[7�����J�J��]��<���B��G�^H�@�"�� ,�Є�w׮�:�
%i���%����������Nj�[��Q�n ;�-��.͛7��7oOJ��%�3�;�R��{'5l��H�'�U#8rh��|
�|����u��@N'+o��C�����`� ��j@`y���Y�� ���pdZuW�L��Z��l�s	��$Q����܊	_����=W��m@�6q�X�ZhP7B������&Z�Ɋ'>�u�J�s���.$����Z5Sk���}�'8h�s�e�X�.�%i��q$��(�F�!����D�g�ol�RG҆y�72�}�Sf�Ko4,�֝ւ;�v��Y`B��
�ƌ����A��hU:�	*�M数2‽���t�b�}���5��/
��n�#Ge�Xm���3;S-R�&�ER�PJa�|�&�DhrK�aF�sbZ�&�Q4z$kv�F�C�"]�L��$�����H�K�S��|׀YH]��N��=Z	���AQ�\B��!����pA\��݋��,�u}��~.�P�D�&19�J�Ϝ���Y�$vm�E�v֊W3g-'����N>�	���~��!/���"��0�B�T�?���;)W���La��f�!�<���i�s�st�l$Ų�v5�K�K[��v�+C~���bs�0�7�� �cS޻(2��O���� 叝Xޒ���t�����Xt������OGgs%0�.$~� �V�w�*�M=�0U���M� z{*�C�J�')~�{���ku��k�t^�6��z��% ��A
���p�g��c�4t|��Ũ-����n����%��8��Q��b��J\oՊQ���KH2�P��VNO4��9�eh+Lfy�1�8���0yw���X��"�Bȳ�?JY�b�X��Vﹲe� �����2񐗡v �w9�?Ȓ����>�p��j�{ˏ��,]�lE��E�@�{�X�T?ʈ�x�Mqڥ�e�ά��R)��a��#Br.n)���\}�� �l�P���|E�{u�T���t@�8��+�岦�Z�$3�����������F��7Q�7
�-n��DQ�
X�v�=#%K�_�.y����^�Ѽw�^n��h%���m����)9��mힵE�o�ɬA��!Ms;�EJw��K�Tp��],���DdR��TkmV��j^�A+�_Hڡ<�:-�&h�N�b��KDч��"���@M%�hӦ%�6j����|u�$>"p�ˮcH�%��Ua(� ���0��Ux0$��kɲ@���T)�?������נ�i�S�IL�K�o��u�TрP�I��l�6#�˴؏,�op�~�#�:ν�ϊ��.���}w���>5�ը�z\sB��6ᨨ�ᬹÓ�oC	 $s)����rOR�UMw��:IN�����e4-e��/])UΚ���Gf�6�ÊCPz�|�}���N�j�R��+Wt]ˣ�������0��[&�	VOMK(u~�"~�@C*gD����9QZٲ)W0!7�}]�^9䒌*&��w�j�ё���DW�>�=�_���d�=/���<�ql�
���p��vU�Y�����}�JUt��U��^�v����N�V��A�I�l�������U'�ᩚrX����/6r�S�,�����Rvl�9����p��Z3u/J���G��� ��.��sVlh�&�a@�
���6�+[�H�{�^�z�s�v/�Ʉ����8���X\%�|qp��4b\ �\&M��#s6�Bb�o����sX��`9L-T�P=|�ꓔ6xzo�nyf\[��
tH��4�^�ۺI�_��:�򑇮��mǯ���Pۦ�c��M\�ڴ�y�i��U������q�h��H�׃�f7�f���#�w��_�X1BY�˦���Ҕ�f���}Ä��ov�1�c�_�a�<�d��^��
�~Å����u��h6j�g���ƛ|}���q&q_���H]�Lj�3rO>pM�q�ݼ{�YQ��#�bƞR�v�O�i��q�?�E��.
m@p���K
��,HV��GG�VJ��6�ߒ�j��]B�����{��lA?�ퟆ�KKRQ���@�ݭ�e�NWʴ9�L�4��;iI��O�H�:.��.�w����<7׽M�ON�������Ww���q2H��^@�G��y��ޒ9�y�un��kڍS�Wۓj�|&��jY�\����SM��|Y��ّ;���VY饌�]���t�ߝ����'jH��,��T�k��7:�#�%�a�?u:��S�MZM7�ͳ��|�n��۟�������M�\��#�TD*7,���z�2�R�����|x�?C>�qW���l��R��,�%ބ�Α��{�]2��W2�w]�x���-q$�:�ku��˔	���b�`�>��î����)�Ц��l�e��]��W!�"w�pw�!̕M���Sk5}��$M��!,U��T�X�5�zw9��aZs�8�����E���e(��n��o5�'�������ۮz[�H�YV'U%��7E��0�������AB�TҾ*�9�#m����c�bpuB1m��!&�P2�2`r��_~�{�δ�.�Txm!!�a0�c��hE�b��r}�^3�$3�Q��6�p�.PWP�LWU�5��Q(['Cq��Y�D�GQ�6���@�^�|J��\�i��n��8m�O<O�&8l�����I0OXj�!��g�v��FdOM�M��<���ƿXG���ӯ?��	�@��!��Ze�i�p�oAgq憕HL3Ȟ��-u"�,�S=��������=���@�P���}���:�Ư��ZHX�4A�pԓ�h�,r�=��K������-M��?���	�BL�tG�v�xx#R�b-=�j�[O�BG��v"����c��t-��`Ԛ%	�:�6?G�̵7e���쬌��"	T�j��g�R�G����8�>�E��P�6D�I�¾���(��S�朮�T��-�g�6nT�,~��W�8%փE+��rKC�Ӷ�>LI���Ηi7��+�|l�u�$����if/�]0X0�"��O�)�٦ϩ'Q �eIhC׌�.
� c��~y�sC9�*�9�l������rR�i�%w�u:���l� ������KDe��1��3G�r��h(}B%�����KwV�c��	џ�o�t�av�蓳� �6z���c�Ɨy��g��-�+�mxt� n��HI��8�]B6�M�}�'�70���T~���(tip��uMetE$���yX�j�4��!������HcB=x�kԠǅS�%�k5�}�zj�9�����]6n�x�@J�ɝ��Af�~�~�?(�ա�5A��w�J�8D�*v�J\�!��1m�C��{��59��c��~7�Yα;��B���Œdw�j���#pŲ×f+�/�vtd�-q IX��]�vCZ��b!dG����j:?q&m�v?q޻
v��.���ߎ�c��=/9�%�L�ɤ^'.��ȟ��tk���F
�M��8�"Qu� ʿB��7��z<P�ώe$�s�*�+6��M����	}�ɧ5zk&E���2�s=�;������̍��Buǖ �=�K��|��(�R��	s�?˒U�9o�+�^7�1rt��K���t�~J�¿F:���c�c��	
��1��v��$ۙΘ�.0&�uؖɻ*������C֖�T�NO�c��%�(\�@�OT�!���W)���vs���e�>�!��I�lhDEбy�s,�`P��I�eRTƉ��d:�a֎�uo<R�38�W�m�f��r�A.ɶf�%V��4I�RW
�VD2�kR�7`��s�rݯ3����M�c�ڽTMi!�l�g��1h>��	��C���QX�9[l1��:�KJ{W�M!qlIy��(�K_�ٿ,�As�}0W����_��^�V���җ��=��6��wA!_��姫ޞ�BDdu�t�i�q&?�r���%��h�I�U�ML��@X'��⤷ſO�~j$40q���[\��Q�1W��,�ˤ��\�-�gx��s(���\ZT�ԉ�l�of�j-����J��,n4���3�����E�ٔ#5�N3W
1�t��_��)8a������n�I��.|��[����uw ���F�	����͙|7k�ϊ8���)����8;�x��{	4>_���_�,VP�y�b�i,�����kyF��d��Jh����X~0H�䧓��T�v���t.�}A�pkF�T"�8\`��$�L�uy�+A�����6��4�^���|l�]�ICk@�j������֮R�뻙g'!q�������9ǒwNG��Q�LIp��#�� ^Z��#dm��}��Dق�8��D� `��&��#�fa������#]s��3��RO���,!�$"�}��Yo�g��
%V�d!���Cn���⇧��kU��s�t��D��JtS��cfL��ܗQ�X�>��'�6֖�re��>�/%�H��;�l�����N�OjH瘖�6���舸�>�cE4rR�3yB���-	[g��������]�~��Iބ�۶��#^�����a���!y-�7��@���%���7!J��4)����!7�q��nz�Lt�x��"P�WG8wT)�ǚ7�L{-����Me:W5�>�S=R��.t�5~$d��HK7�b�7n��$W{�(<�v�lljl�h'(�@�����c�`r�_LK��U}I���`��պKW8Ѽ	�Fn(7*D�ʕ,����u�蘆qY���~[X������M��r���!*=βea���h��C5�H����_�ϲ�C�&������~E�n�΍{$Jȫ���r�䐫�?5T1�$���l�� ;�ggy
���63��X+�ڒ~mRU_����w���FpD�6)���-9'c��i��35����;��,zd�����O��%PT���a��-�j%��1 x�< �WVS�k8)�I�'@�{���iR<�E؅#��,p���|�ۦ��Iu�5d�嚊�������]ڽI$��ݐu$�H[��g�s�-IcaP���~60�+5���T��� i���$��>^`ҟ��L���?��-�7�pR?P3����wε<�e��,�0
��i���s�Fs]�n��$��=��e=t�8R����
@kn���tЦd���:ͣ�޽��Y�j
P� �r���'��UW ]=w����X��~�p�FfzE�}�I��y��
�/��h7�J��PT
���u]q�-{���j��yJ��W�y&��$���Y��)3$�?���յݯ��I��隙Yg����7�/�P�V��}��$����	���/^$n������Zc�"g�r�??�����:��o�lς��R�
�����)VPЏ��3oG�#ҙ~�
��A�I�Ñ��Ɯ� �gO�{1���ģj	��y���)d¤��f�݊�r�-�.��g�M�������/�ū��J�z2����ctVɧ�s���fh������NW�A;?�"�|-��~�j�0:��6�Fͨ !<�⎮ҫ����K࢑��YX�3)lE�%���6R�ڜ�?���~ηؔ�B�.@����i��N{S�/�2���?�%���NC^�`�<q�~�݆���c!Aoo��d�gI|�I��)���|��C�=��rf��Ɨ��� ����=��Q��7�L�?7���1�Kf��.s�F��.���!j%��f�n��+�Dl�>�b�l@�7�i�N�SH��)�a!ǥ����7h�X)����-�I�Y���3��	��C���+Q�#LW�7�����ȴ�fU<��6����d�[)�?����t�m�&3��� ���ʎ�Bz��V�4{^�@�j�N��2LT����ѣL�����2�٬h��[u]�;��jR�d��6g^��Lo�x�Y�+A5PA����i�<����iBP�N�����swP����#�V��a�6���*���	?EnU�K�da q^���}���'����ALD���}��}qZn�y�y�~��Z*69���?��V��S��8��o���.=����61�~�[��'�S�?�==J�@L���(ɟ�?b�]Rj��χ�~B�ws|:�*6�*1Y^7{D4���|w˺�)����_A�Ǳ�������|vs�e��m�Z��Y���<�i�7���*K����*��S�7�P������6x4գ>Z�p6�y��gzb�<z�%�N�����2&}�A񿗑t�*S��e2�A0m�
�ff4g5ټ��4���rd	��>����� L�a�H9{]T�^���˂Iv��F7O,�H�K�g}\�A�>�ȣ]/G�֣��[F�@J���}G��H�
.\%2��扯�1>�o�T{������ķ�*�RP.4!;���K�5N���C�
�6Hia	w8Fv>���xQ�u-��e��E4�jy�6%����c�ƮQ�Q	�B����Oh�">mو)�uy���
���St�+`�{|��z��h!�W����ݖ#1� O�sI?5��8��_:�`Il֟	�n�/9I�s�B���kt��P<n��U0��cP�R��(���nr�X~���x�n�O���E�'\�P�r��н�s<8[�5����1�kM藫J�w�Lo�|h�,�`�H2����5��kQ����O�fЭ��X���WYa�	0g��'�e,2��m��hE���geb/v�Npe!����Qdz������[R�?\�8Q*������w<9����y�4��0�;�[f��y�~�tn)K�.b\����[�=\>�*Z�TC4�d������u,Hͯ�->�vw�9�9[K�þ�7�M�,������߯�U��C2� �8U�8����ef�<z�� T���*���A	��r����:'��ĨW@t3����G�O�����7�-�SX�W�ٴ�[[�B"���=KS�ܳE�s�ǩe	*�L��Dg.ܛ��I��â�I�W@���y3�U�Ws3�MQ*ڠ���eHwhD��3�؂":���Ɲ�4��２�^������F??in�
����<�lwy!����	��e|Վh��UP
���g��X�7��D���p����C֔P����8��<q�����w�?��	r&Veqbii�Wz�g@��	^��W�o)<I6�R=��>i@��#�?�O\n`���o̗sM簹�䕽����L!���hA���s�Su�s����i,����y��٤XJ�m�WK�J t>���O5�v��
�h�j������J�x�b���~�j�&�Zr�����y��=!�l����ţO]F��e��<S���/:چ����{�]5��	�hU�I��A���n��E���cjWդ��H����4ed	�����G����������Ԓr�ܜ�S�^��ӷ�����V�C���� qJR���F%�0���}�2�f�ճJ�x�G�t[w��N��[�{�K�#�0@R�]UQ�6̀���T�-%,��H��W�Zs{�J���s�78âS_�A�5�}�'�*�X3���,��"_]���,2�#<!�k^��%	�ϸ�x�)#��sl0�Vf(��Ӆ�"��}B���a?%�')�&<(#����F@wRy���{��gf7"p��d<�"�#������屿���~	RNI��ED����V�yz�~����hN��\�9Po����BE��2/�����$7�$L�X#u�p�닚.������d�`T���KT�/2�K�����ޡ���%�0�֑�V�<�ίh�W
����>�w:��`�#��M���M�'�|=mJ�@���=!6ީ�q쥨CT�(�uwtE��І%~-�*��u"QW\���2R'h(i_�<B�~틁��H1oN������V�D���v~>Z��>�qW����&�P��^�˝#a�Fm�n����P��5O�����ثs�S����!d�8�Pfs4�h��ώ��:�c�@�����4�/��s���R׸��X��i�̍���ա�c�FJ'�	ܘ�pV���[��!��q&���͞�}���{I�Di���7���֮Q�.-���ќ5��.yTTn#�j��̠�ą�6��AŠs�®�n�vĻ�흭�}\�Ys�$M�7����J��(D���W�m�/����˯a��l�|���WKJ���Q�/qwy����g٧wN$�y+t��	�Ѯ��I�BU�ݓ�N.���c��e��Y�X߇my���j�7ɟ��J�b.�>/�8��_�~� ��c����siC��*��f+N�LB1=D�X���u�ng�������yj����L�����F>Z�#��yM�C�L��Q��a������leUD]����!z_�	Ս�&*��`H>�k�'-!���6�^q��bUp���� ��"s�=&��J�)+��?tJ;Zka���˅u�A�<��s��7�X���$	�����O| ��+�P8�\ֲ�D@�������F>N>Ƿ�
 I�v;�1�3G���ls��=�ڔ�;ZG!� !�����,A����_v�x�Nǂӽ��C�G�j��Fag�	��2�����Z0��A�[D}���-�0[��2bT���I���������ӵ�]d��9|@�u�~[t���N`�rye��D8�Y�����H �w0�����%��r��xi?��g��ld�K�%��:��r����q��]��m;�<��Q��7e��m�%��&E�f��ǚ���B�K�@
Л}6��&�%�y2��)��g��}���eW�X$F��L�n!�,'�V���D�"{.�$;*��^PQ#�2��=�kXl/���i䅁��6Ƭs0'��f��O��;�W"����Cd&�]S�c��hW�����А��O=������m��v���IN�6��M$��j�"�1���.sܢ�Ѻ��Ⱦ��n�)�8�zLAr��'�=3+���Su�L��!���,t��m��(�YU�['N��^��cl+0�tU�����:�fe�D��6ǁ�O;s�%��
 ��Ў��Se��f�G�I����ha/��K 
���o���������XԖh��*Y�r�?�A�M�ڤh���,)�Xa�FM��_���>�:�tU�"N3҆�20 �f�^Zl�P
���G�t�M>a���&����.Q�n�Q� ����`�����*4M�����=�|�f%�8��9_�XU��+0�A���{f���$� c�×��U6~i��Ks�_�eû� �C�j&��V���T'P�����2���,UV~�Z�YEP$���U?*��zє�!F��/E��<#鱺R/- 5���R.IX6������m�{�I}$��*Q�Ӱq"�E�o^R!��&U�צ�a�?�>;ϻ�M�����4��X���>��G�u[�C��J�%�o��]U�Z��[a���K[E��]�3�+�3�wS��W�/��� 6�|���w�'��f��D�-��0d�y&U	��%59慷��ޒ����8�棠~���;I"*���a\�>�����+�?-F�dC�,@���6�ͯ�5Ў.�^�y�[oC@�|]u��"�;�$�թ��@d �YA�oF�a4��#�h*�^I\��k�H�/��cM��)�7�\�TH��{JZg�r����8O^���3�th\BB������t�ZQ�W�Ӛ|&a��C�j�ʟ�O7Vh�C*X�W.��&أ6��\�5�X�w3R� ��:G�<����=}X�Ƭ̢����h)��W��]��|�W�%ܼF|+_{gۊv�]Aw���v��'%)ٍ]]���"<F�ֻ�ύTm�����s�&�8�>;��3�� �����׊���F�l�v+ ����I�܄7�M/C�4=/[s�*Z��{�Cq2p0W�b.�}�.A]�Ԉ3 �e��4��8�����ɀ5u6�#ɘ�H�m|���c�w�z&\g��v��j��ꌚ&l��#�ĩ(�����U��N�,�&�����j��������4��L��.h���w�s<{��pѤ��TΟY"�߫[ͦa�b�dHG�J�i�����a6�3-�rxR,�c�$EJ��D����0�h���׊F\�ӝ'�-Ϋѝ��I�Y�J��/�g֤�r*ۄypa���\�H\��Z�C�(K��2�]-O����,�ڑxє�t���̐r�U�,�9���?LAW��0J�ӫ�B� �0����]>Zs��S�K�-jw#ٟv�O�*��A�AP��,���������q�E�5 	��8Ta�7#޵|]��q�d��������+�8v^aO�J.Rsu�]���&�Yz,,a)�tEյ�G�C�N�Tp_V��l&�H��������<��[7�|���MfC�O<	�YVN�D ��*�bP�gY���I���ε��ύL�#����s:c�x�5�.�*�!I$6ZL�S7���K��y������jo��e�D������o`r��x�GR8&���14�'\Ƚ/�l0�$:k��.4�Wi{�c[�J7��4T��.i�E�@+R`F���S`�+�zCEC���9�s?�,T[c��5�����T�(�;O��*nI�^�S:�e,�7��"|�vl1��=D[�!�S|��C)?�ӵ��� p
�縣�`0�mE�sV���MASJ�r���,��R�+W9�(��&��"�љlF��f*X��淫���=oj�s8ߔ��0�&��X�ι��6��"�#��`?�R�{��^M����/�,A�r��VM�r�b0��0óQ_��9H�Bժ/�Dfe*\SRGT����":vI��t�8�*� y��N��c��랼�/Mx_!������#���\�g=�"+���5o�'��[3F�V���Ay��)\�޽�m.*hyB�f�?t��`��Ӈy�C��&Z�!έ)�_���Ul�W�1ԯX4�8qn%�t,����f�w.��Zk��"��K��d����@�i�}�W#��-)��9>�k>Z������J�Ypܥ��@$�k:+)Oڎ�܃�I#�΢%? ��'�wyq��l!g�5+��X!�F������&`�&lJ�F��d=���ރ��x 8�M�q���g��r���uӷkh������	�5W���s�Źp]� �@&��Pᤇm?p����]��i�G��HE?5�;��*��
��v���D��<xIٕ��_��� �4j���=���p3�������
{����1��o��iؒx��K3�ϣn��7����q���Bj*������T-�ڵ�#Q���՘]	",b��kƳ9g���\���^m�x�5548%x�G�VD�Ng�F����kcW�X*_�G��X���ǁ��v|t4�7�\���_�I�#/rxigx��PR]���A�I���ݍ���o�BTqo� ��`~���u�2TMQ�柔4g�����xJ�|>��Mg����X�M����L�I��MJ��������վk#���|�M9?!��z�ު V>��F��iܣ �U"�DY>��#%:w�E�h'Fe�A�����Ʈ�Nu���f���?r/�s}�o S�z��Zrd�k���&'Ӑ>O_��v[˹XqTC=�1�[k#��F�q��F�O�h���i�b�/�5����35D����]�؆�V�Mƃ��!�����ʍ_�yIH�s��/Ɔ�����3�M�v�G�$L�������J�?1����E�<	D0���ǔ��CTpwY�u�2�↵��Ō1== ��=I�Z|�R�|Z�*����^��F��)7�Z�79�(ɸ(�O�B��U=��B����](�G�X)/�i�_�:��L�s3n�C�͂�mC� �ŭd���ArZ ��p"W(��@�L�fL�nǆ��,�i��f�fm��n��^nb^vqR�C�f���#]��}fh�NN=6�WfV�{�U�G�(�^��:4���J{��[~u���%�gI$����w�T�Y�H�XQ���I!B�ȡ�X%�����/o<�-���f7���g�X�Pi�6�r��Y�&�N�	,g>�w�����2��tMf֩	�E��%����N��D���.(.C����b�X��Y��@'&��Xh>�'��}g��o��|��[l�jL��3оwN� P���ViW�m�7���׼"��9�o��n�L5
en��Mn���>2�
�=]�g)��TxO������R+W=�n~���ަ�^����$'$d)Г�(���|�CL���ch���Xo`��/7@�EM�����T�v}�_↑$-a��p�/'!��}6I\)c�x�V�j��)��	� ?Cf��%/p�%ƒ9[�Y��z���l䮘Ai�RbJ����z�q�p��ϵ���Es�:��Q�>���+����Q)��^��I�P�N��3�[�״݂�)�}(�*r�C�}��P�1��d��t��;H�b(f`���{5>�����0��3\~d�Ty>#>�v^
H83w�h�W�W���O�/��i7�N[�E��)��O?��F����"���c�:}=�����ˠ.L�Xӧ��n�3�#%I�b%�-2z"y��{�|��H�co�Z���0���7�5M�!��;qA4�2�R6B��a~3�b៦�N�)	>&��~NW60�k����������8m�q��ܹ(^∼	0,F���AN��f�5 +R�+�B��7x�7�N���P&�J����/�VAz �X���&�eV�.�J��M��'��k�*=��ތd�Y�x��ϐ��YP�Q�P�>H�E�� 8������V���3x>��;��R��X&U4VF��a��	ʹ��d�sq!��ȳ�2��Î0x���5��|�H�� g8S�K�<�ns��.R�r����\����b��,���8�L]�{u��3j�mh�Ť�#��Zټ�.O"΅%_zt`_n��0FqP[�����K��9�/�]T�|�,��Eym�^�U5��~&j�t�/�E�us3.jۑڞd�T]b飲O8�~UޞƓ�}���	�����	!7*�2�),Mk?�Z���!��
�����{���a�n\�ȍy$���D��)l��C�)(ve`��͍�S@vKX��`�vPu:�6�g�+����A������<�������0��$~�?,��q�	 '�c7��	~筸c<(���H&�E��t�a��#���0/�qL��Y�N�q�1[P0f0B��$�x'r?����V0����ˣ�&� I�GH	���:�7�&�͡+~%=iFZ�P�Ɇ�g���������u4�M�A|Z����4��.�/�}-��E�5�I_�UFm�i7�gKԡč���� �U7��~�0.����0�W�īae�h�^O�lVf�����f'�%���W4}b\0��R��J=R��Aˇ�}�1��Gjȱ�|�l1����Y�w�vi��M��c��jq=�3��6��9�����,B�Lڭ�J�6�5����\��y�%Y?���h]͒�-3=Jq���`��X5w�J5~�]��v�z[Q��~��<�=%�P��`Võ�W���<	ai_D������\3k��/��UrR�-I��1_C=��p��Sj;'�P{�}��2����TD����\�K�R�!�́�9 DA�:�ŧ._zc/e��&wܥ L�P��oH[�Qv��p�Z��R� G��Lc�h3AQo�	��T��1ׯ�
S�.���kˍ��e���5�֋�$d-���a����'/*o�ΈY,�(4�Ƨ�ᵝHr����'�����{�	7�ҫCM#!�r��YU��ݨ;�%����LX@��D�1����X�d�\5]��>�#�nއ����x̭�6\wߞ�I�=�6�E�0Bp?вfn�d������u8���q���|�����~�Q[ւ�dd����!;pK�$� �S���4&��,�R��Wv��P����2�5�oI+9�d!���t�~���#�kC��(�" L?�n�\����Yp.���aw�@���e��k�b�lI�Ύ%O����7����a����u����Ck]�P6��\�D�$;o'�2C���H�1j��)�l�+s�/)I��Fs�3ι�o��\�E-�5�]�1�>n�FCN��) :B��2nP���+��:�'�G�z�����A��5GkFN�}�ZE�k�U��0�uR>$��P����y�����yĩt��Q��Fұ=���j$!ӒD9�KLR��w��.=�ď��v$,|�З���an^��L#��7�S�9�j��SJ[�Z���2�X�.�["��~~��o�[�w�L:ܧ�o���*�,��#ĦX�uL��X�NJzi����Y<�q��B!�"��.�:Fߑ�]w�uG~m��>a�V_dS��WGUY�嫾���]N�:�����YU\W�E����r�.�¦��B�k��ꏲ�`���oĒ*�$R��,�o�������@Wj'⃂�%HA�]��F�tG;�R��5�j����90�L�d7�u�L����%
{�1s�T%\MEL�t84K�;z�s>��5�y�)��Ӊ���r�}$�r�#R �i������,c���[�B�A|�|�u[!&V,q��
����|�g�Ӝv%�*��~[�[l�?���my\��iO����a�@j�Ҍg���}��^t��ҡ�[�/�6���탒���@���5�V*�C�iT�L�,��p�YM�b����n��R�s��5L^mO�RNd�v˙r���$w�t��5rF��m)/X�,�_�jmZ�R]3d��x=np�7������ʐ��9��y&�N�=kTIj��(�����Ò���t��U�۩X���?�T���ǁ>7�I��+�иq,�7�i`����\E���t��czM��BM�n�f뀎���W��:\������N��~�����Wۯ���*`�j��#�z�qʐG�?��E�V9�	��zՁ�$����I+��XiV �U�ި1��Oq}i�*/��!\�.��'�$�kF��G�w	)�j(�� ���k�.`v�������Ū��M��I܎�{���z��8T�^ʾ�"�͝L8\qA/�����bJ��&�*�O=\�Hk�����|-�('�� ��~�r�8t�]y�EG��]�ز�҂vvGo�C��=�������v�؎A��Y���ɺ��p���o@[��ׂ95xB����3C��J��ǉ*�duW2�fPZy[���-��V��L��7�	E��-90��"��m4X�C�;�`������x�� ծ��,{c�A�_�蛡�"H�X=4��y��7����T#Zs�� ;.oޛYU(�u���� vOv�#����V�A}y���fD�T���m�P�ׇX�R]�0��.Um?���<���(�f��#��q�,�E@�׷c� tz �x��H��s�b�,���;2��5�e<a'\�%W+�+�o�^+�'ؑ�9��SA��\��:T�lzW�����T�A'.�I���LO��g�n?��3�Y���U���Mqm�Q��~a�[�Q���W����,�U�o�j���v4�ܣNJk����2��@d9/�1�6G�\�+薫��ֶܺ���p���p�sUe��E���6�:}ZM�Y���k0��qB�*�p�|�F~i,��e�����wF��AA�j����h�Xl�G�l.��y]	����y�p�;yCRY#ex�c�jb�����Y���k����*=��H����c�M�m���O�ć�R�'�?�s)`�v�/�&u������0X̖&�fm?��uCr��:��z�֕����h�뻌�?{��lsr���`���5�����:�Tnx�6�tN�p��"�m���ʅ).(1B*P��l�b~Ƚ=fn�ˡ��J`o����j���Q�s�7&�ScY+˙��#v%7� 	���K�p	�V�a�
�?C�S7��;j��3l�n��;+#��3k��uф>Ң�Mݴ�04��\��G}�� o}�ӓ�ͳ�M��%�+�Ch�O�F&�_�jp;t��+SX��?G�M�G�(�9�9$�hl���L>�v�%8�V����T�t	2�ߗ��5�r�6�Sw���p�U���7+������T�a��"���x�7�ebX��su��'u�|�^�bR�������G��-f��x�﷯�)!�߲�X .{-�Α.�y�([�� ��D���"��o���)�Lt)����Ы�8�5�������_����FY~�CY�}�Յ2�n�&��ʗ/���
5^�.�ۘ�f*o��;vƢ|#@�/z�R�M���'���������pk��U����͞��a8@�����r���r�S!TG�5�+��m��İ[�"�!�Z}�l���Õ�\�UO@׽0�w�0L�8���v��$�\�(������ܶ�g̏B+�]I7�Ԛ��(���@�Y_ɉ����K�LVu��sU:�d.ڑE��*���pMŴuW�3�����矢 J}� 3x��O�L`�3J	Py���V��T�0UP3�6gUH�Q���q�ց��N��m=}�7���)U��E�MM-'$,��P-}e�-G6�L��7ۚM���q��x�
�'�.��U��W9*�[?�,�K�p������[�o�#Ek�eZA2xi**b���P�|��J��ҙ�%e�g�*0�Յ���b�!�{2�_=[�O=�C��Rd����r;����Q"���Y�t�G��9/g"�j�R���Ź�J	�����'��_K[��".a���z�Xά�DZ���I�N��귧$��_�hf�@���8ER�bL�eE�a��&�^��_T0�gӍ_^��،�8C3�-k�ϫ�Gl4&ь` _,��������	���ߙ2�)�W�o��C�X���Ǥ�ݦ�����Ե����h��~�(T�'vA'rǷˀk��h2}�|ܺ~�#�T%}�si�+yH|�6M6��V+r��g/�'� ���Nݲ�����'k�*��W M��$��/%�q�0��%�b���׀�¹ږ���P��S�p�cޠ��E����0	�A�8FȤ��C�$p�m�*t�B�Mp_Y��$I\~4�sHB�c���i����	=�� F2�m*	̽o�!\M��dZw.������U�8��N�[�z����fH'����t�)�����,I��F	�?�����Xbc껒4ԑȻr��y�c5?���)�j/����6���ܚ��}cY�3�ggDt�Z��	.��x�_���SlL������OƆ\�{7���_yy�߹d2�kO�;��ȥ�� #H��;�I���vc,H��L� �΋4�Z�/rH��d^��I:�,������=`�ӗ�!x?Y=Tf��+5{�Q�b-�&j�������hvA�޸���2��'��TQh�
�" g���>iq��Q�b��AyD(�B�����>%�ڡ��=�G�m�Iyc��/��?����k�*E�q~�
��,��C���4W�b(TJ��fh��"pm�,��H���%�O���J��}������z�`�жFo>�X.a�/i䀑�1���� Q��1/�$p[c(���[�<�8�k�2ɗ��0�c'�ϮG#�����ۛg@���L���W7���p���d��qD��]���~.�C�Y}�%�oC*U��|�#�rbD�]ƝB�q�`�&�%�u(OC��/�X5.%v��u�j<i|����"�ޞ,nb��8uy���# �k:����t�XV&�llyN�2�L0���E<�0�cxc>�D��N����aZG�Lq�y]kF�etP��߅�K�A%�؇#CH�,4I��C��R�7��_?��WhF.�i=�-�	r��
�������:恜���XaqX���c�ջ�[Q�	Z'���ـ;�,{{M ]�ym��1��u#$��mY�� Īt���o����t��q�e�YpI��Vg�=�������b������r\ �O�q�G��0ۋ#B�̟�`�l�$"���z J�T�B5��g =�C�s7C��.W��ں��|��raܟ����8�n�Rl�H��9}��d���}]�q�����nV�/L<�Vԝ1U����pqC������+ѝVmG�a��{b�;��`��R�����'�ᰚR
Q�*�8�(��f[�t��A?�L�.��Z����-�gj�F;����(����fJj�0��aEe`���Օ����a��#��A|�磯{Ǝ����$,�Z��߂͸���t�@9�Jyf5�EƓe/3Ƈo��hmi�� M]�Y=D��_�P�nly�B��}0~�e�y#��[���勃��� ����R
���h(H0��j
V�>ʏ��g��P0�9����v���^N�&�D�#�5V�������}���B��̃;��Ͻ%O��>���t��Yy0�b�Z��aaTR3��w�
��Py�#hbC�?
�<5�J�E����9���'�Y���k �N���u�J:��� b�*�`�`�=����}�ê#�8�''v��e��N���~�.�No�H�<YY��-)���wu�-$�HR��c�(�k�Y�OB�{��Z�(�
E~-�x�����RR=��۶�0T��"y穽�GK��	���CJ^'1�J���sG��������m�I��%?k*1�Wm9&��R��~� �xB(�]��
�	�_�D�c�v���|ee��+2��5r4�RC�X)�4f�ݿ)Im�eE�R	!��*��=�X�8)�]���r'@�Wg���_Dhd@ķ�N�dB�V�����;��l���	���C�	�ꖐ�L��(L��Γ��Pq0�-V���n"��a��q��f�rOX�aM���m��.hT�~�y5OK��K�g��Pc�O�	0C�� ���4���P���/4`�� L����u�f����@��4x<��i;����{��~�?{Al����s��!QW��wg� ��d��t�Px����QF�є�ӿJT�U��|���BX�k��デ��F�9��x�*�v׈�ێQF�5����.��$�
o'�/�6p�̬i���4��,�h�������6Qݬ]�5�z�d߸}��0��)BVRN5*g ?�<���l	ܱ�F��=�S�}*��A�EZE��%"�v��n���+�����a�C'�iY�	�O?�T�]�Զ��Z[˰�f���ݖy�9��J���2�c��1����w�.sy`:�d�0D6_F�� �O��T|h�����Ͼ�{��(�e�.�cc����K�
��>�]� K�a��{�Sl��H;�#����ea�Qτ"dя����v�
+%�y�R���V��B58���Z8��>�~M�4���[�%��Ͱ����W��z	r�ޥg�\~B�yXڽ��l������+���U�7�*�^`QIuC���=3���(f�~�ؼ�Ӛ�e���F�5���v��S���}^=���U@�'�;v6��5�:oLe������5Gl_�-9�Q�߾��I��ĸ���L����ƿmC�$Mm��*ր7�/(GXKyq0�f��E�b�&"�/�����+z̻�T$Zc��'���f�<����U��G��jz^�|lq,(�_h�=L� �,q}BT��+��Z	p�����=h7F��^�k
�.���Vh�a�8�\ʵ���Mk
!˰Ξ��_�4Xy�- 4�"����3
{�����"���R!w"�ջTT��{�e�}MR�҂����*�]N Xb���AR�����I��A��J�ɧ��:��Z�S�P���z���΋er/~`��t��9G��7�l��f8�:���Az�J0Sl��k��p9���:N@�%�U+�LS�Eb�&�oq�;�q+H���
Ӆ��M�N�� b���ųq�9���#��IZ�>�*����Ŷ�	��ir���1�%Y�˸��v���
��
̝��4�]ب0ޞ(�F�3�%ȸ�$���}��p�.?�Pc9�ݤ٩V���#h�':rԬDD��4���&vP��`6�ކ�^�ۢ�<mX�˪m�I���78Xxo2���+;��~�q����
be�w-�ׂ��Pf�H �����E�۟eRWj)m��:���0?�I�Vn���iw����|����@f}�i.XLI�#�j�q�}"S��x}�W�jK�ʹ�I>�����2�\6Aq�����x2�ô�(� v�6���ܹ��D_�|=|��g�O���N��d�A����1陡�0w�԰ZvA/��I�P�b��11���\�$Brf���
l"��@{�5O���e�rFX[��ޙ���D7:���f��M�T�q�]�� �y#�jyl:��)�����JZ7�T�g�CU�����,O�Ѓ����n�$a��귎��P�-����_ٴ��������͟��@wn�ý���3O�fB�'+뼼�a��g�`�\�j�JM �Ȣ
�P��0%UNqʒ�O��Q2�Nc�a_�$����|A�Z�C�����g�2W��@S|�����-��ĪS��>��H�����²��ub��8��@
��<��t�s��0�qv�N�ظ��ɥ��)�[����4=�N�:QSE^���+3p�\(����U���mt]�>�9]�K���T$�:�0���t�����IE��|�g��[Lfq�S ����0��$I-W�VЁq����r#�-�E�'�t�;�W>R"���&��,��S����+�xF�����xS�B� �&~'BG�yiOoLU	8��4p�LW��ޖ����rt��T=�U)}`��Q��bD@�t�^��
�5��=
�[���eB�z'_n[?~%�n�Ռ�Z�Ҧ���̀��0k� �JM���v����� ��<�m	qۈNͫC��2�7N�&������Xsd�2�����ē����C���o�\�u�%�3y�[����j����hN��!�x	�&e�Z��$"h���/ʲ�KĤ���e;�	�Xpp{���a��V���Es�5DV���V΢ݴ����W�\�I�"��t�o���� ����~`�q`�tԸ���;~+���w�֊����+fK�dXrvi�!�BĢ%�L3�j����C
J9��\�S�0�g&U,m��l���uDU�cڮ �-�L��F�(^!"�T��0-�� ��)��gɚ %`q����ə˘�S,����?��R�f�eѭ���3��5-��q@<S�e�Q�~��=rR��^��ν?���e������X��AT��>���,/���y%l�e^��D)1�9��i�+{�|�w��XH�J��(���$�:Q��>�٭(��0E�*!P������6�QY�1[B��]g�W��YM3 �����7wo����q	/۪�z=i���U.�L�C�d]=^�7�uG�B�C�-؁������~���H��2��MXc �P,&�;y6J�V{G�j�����A�ʂ}Rp|X!��:���A�������tS�%�^����R�:D��#���ϟ�B�/���L��c&����8�T��v�;�E����O�%;"�z��%T���Kz���hj�5��/}1��*jb��\�]�=w�ň~D�RE�;D�"��k�/K-��"�O��]�fD���cxD�җ&��]����rW�Nm�j�h������?(z�P&��ĺ��#a��
wMa��왐'�hݯ;��_�'����\���}W�#�1�w#��P1ީz�`q��gs�i�ʱr^/Ym�~Oj�+&�����J8����k S=�&b�u�ݐM�i�e���n1����b� ��<�6,P�b�f|O������=�I�)vm�>`�ao�+��:��3b�A���] S�u��y��G�M���U�C4�w;h9kaBCK-OM�&`�Z�¿>��P���F~��շ2�Q����xh�{��mܙ���79mG�8z3�x$f��Ȩ➮��I��f�C��i�5�m�<�-Nf�f�̓������	��:ґ�G�Gc�-��!�	�w�#�Zk�N]"�a�<��9����'�~�Լ�H5'�&�ɽ�Q���㝂c�<�D�ӳ03�Q���_q�nc3�*�_Ga+@re�/ЭPXp�@[�[̭�S{���A�=�KcT���Y]�� �sxi @6uiBWF��Pl�N���@�����Z\.�	��Anڕ�xx����X�����?����GǬ<��|&o|���:�ܠG�d}V����=(�.�Q���3	�q���R��� �7�M����v��0PoPs��9�~ߟϹe����.*����w�|��m|E�?�N���,ZM�\�	�&nF�up,�B�n�n��9�Jy/��胨s�@t��OF�1�o�G���KMC	}�E������>zy���i���z���2yz}���&$�m�n��7��c�����v.>�l���,���%WY��-�A��{��E����*��.�+~��qF��(u���RCHGF/�/G�ՃⅬv�yp����!A�;�m!��NBER���R���I{���4��=k�(��i��2V�dD�����ڋx� XX�Ï�X���-0A?f���ϵ�W��p��a� ���A=����8�.�U�0��P*P�J4aM�TFT��@�$� lA.�LL�h�� O�Wqka���P�u��M��G	��]�p�2�6Y��hw/F����y�V�苺�{/ȁf͞�wl�a�Kۢ��C���!�^��$����m��@[��v�\'A�fޓ�N}���!$�î��l��:�ӭ����I9��	���W�K" @��N�<ϧ=d䣐�l�F�5M�>Ze_���C>Q?�S�Tw�`k����@*�Rh\����������I[�S�J���k�q�E��t�KD��ھ ���[~f�G�QK��&�@t����O�:꣱W͕^lhs�)�$����jHyn/���J)��������W��#2�h�>�i��j�����������<H�.��7�L�d�C"��67���-Տ���ӽ��T~�a:��aD�;���lfr2���SG3)�����Jց����yUry��n�j�Y�Yi��3�RǶ��e�����"�TɃy9�U{�m�F�����)� ��c�8g��yZe>�H��W,a���(������= �L�Z��Y�2��[`I����w0���T"m�z�!�sad�
/���>�*YVK��n��S�T|���3|��w���
�V���W���i�>�v���,��^W[񆕔�0q+��F���/��n��R��N<��j�]p���N$�E�ΗN�1H�V��!�HRE����-����XL������AM�s�fF{D4��j��/�*ޑ��U*)�D�.�a#s���B�2����l���<�_-��!_.)�G��ZYKg����l6�3*��`8[ɹ�����z�����e���t�4t�f��M��ȉB��vdR���]��O|[ŉ%ϾS:E���%j�r���I�(WlA�U�N��BL@ҩҾ����&*�)7��G�f�*�P=��}Z9g�`7aG_�0�S�b+R�Qo�����Gc=G�ʀI7"�Q ��Y��	y#=��W���j{g���94��Pʠ�b7Mū5����GL���.�"������i-U'�p���i��K^�m��@�g��FwIPP���̛�G��5�5j߀���������l����x �怷�0ti8��K&_: {�%oR�?��+]}S�u?����p�5��ػ�T������Ʌ&v�a$7�.#=a� ��^@3#^���qz�FN H�T���2��r�[�z5��I
"�E�����|nіViC����RSޤ���p -�.3�)
�-v�W���ߕ\�A�9!r�h�B�jk��,�-�������Do�<�V��Ss��DD
�*���t����(�vTh��V���t��u^�	[�zZ7km���%h�4O�IA��󦐏�?�����U�oP��$�ڳM����O��%dӵR�u�{��^�O{�{�7f�i�ù����V��'9_,S�]{�t�&��+�2�A�]��}w����͑��@�̷r?C��qH=��ڴdV>ho��������#��ou}=sD�b'�ۀxR�g_�Ҁ��p*�u�~�	�Nx����?$񛴊9�A_?]��<��]ZK�U�3���eJ��ܶ8C�����Ź0�戽Z�mP��Ykc�X'��~+��YiR�-�]��-G��$�!�9n���2}n)j�-��5Ϣד.�/k�|F39�����Q@Y�8&�i��O:&+E��f�O�o"����`㥎aN��3.9�4�`�gԖ[���j��򶂮��?��ǳ�y7��h$�^*%ۻ�48���i���}�d� [��[�1�(����X�}��K���al�����f$�t���-4"�H�w�;�W�S1Wb��j����l]������p�]8o��c��y��o�;���:�$�UM��Z�$���)��s�Rz���_�q��D
�uZĨ]�7�06����5��'�4E�Dn?�a4Tn�F�js�3���{n:_F�"AT]�x��g�7��oHߖ�qr3�_X3 ��B���X�Ye����<��u���I�
��?�c	�p��k��̌e�}���o���W��v�#��;��˂rr�g�vU�3B$�  ��
',��VL�O ʟ\d����kh�?>�g%���zb4�|����0�E��	u��C}�ݭ@��j�M�y�;�Ua�O�1m�:�:E{���X�a�R� ].�#��{���rN;f��1�D`�X����\��nj��(��8�@��4�k�a0Г�y;5��h��w�\P�:]��i}Ra�&_	u�L���� 2�Eyc�ǻ�Ҝh?���V=���/",V��8�S_Z�|H�����1Z�!Xo{I$�NN�&�G���U�Č��XAЄ���7GWPUk�4���+�x-y�?��K�7�T8^t���	�S[|3Bd�j��Z�p�b�-��*\��{t�kt�(������5�%p]�sZ��{(uO������Mir�5c�qH��;o��C��N|�	'H�mm�O�i#�M��[Du~cz�z']2�p#����_G���K	q(����Z)�@ԥ� ����q�<�[�C��mF�@uSW����܌>Ѕ�$f��&hY�����!���ʴ�u%V�J�N��`ޥ�Y��f����(�F�ܕ�CV�V��b�\�K���v�賞�E9��:���A� %�.�� ���"Ć�D܇�W���n���gCv�����q��?����F���4D�^��ybʛ��.'�����x��#��S����;Ȣ�c%1�+�%?��e���l�W�n#M�P;�nvM����/�*B&f5'S;h�k��k�	���P������bQ�n0fαك@�b_0�UI���![�⠍f��,�C����f�����g�h��A��'xs�I��p�w�@��OG������Da��n��Qy�r�w�Y�<M��T�)��r��yu��"�����X,u�20<@s�u�>B��G���{L  ��/��7��M�/X�4�\ �1����@�C��7-�+���-��^�}�F+4`@Y��֋}p8�R��Y��*�K�{<̳���$*�(F���Q�_X#� �`�e؉��j1x��ѻ��dU��s���"�M2̵7��ĳ=�mCv�b�ѕ����'��^��_T�F,�H������)�����"}J���=d3�ő��B�w~�	[߆���T:�}
n����7m�cO&�"�XБ,.���!�M��̆������3�?�j�y��7������||<�T_Z�ci|�ޅS�h��[E��τ��l� Ў��	��
�UN)I��	C��b���P޼:�<l,���S	��O_:��O�|����>�)����)��})���%�����@UఠF�S�,���n���v@��ʔjy�$+m�HT��wB��d�޾+�I>����yo`�6s�{�+��aӦ{O�	)ǅ>>�����&Ɩt楔w���`Y�e�5����F������*����x~{����ێͺs��q�bh�/�eb��2c�]ay�����Jvd�JF���?qP���Z5��D���FԥU�4�H�K"=���p��Ȩj��~�k�XsU�N}]QF�eA�[�j8�hF9cIW����5Wr�9O�>FE��'���A,D��(����}��O;������8"@O[?�ls�x���FңR̥eC����`���Ź�/���Dr��F�(�&vE���$W�������ts�؜;q�ΣsǙ��>+�ٳ�"��f�L)ιK�ߖ'���T��8������P�4�[.NJ0ǱͻS�-{��rXvdVѲ�z������`�n�4��l����0he��\�^��b���̇�J�Z��3�uP �s��b� �o��)���oYMT�1��#t�m,&l���DԐ�gd�x�,q�	� ��P:Oۮ��p�q�,�&'ݪ8�T:���:[zV��a��R�`Α���k� �j$���t�D�4��4L�42�Pix��Gx?�=��L�L�#�^������&%{礳��'٨�9w���>�2��<,d��U�~�׭#��sV�އ��s���xu���J���I�@L�E	�b��~�Y�[��M��擈�^�
�w.��6��2�]������E~��C׎=��+�G�h�o�Z�)E�}A�
w�	=���댣�5?U��,K
#[��+�K1����z��(T���N�*#=������R*�3!���T�K��Ma�� ��h���m�#'J����c�x�?nG�hV�Q`���X�e�WuC���!�"�TsW����"��S�W<ģ[`��ʡ7���P'�e� ���kk�}�f���+b|^����͕�E,��O���;WY#�6a�$A��L�3��6�Ez��.�c��?�2d\($��ʬ�x�D�H�M̅�i�͇i���;XA6����֨�>��.���K�ea�Z�\�:,�R4Ɍh�^�]�A97s��-lՃz�.=6�{r�rP�y������Lmp6� n���c�$��#�pw�!�6Q��o�R�oo$��[:��H�����A@��*�.�r�u���2�Z��ƞ�������A"R�Y߻���׷�+uz���C,mo�hy���[`�v��2_�6��w�io����U�-C��h��So��,���|���Y~��`�I�hx�[�G��_]��_fe��C�s��孫
x�hK"q�&�4J���$9��c��3�|PW���V
�{����}��'\����Z�S��z0M��}~��Yl���>WlB\3��;%f:���^�Z1�r?��+L',��[H��З
��#Z��4N��lq��.�O&�WO���vH�0�ڙlC9T����I]����o��������&uRW����e�d�Kd8C��&����>�>G	z�����N-2+J�Q)z�W%��>Q?�\IA�=�6 ��wO�XF�D��E�z2���V�N6��ۀV����0�!?�������X���k�̡|��[Er��)l;��}KWz�F����[�n/�����b?<fsO�]�5IS.)��5Ь��[�~g֍h�}h��Q �'����xE�)�^]I�t�/,�C�f��� �,���hQ��\V^7BN��j�T/o��� :s�㾀H��4U���1�;V�?��V���8:6ղ����Т=llRP��kA&YsE�V��2�KD~8`�k@yS;���fԭl�4���������8[�ɵ	�t���r���f
����QBsnC�]7������)(��WA���TW���_|�Q������
�~�V$N�!֝SGY9.!�|�'�������ugs7V�gp'�C��}�iueE��?�C��o ~>%������
��`k�h�Xe��"��$�M)nߋ�gØf=(t���0JtR��c��<��JwB�[Z��ථ^�^�q�s�9� M���yyȄ�n8�t#�%����1����l �pL.{�,��µ��א��|��TN=�bM}b �L�-R�
f��H���Zo�F?��5r�:��qxjt�����1\�O�ɋ�� ��qc�@^�]ˎ�	���άD���{���H}���>��XI�h��~� �W+E۾��N`�ku�>n�O���T"�2:Bb�B�;���7t���D'�gR�a�0�]X��E?6aE����/�'g��sB�ǫe�����z���H̳E$Nh�Q�}MRː����,��s�e��|N "��(�p���n�d}�KUS�2�5xZQ������Tܘ��~/ 4��a���/e�|��e�Ȏܯ���$ARt��@���T�!�̴���L�E�*b/)'H�W�ī0�q����W���O��:�ҍ�V�{S�����b� �;NB�=a�/�uβ���f�H��s�\�vH�
�3%���1p2Y�w��ЏUG ��L|���(=^H(�0GidR�'��g�]��������������+CW� �%�N��j�j���c�����a�k�4�����c��r��ߢk'ԝ��,)��G�
��p�<�聠Q��5YE��d�k�*�a?�/-<���W�=6���Y}�E��Do(*W���[�s9���^�rۦz�rnCܸ/u�?t��MOsX���\�V�Rq#s�MZC���OqL��OԮ*>�/��C���	����j>/��fi`@c�%��p�2��:	+��7>K_�bJ�}�E��b�r��)�����s���4� �d�^;p�Q�H��M/xg��/��@S���ա��ZQ���P��%�B��v:Έ����(K�r��+v\n�2��@�N��ի�u��Z��Qnڠ���g���W�Ћ�$A]�0�?Y���?�Fͩ�䖃�*�z�C�7��;��`�	֪y���>�X���>�/C^G�Zpj�����F�\��(�J&1�ȧRQO��ܺ�-�Rc�	Ao?�u2 ���+|����`��0Oo�����̥6j�=��IJ�1�~�T�q���P�NQ�<�����iI�W�S��>tk����{J�wվ�����,SB�A ɗb���.N�F���>��Ӆt~��<|�h�?
���9ɍ֍��Rv>x*��܉���$�|��Nޔ�ȥ8f$�"�@al뇠M�h�>8\\�QX̼34�{|w6��#bΌ�L���6��x��9��Ew«�-P�M̍w��FA��ϣ��0��_�0���x�cQZ/�Pz/G��'[��dq9$U|�S5FF�ހ�GR��dy<7�v�q<��Ka��0��Y��dh!��$O���2�B�'F����p�:��ᑙ_Q!^�/���<͊�]w���M�O�4�`:w;�# U����	�˟ƒ� Q���Bm�o�|��F������񴺭[ٍ_�<�(3u{�/��WiD�j��/��A�O8�Z��L2 9��O�[n��I[(�F�2�a���	Pb��f_�H��rg�?��4��xϾ0��0� �:��xzzhC[O��|��!���@�g�f3�����N��[��
F�L�����e/ �����2N!��6�����b`�Q��Ǿ]�F�ߩ����,�&��U��Ϩ�e�8��W-��BpD���IY��zD�KB�����6|yݿv`a+�+3�8���FB�9;���B���TZ�����U �^3��վR\Y���b���G�C8�ͦ��{9)8���r	h������*Tz����[�l)��_�d���b�/��\{`?4G�(�[`��_'�Ç�m��0����PB��m�������Y|h���;̤�����d�J}N�]�����4gۊ��J6�rY�Ű޹���۲���!�㛠�QU7��Re!�*'�/*��!vhm�9eW�zbpؿ�|�p���:��G��C2�s-�X��n8�Q*�s%hS.�� F7"�%�S�X'�J��eQ_�� ]��%�>Ѐ�ٛ�c`��үs�syZ��� �0ix`z��%�\/]"A�>�Ҹʊ�����=~�}�;���%��� �KA�[6-!H!��i�&;�"}��"����r��<���;"B����F8����8K_|D�~�Ѓŷ��򸜉��P��f'D)���(U�<��j4ɲ,�� IGʛ���]z��}���]�#_��ƨC`�FlU��+��z�W�hZ�MQ�=�MW�t #��3x_0;��bX�˧����E��L�b�	ƅe�|�AB�̍��R�P�n*.�4�#�W�$X����_����-��ץ��P��]9=X��S{髯����m�>+s�u	�RƝO�sf}TC)-����щ����c%����Tt,�1y�����Rq��U�����_��ٸ���:E{gޞ
��n��Ou8A.i�Y�Zb�.>�vn�2��jک��L$8��'�K��eze��K0�S<�
��+@ l��S�L����oDdF��xՐ��uY�2i�u���q�[�?����q=��P�-i*˝�x����Qz����[���7)@���Ս���BE��Xt�R&u#�{�QMe�c&a<F�Ϻ(�s( �?�B�3�T�SЌc���m���
%��چ33N-��?�o�M���O�^*靗
h�<���[k���¶�f�֮�)�H�E�C6O��,H�_�O����g9�*x;�K�ZI�#���>�_0�`�8��������ÃV���;=����l��텎Z�L�����������ny�v}���p{�!��)��	n�4����[��q
�@�06�CRp��j���=k`˃�צ�rn�����_ń���6����[RCz���F��8�!��m�(¤��r���{>�ȩEփ*/vz|���"�DH���j���H�c�����������z~H�����df���7�c�Qdf�"]�4�8.~��Rv�Q@H�-8썡�?&�5���ǓFL�_^����4e��z(���f�����A��|ge>��݄�a�����Q��ܢBb�I��P����a'�h�F-\�Ay29��`��2�͏�~p��ﶪ�ە�F2��e7��D?��9�tQX���YH�)CXn
���o�[��*^q�>�K��m0gº,��|���1���+i_�s]��K��L�R��E��1c-�2�!~�h���R �����@�������P(��!�)gd��A-�g�1���Y���%��0h��Yh��Aϱ��W;��x�z�2�������#8�����i)nkm(���X����,��}	B�bȉ9���۽aQ��с��\VՓW�CYH��^m��?@�	V��,�8��ڪ{+f���"�k�#����%opptg�cn1�Cƞ�칗Qmc5fv���$ (3�O�1�7dl�1Ț6;G��l���gƋZQ	d��)zh��9�sk��-Ӓ�s��e4$bz���:�s]x�K��}�#a�O~�95i���	Т3����{J_=�l/�T'>���\)A�w���Ov=d�߷ ��w]96Ŗ��i�b��x����, �*��<Tb�2< �m��.ճv�,���(��U�%p�t�Ӿ���|z�d@�1_�@l��U�{�,F[�W�$({�Z�ؿ�,��Iɫz�DEeA��`-�9�!t�7�l�C�
�o�3�!���6*�c+k<ڥ�Swf�c���'j��x	%D_���[��䤘5�u�T���b�	�5+�Ґ�I//y�<�_���*h�
�}YNsN�=S9��h2�okY�)�`\:��02���>�q�%u��:�f�\:��j������Ҽ�͚��Y��7�na }����"�y�W��"r�
?�&�|r6@�7�?�ǆ���vo����"K	�NĽ .Űw1���IGھ��>��F�G�m��B$��,e.�Y���=#c�t-��-4��BPv~4D>�����52`;�Ml�xZ�R�ɼ���.*�B7�\�B�jJf-�fF��Y;ᢒ��&�>�-�e�:�4�{��Z�y����Fi��P�z.ۗ�����v��'#͌ǘ/�����R6���d|�k�_n�x��m�����(�VL��;��	Gل�؄4b@�� V~�� 1�V�Z G	Jx�v��,=?&^1���W~N6i4�O����3]�M|ڣ<C��R�
ݶȧ��OU��O�thg��1O����(�qN'n��?��n<�������ql��iYq��l$��`9ġZ�Z�n��u_��VM�����������;�O����aܤ��X�E\�"���S�\^����S�E�l) �ޚܝ�%q�"��XCژ�G�0�F�s�"T� �W;�����k�0X�b��,�O�M^;͇���%Ҭ�E����+��=6�p�������	b��/и����(��]X����e�*j���:�W� .?�k4��F�����I[�� ��Aܻ��V���~��X�LVT��C�6O^�f�L���0�eC����5��s�v�۶�cڨ����%b&����h(���Ҡ��H���d��l��l��m$?���Y��Ә�|�CݘmP}��)�����Ey��Q�j]�{�6㗵h�pnߡ��7���ׂv��kP��$�Wѷ��x���T��h:��Umt�\J�璏����.�6o����g��HS=�_���
����ޒ���'D��ȟ9TI>w��������g�R���L*�����F��'h�J L�s���1��W��"�V|w��3j̖��m$�T��1�[����ǃ��p��ˋ��������a�L���@c����L]Xp�UG���.p�2���|�qr!Η�1U����=)}�!V��6��Y�n����~�m<��A/"P�kR��:/[�虆�����j���=6�(���^�ƫ�r�I����Zn�u�ٻ��o3����Q��n�r@J:���B}���1@j�N>!"�Hh��G>pl��2�L�ͮ3he=�^��Z�h�㖚4;M`'�4"����*��T ޶����w��/̬���:bP���^�V]m�f���C�9�=b,_�C�X:�Zٌw��j�W����M)Җ���@�Z�υO[�����^�:���ar�T�u1�ū�_���!�����P{��{+LJ�~[Q�S��	���D(2�B�ɮ�l��(@(�R$�[�@�Y~�پ��t�3��dɲ�����o���{f����r~#-�0��X�YN��b�z�K�I�{��?�N��v�vX_z���T�����P,�2d}돹�}ޜ#��VI���ٽO�}��i�'�K�ƫ_��\`������T�G�,سKbE&+�pY����g ���L01�?%�'5���i��T��y_b���E케Ʋ6�֗�Qߙc�'>���6�?�, 4Zq+y�+�!� ��޺Z,Mb��_	��@�yoP���:��E�?�4sM�b����^��ie�v�#j �H�C: �v~s��r{Y�eÿ���=�H��E/���89P]p�d�ĝ;1Y.2Q�$�_~z�rnL[�L6��G߳�m�]׀�y_Z�N�^��T�=�x\�/�-=�M���o�0ֳ.�Q���òO����
�2���ݙ�\Z_����h��1+f'&.HY��oK���7	5n Q�Ⲽ������W��lO�-�A�@�nA=���[�%�<b��������e�;jAG�U$�>�ⶪ����z9�f�t,H��h���jj�4ȶ�1b�8�-�d�_ߦ%��NQ�9Cr����l�z�^��uf+�&V:���s�ܽ���6Ȫ3���3zmПQ�RX�h_��i��Б�=��f��~�Ǝ�~�0�]/@��1E\/���,,ϣDJ���+^�\����_x�&,ʾa���}ǚED#�=���k�d�@S���d��F_����Fŕ,�����p�C�I������p�Y���0��;$C�!�w!1-X��(Jt���(���rĤǖ�Z�B�b��	�^D�� �M=�L��l輇�q���@j�YgC��W$������R�kV��/cϒ���Li�s��*MT�n�h�r?�v�e�-;�okn��	���ʸ;ae�g����%����hMrfr��EvS�:'ɭ��r���I5)�y��:�fз͕�g���3m���?�<�"�V �?Mv���z�?�v�
�E[����M����v�ld�A�w|o���"�P����n�:_3t�뀴"�Lia6�d,r2ai[�%H
������诮�dd��*י-3h�]�[��S�L��X��v��W��S栏%GTZ5a.�L?�ERg��d^Ԝ0)��E4�g�w�N1X���s�U�������APH�6�Z^�Aw�i���;Z���d�4��:2����������QGBl���+p�^�a\\ߴ�D��{a��+	�(�Z�&�m��ͽ^�ׁ�����g)j�I�eԀ�a
l�>��!4��Ef/��N�A�:�d*�y�_��h˿�Y��V|[��=3 +Cu�{�=U�\�}O��t��M�n�#� ���Ko���pWb:���X�'���(�]�P���Dn%q[�W6[�|Xe�`$������}J"´��&�`�㩐��k�����S�M�����>c���c<&�M9r*���VN�MW}=�����D�:W�)����� iX�)_���T�D���F+����m�k�N����*5�vN�,y?����@(K}��&�(���V��6v����JD��*u���?j����3t��*�\�9�ޏ���>i�z7���݇7�
߱�a�Z�[Ā��o�͑�_�Na4���f�i#��F�P̟|,(+�,d1�+����)�@����>���AAs(���%xS/ƹmp)�
��Y&Hw�g�9�N:.\ȆZ�;����B ���z���W2r�ԴW�ℚ��E�X��	zb+ɼ��}D�@��A�;�pT�՘��#�aAd��X����t��� �B��_|��b<kK�+fz�Ԝ��������^�J�y�;Iٵc�?�9#C��h�(/'�����k���C���~��0ȟ��e�k�,PzN�AF ��=����r`/a4g�{��X�)l,�"���c}w��F�!H/���>��d3I�@��m�i@T��^�Rs-%�u����.o��_�i?>� I���N���7��㬑�+��Y�.������riYx��~�����̃ьG1�����4��V(8��M���L�����c�W��-�y*�15_�1w�?�e��J��]������JG���K�|�))n�J��C��x���1y��(��B�
r����>r�oڨ��N��C�����(�A�M%���Y���X,dGE���=�r	�*�@\�5����G�����?Z �[�O�2��oE�P���T��J�}��X�L���f������HѯʰXI��qs� �zI��W���`��w��9�u��T�?dC�1HU��i>�j��P�셉��L�2���1~��ظ���g�ЈF%bd�C�%F	zgf�!�WLmЩ���zG���WN8Mo������{�ZV�,U�[���0��9��Q��O���`2x����^�ƽ��
�+ъ�E�#�����.������E�ey�����H��v<z���#)�D���yͣ����u&؄A+���Z��/���$�S{zz��4]EX6��%���2��c�w��&�$.*��Խ�(@�i�l%����T�.2�֣��<3�1QGB �ۇ��v���ܕ�Q�&_9��^]{?�>�+��@K�3m��s.� \��5�1Ro�(�z%�,��s}x�.��m��%bA��|����R���`�C�_<1��y���9�+�>~�C����Hd�+e7�[&e����t,�k0��R�>�6��fʤ.�$�h:��]�O�<�,�{cqs��R���dQ�.��t�ϱ��n�����x�o����	��j!�͸Z�x��
f�E΋-�Xs�0Lr�c\@�ӕkN	���ۅo>��@傞�U�����R�b�a�Ziռ�OEQt k����5��C�<Q������<�+ӊX\?�H�n	|������5�y���i�znW����4�7�Gc3?9���:*b�(
=�^��d��a �U�4nmZ~\"�l�[���GX�x�tW�v`����ꨅ�A0����;8�"�o�-&��xL����+������Z�'�4t�ㄅ���Eh����X���-WkAp�,ə��l�-'�|�1_��k��N�`W������(u�Ze��C�-�pm�b^�k$`�(s$<��G�4Y�po��c���V�j0��'1���9��!kK�MK0�a*z�w�&5̊/��ufm�B��s�.��&����ܠS�ќ��Ӹ���Du�Qл�Y��d���X�'�n�B[F#b��ɷ�����2�g��-VL|��W�Rr�G<͗w_Zeg�������:��-��KQ��C���������v�S�N	YY���_�u��6����;.����L�?���#�6�Qm�nx�m���v��T�B��0��ƴ�}V�!V�:��S�����U&7�K��F�r?�Wތ̺������W�%���>5��4�>�Լ�#@#�����.�'��]g�l��__�MZ���I�G�un)� �;�����~M���-`3P�l�>�y*G�p�a��uq�dU{�r��G�|��RI	M�WA�}���Cve8
�"�X���W���@֖�N�/���*�y~s���LL����A�χ����?�s��^����GĔ/B�U��	��3�G�9+LĪ/)@���]��ު�P]C+U��E����D�;����~�]��so�,��������F3B����_衫T�P��r�$9β������-n���+���h4V�ʵ���b]����~k�&�	D��	�	��7k�A��X����v,��'�eڐz��w��U��k�r$·��x���Ī*�2=D��`�����"��O�ߤ�� O��݄����x���1�[o�Մ3����VϘ}c�$s��Ps�j�
-�H'{J�,����]�߆���=`�i��,2�si9)�=|\�{Cd�R������u@a�� 		�N���ElRU;&�8�$�opć��]ڬ��J�r��ݹ���WE>���?%P�B�����Z� V��~p�}�#zy��-���~��tH"�����[HV��?�` ;$ ᤚa6�x)}�>��/	�Y�v��8���Ǐ��Ч�3,B��Mն3�W��hȂ˚я&�,�C;2�/�J�ge�q���+V|�9!�qTB9�yu��h	7��T�a� ��0� �)8J��)#�?|e}��Z'�R�uwrD�
��'�Q�-��?��ֱ��axc�2_"�sn�϶���JpU���.�=�k%�@�'鹿� ?.W��lI�A�>AAO��5��^�a�� ��,T3'QA#��S,���>׉�Ca&0�H��E�[(icK�|L:��i>"��ۖM�>$N��@K�tK+�<�v	�-L�d�]�̔�Wn�����Q�9��I��Iz�p
�-Nj�	M�hՕVƳ.�4�t�VNY�����8�~N���m��s����M}4���I�AO⣘�F��O����� ��.��j��F4JG��px�v��]�*�W�|%�X��f}%��ށKO9J�Du�R�\Ǚ@��Q�R�Vʱ$N�6�0��e~���~���U�".+Tt;�?���8]�p�����C~9Ï�3��'���T�^���� �2�6r�_�Z& W��֫LTH����ɭWl�±����Ś���e�?؍l�-�>�lo�HLNI7�6���T���>Ż�,�0�߃���A����;	���������A��FȄ�Kų1�C��|>Ҡ"
:s��K�1v\�"�ő?}����4M��(�I���T�����e&�4���:�:T�\�z�ް�՟$������`=��tО��F�9�ZhoT��g~�&�g�~���\��mWͧ,G ��T�S W�U_hO+,���1q�	P�	��� `�(�r�lL[; ��H�ׁ4�\�+؎���E�s4i�(�%�B)?�>10�j������f&s�Ȗ-k�iRk���:'(��y�֭b�v
rn&����^sHE�=�1a=��� B�3���0`;�O���7X��9]eK�Y�ݖ�����Z��*s��X���U��M��"_$�Cs��^7��~��>7�1��*&�c�#rt���~��2d7�QW�8��THD�V2�q;�>Ӕ�4Ԅ���NS	ǇX�LYt8���J9m��>���Q�os��a]�YE�<�[C.����@����XV��O|&Ѫ��P���ޘt�_���uѕ�a�$�����͕#����~�]����ٱ{�>U��:\�"��}%����0)#�TQ�����U�9�����_.�;��0�o䱑>״���j��bU�U�߁%�g:��A�	���е.�����c�� ~s��`�4ν�B�s�ހ"|��nFL�o��y�m4>��vYu�����Iŗ��>i��u�V��g�9����Z��@�5	���-O���kA����*��PuPYް2M�gy.�3��za>+�aS�E��ĻH4��d�B�X��lm|)�RD_�����G����jQf�u�ݲ�UCCF�$��pT�v�+7l<�/'v�.�p���٠=��d��4�3����kC���7bbR�:?K�A͌���3�s���ӫ��+<�`�>��U���7<H0r�����S�;�Y�Ċz,] ��&�������'\�	xύUЋx� K����x4[��]����?�������4�<���ո8�L�c�*;��ݬ^/;P=��ڌXn��������� 4%*&s���`��4�pe&�����(��{�'��"�
�����/�p�J�3G6�z��,�c��wc���T�;	k�9AƖ�i75������ӹ4��eb;')�ŧ��?oZ@b��� I��Ч_�	��*�������f����xC���b6��W��$ƱƅWLY|�䩱x������j7n�Z4y�(4I���C��I�bE!�~p���@�� ���Э��[@�}��V@B�g�2�	���t5́�-f
Q-���G�6|�P�g���	�\MP0�9f^.�ph��r���P0@���{�v�-�t!!HwԧS�T�~�k��� �E\uє�)�E��7���k�dÂx��X5�TJb54p�j�>(���a�
���n�EE�ʕ�P����vb��N�2�#�W���h1c1he�z\��^�:O �}���+T����J�z��K��E��q.�ԩ��{1��숱�������p�J?��  i/��GD$��@�m����%�6���?M���~c�4Ѻ*p5)0�b}�Ji�̾��剮�E�#*����(XWD'#��}G������p���(�� ��|!׊��D��n+���d�s����\��mԬIT�i̢�K���� ��Ě�'�mC��aL�y�_)*0��ѷ����o���KMӴD��9}�
����P��$��i�)[,�u�F|l�=���պ�g�ȫZ��� ���W	{�	r���a���E�X܄8y�q��;߿`��7���#�A��5"�2�>���=�:�#`|I��No3�M7�s�����/45#dȀ`�&S/��j3�^4�G�(�T�n���e+�}'�|�W�뻳���d��j�t��*������m���y}8�Xw�%ȣ��'Gj�J�TX�2�2j5��Ҍ�Ad��8N���H�Dy;�N��-���Ԯ/�VJ��xj��bKvHłL�?g���K]��g����Ö��Js�],MT�?&��5)0�d����c�P��ȥ�R�$�c��#&J|�xԩo�\��3`�����~D6SWF�}��Ո�*H�ƨ ɻ-H��
�Z��"P��(���`�ƶz�pRc�|�T_����U{s����<����vF� |�ն,��ȵ��'�cUn�dt}C�2��i�Pq�Yq9�����$b��?��`��i�j¦p�B,��Mt�	<� ί�!
ރC����+S�y�Is㑀l�Q~�_T%_Nji�⌙�fy]����!������'��W���V�Q��W>�Dwb6���303���kL�T�Uó�vcf)gŘ<fm/�����|���w�ps��Hʋj��Z���abKqv�2t>�+�/�I>�����.e��L��í�ϗ<�#K�H���^N����;H����d�6[��RdV��ۨ�y5|-�@��;
�d�Y�MQ�ԥS��:�U<0��v�w<�����w �g�7�3�ȧ�l��Wc�ѷ ��n|��0S~�}ki��v/�xj38ajM<��Je���Y?A3�'��u�"���f����.K�ݲC�|y�����D�")P����=��Y�$dr��8���_��<{�K�
��W�pJ䩛k�Ԁؿl��pV�|���4�,�W�~�>|	�z�g>�ִ�<�f�h7�\���@��P�d0��J�+6(��j���%R׀6��Uz�BK����k��v�t�u�GIY�s�p�y�!�"���<�*���P��4��/U����cS���@tk��.C�gLљ�7��l͑�B$�H��2���l�1��MZ�=��&�|�@�J@���d_�/���7�������6�)ѽ�7w��m3;�Lt��%���B�y�\��brm���2�,0+�'m�F�ueJ�������s������[!��qj�7����
,a�|۴	S��2d
u�������N�!m9ςsm���Y��"�Q!a���eqa��P���F�,.>����'·J��Q��S�J!��S���E�����,?F�)*�!C	O�IR�:��ᗽI@�������J��k,�QW]�I�N�����4?7�}[�����9���J������'";pEz������tv(�+X�^���O`�|2�Cy�-q�`�D9�))^(�U�C��'!��2�:��<���p���͐}�<x���x�+��^�G���Y��2h"Y�A>�	��8�R|��N��J����[䙦2�ÎI�ۨ(k(AM��a�/�7G�ȕ�/�����S��t��{���ktL[��s��!�������� %o��U��{�C@�"�F���p��M����!k/��H"��	��&�1
��h=	��uҷJ�Ctk{��x�C�J��QaW��B6c��x��E��ȩ�?^�ds޽��O6�������:,rB�}��ϗ3)$�H$A(�{5=g�d�~Ru}���o�p����xι��M!D���N����������W
l�2����S`j��x�0�﫬Q�_^?D���}j=[�#?=����v Bv�j�ǫ��6��6�p#�s��-�Z�#��0q��H��#
�T���rW ��R_�����Jd×�h�
�!�~��#��?Y�߇Ϭkf�����m��+29^���`��״�4������F�:lC'L������ޓLo[�����6�S[����3>���֝�����;����V��_�o�&)ǭ�r��ޫ����YJ0M�_zpʫb��1�ߣ*��GS�`�$����2��U��cq�&�����Z?�,�R��LN7����'n�$s�:ˋ�X{�J7d_���0��Q��P\s���j�X%�9�W�(*�O3�u�_]+T�t��aa+��E���ń2�㯹̭\qG���V(����']�`�J��5��Aë�A�[`R��p����u�!�̪�͗Nk�Ǟ\�ƅ�#��B`,� �ۺ!tC���C�GI���2ʂ�����u�M{�i"���3Y��V�c�yd�R�y�&��M�00��ⷋ�LF�q QZ�LLc����r.�+�^��S���3ؾL}��>��W�0P�Ì<!$�jT#L��İe�9�Ǥ������1i��o=��J�.�@ݮ�:N���W�!�,��eޯ *O�����`H�����va҄�I�T[�4m5���Um��q�:cr�U���#�փT�&��B-��ޝ)O����dア�NU��zp��;�%:��<�K����<��1P��gX�Έ���JN����X�c�����c0.%UÇ�qlk4�є'IXq�T;�=�:oY�F,���㓃v��
Id<vU����`��TH�Cꉕ�JD�* 7f�*�5�f}��'$���JF�U�\��z����������;}��l�	�����j���#�|�F������t�ӳ�����,/ǟvL����La��c{-މ��11R>�$F��Y:�_0�{ظ�n����פF��$�5�t�Q d��?|��-�4��v"�R��ڢ�(z!\��h�u���+w�+@�B{�p������m������Ȅs0
*��L�K�E�Ko/�*��Kod���-�����I�V�W>r���7�X��Qt�\{u[�<uS���l��G�́� ����#��5t�Y&�t���6�un��S��]���J��>4����Q��pد��2�ƾ}EL�M��6���fӤ��Rs`҂PS��>�ؙ�m�(2?F�Iû�/M��tT�K/��{xG�hod�0��ǆ�іEe	��ѱ9uv$_�&��S�wʸ��1r�U�e?8=#��ݳ�p_����J���߬�y{��z���:'f7��f�zޖ@"��=?�����-�2P��g�n���E�^|��%���aô���d�N3���vh�A�/Ξω7˫�[� �$nN��
jV�\8/6�tJ�NU9�J���@�Q�<A{�n�)V��W�������F���6�� �+�m'o�ޤL�l6��B�S����s�e�5Ȗߍ�cA\4�>O1�
������wg�/�=��R3�� @M����
�lj��Ҍt�]���	���Z[5��Y���y��+©\�fgX� ����i,�j~+�I@%���;<( �C="sQ�c�pr����QQ�
;o3yHo���� ��>eI�b}N��ǴJXɄ��Ú� w��}]��9� ;��l��.��l��v�㯷�@�_��Ѓ>B�7�|S�,mL2t}#� �tS���D��K*�o!|�N0r�Q��Rl��:��/h�>�+U�3�44�� K^#�����7��m�y����ETCH�ދ�d���<*��z���������p�I��Z�]�Q�%u�$ûpEJɜ��̶�\	�(���yR��0�n	@#���a5�Ŷy�h�8U$V��2�Q3��H�Fo44�?�6�r1��]�~fF��c���x�~~��1p�������^�f��!�-F6H k��ʻ�E0�o�P%JҘ��O�^E�M��J���ث��dP5:��b\,��S���������إj�#Q��N��
٩�H����"���t>U��V����(u�$��e���z!8E�fH��JW��b�T�8xFN1�	��̦�9BnXo�s���xz��db/xk,�O��:r����`l1��=W&hS�	���-W*��'��7�٥ GsGKN��HRX����u'㨷,�Y_
kHL��S�m�8뤿b%�͘���`]F�!�]J2�,��ĥ	1��W�$U�+�ߟv����n�Z�j;rbXoO�%짴{#r}r�̈́�6�S��YH#�h2'bY�3�24�Pk��j����)�f|5A�C�do�I8��x���>YFB��A�eH%a���iD����fe.���>%}�L��UKV��
M��3��k�[L�G��ٜ�TFb�z���L-�<�����^^K��%����UF�޸�\�Hݐ�3ސص�W�0c<4K-A�&�k�A'��+0�2g���t���c�;�Q������$��1*��	�'Rɾ�ój�����s��ƚ�[����ShL�uZ���~��P6>7�~�;�Ѣu]��Q�`����hԿ��`��˗��X��Z���a�#��f/q��c��~ޙK�ѕ8�!����w_��P(��~�0��m��Q%5~"����=��S'E�M�u핂�n����z���e��ElZ��&)*BF��J$b�T{s�O"���gB�Y���됀��4�ôה����0M�^g��Ι[T߫sS'����+���w:��x�~��`g���K���ea����{�cm�Mp��(5oLH�����9R�_BJ�i�����mdi� [�o+?sN���(.���C5�g�e���	�ѮH}/�Ca��ܿ�����W�Ps�F<��у�p��1��J�n�i�Y��D�i��d�G�3�L�-C�;!��n2�kA��d1��T�0����,�ce���	D@;��;�2����'[��b�����1m��L9��zF$r��/c���&��b�P�����I �^��+Q*S��Sry�;��vB���ĢhfC��I)�����k�n�h�PKs2�9�ql?j7�0����U��E#�F丈�C��oN!��?6���fb�9;ª��n�۰��[�^�iG�Fn�����r��jQ�^���
�����M$[��_����S:^
���fM]R@�.�N��9�3�[�f���ev���L����>��[�*|���=��_6�� ��~У�]P��4�M��׀��Nv�]����&����I��j�1�����a<���� ��ot��
�)`��G��+׍��*划�r�M��&[(�!��yYk8�۶���*|0�)�q˺uHH2�?O4�ɧ4��蔽0���~��ű��a�B���p��Ҩ�E�jT?M��h1ʵ��욾�d��$�ˤK�P��;6 0��0�+��E;#�:P��zg�O�H�?�<jwz1%m�-�ܰ��i����fmǁ�U">�>F/<��V7��o����H^��[U#(�R�կ�ֵ���O�1p)}2��ۇ��sFˤyA9O����A���u����t+����r1[�F"���^@�sV�ή}�!3?r���n��ͻ����/d3�Ŀ��k�u�?��K7c�K-~��v�E�	a�Xg��(Ŝ̲��#��ҩ
ӏ��D� ܝLX�3�n8A`���]g�WWS)t��s���HV��5�"����E��%*���4������a�u�F`�7aH�(��2�c�������Ņ�çus�4<0��Y��a�]��J�K��gh�*%�6�>m�],p�z١�"�x>��f��t�M�U�<�,S���I�G�Do�d�����߭&;#��fh�8��ȋ񹡾�b�~#�i�x;�Bm[��yzS�I,'�Z��[�,��/xXm:���D.3� �}�cv|��;n��h�z���e|��UKg���y��{�ˏ�%X")��$n��V����{:�y���� c����kE�2��E�m�D������:��W`ζ{�n0!_���y,ȏ��;�'Ө���*�k*�\�����|�x��Q\չ�"�6+H�tPnn�e��+M�-$n<a����n.\�O�U%�1��w^����/g_��c����!���o�H^
j6���_��i81-�����;r��@�4���u#��$��m�����M����B�hۗ�~Ɋ��46L�u�|/,@�I�5),�>�/���ߍ�܋����׸$�1�8���j1W�B���Z��IY]q�Y�2|��H'�n�8��|�I ���f�#�(����}��JTD�	�~���=o8)�9r���K�T�`V�˜Z!RȐW����"��� ����D�SӮ -��i����+41�#/x7���\R�S�u����g���l���W��<5(����^a�mF%�l��Z�եӊi S�t��������O+�������<
�ҽ����'AP,�VI}�U����5�\�4�{���݁7w_R��:�	~��xR���
)�Y�`@��P�l�@�Ո `�����񴷣��|�h��rp�]F��� 4v`�K�[�If]�_@6j�߄��tx��u�fQ��5D^.���O�R$[U��Z���!Ķ)�"}O]ȶ����H>�R�$��a�0H��tg�R��@V��\�  :ŋ��mK�[��sS.�n,���rr�'�(�#r��CZ��?����çކ��S��**x��D�d��k�n�kb�/�Ka�mj��X�n/���G���ֿ޲��"��xH��q�&VmϰdVSL`�CY�0J����פ�,�S���>\60RC���.�݄�A`>Ů`��^�@mI��l��g�Ӛ��z�ݹ���W��_�/۝�����C#�f�̲���7\�	qc2�AV5�J��D@�$2;�| T��a��J.��+��0����;';O&��sy ��:�vs� $�RZ۟�X��U<E����p��H�T����]gmF�BO��G�.�X��I���a�W6�n�w��R�T�@�]�8�k�{g�ML,:�dN]����oi��Ǹ^�u��4�P6�i���ս户�T���W��j�^>���D�>�W���V�#��%�ڮ�`��C�t���^��*�ȱU�U��5G�b��y�u�D���=ϊQM��>=)=X�h�wRX�S��G�>�b�]^BQR���ːSj�!�ź�$�P����g�	�_s�լ$���"ʚ��K�E-h�-�X�b��c�)�%��"�t����jȗ�l�� ��� $�X�"�B9Ug��Vm�S�y2�b�;�͈�n6[Ω䠁�˓-�u���Wj�e5�As�'e�N�R��V��l5�^AǱ��ҰF4��-�$d�������a!�.0"ȇ󷄪���pe�WS��W�`|�ltJ�U�+O�v���+����N�ITjo�w����{׏��&�����A�w['�N��m�f	ȝ%DA|��I<
g�&̦��	�kӜ?T����rRB+��FO����"���O�Z�4�$�������I���@�}:�SAAx�9:?�
�_�k��-C��y����`�/�G,��ԡ�ZxGkb��#�AX�	N�臰����}��=�_%�#�Bנ���������X�󃴦ܛ4�Pb�� ϥ�b�&fm9[ 
�����$&��]q�[&��(EpC./-P��5!���+ꈬ�a����9�G��+�Q��6Gc-����i�

��+�
c��vzS�F�:@^��q$L\���������Z��$=�=�Ğc�H�Iv�������jR�=W�kC����K	YkKUCl d�B�W��YβU��J���rK����x�����w�/bg�!�Ǒ�� ��.C&ܶ`)�x�\�`��N��ԡ����,�tK��oHk5Ϙ3�z�-e�� ,�ߪ��|3�͏��sP+�΅����/	�`�MEy���V-%��~F�Htz
�|/��-E�~Fp4p�d�'�c����	��	��,�f�9�	��)Q��9�*Y�3��[�[�zE��A�/SO��ȩI�0�H�L�_�^��PR���k�$�W����Q%�텞JP��B�Q ���MjZn*�Z�~1b�MiE�U9�IeP��(��w��,!ƍ>5�h#���A��<�ƪ*�'�~�����}�cs�NA4��1pC�˛��Bx��zR��z>�4H�s�X�^�">j��pA���~R�D��9�Ϋ�����b��#.J�y�Ku�J(h�S&�?�|O��mn.|* �Ofμ:�7OښP$`1P���|�w1��	�_.�V��.���/�O� �L�U�Cj�=k*:�7>�t�k��~��Y�n<�j�6�f7F��G�E����gh��owH�02��@,S�\ᯏ=���Q��-�6�	��}�o�W��T[g���BI����YF]�M�9�8�g n��������_i>��h5,�޵ೳ�� ��g�eck=g:��!��V:�=u�^����j��C�0�6�l�}:g�;t�:̏�eo�� iB6|^fg��+\��Z� 6B�8h����S|ԭ�o�4@���4����ɾ�A٨�(Th����� ?�����ۈ
�U�� �����4�y�[ߍ Nd⫉�wq�8�V�f!y�;���/)=-yO�J�TLi���{��H��UW��N����C����/&s�l� 6��nl�vfyq&�e� �� d��<�c�K&��*�aG�	Ōq�Z%�2�k��{��GZ�=ۀ����>�j ����A��w§���1�{Z	��eҚ�h�v�p��� i�=s�RQtm�S1����y)bLw�.���Myz-�aj��9��'"6?��L��A��gw��(�W���E�v�t'8�v�8>8|EL80�@z�v廪7N4B�W�2��jQqG�b��T��#��*�q���8p,�%+F_T=R�҂���b����D�qk�f�:X�q�{a	�1�4�d�[=��\�ײ�x��T��E��YCv�K����C$L���Y��nr��P`]Х�ȥzvJB ?%���P�-�+_>OyH� o���T���1W�%4��I��ҍu�D}�=�F@���������55�ά�����-�~��*!f^S;��n_�v��1�'B���ihZS�\�=��_pw��d�d0c���d�0�ҵ��_�������_i�������&����u0�ܸo�_�@��:�q������x��Ą^MF��t�P�yO�L��t�[����g��qV�z�����:�X+�pL�h�T��n��/���w�	ʂ�\�h���G�I�V]�b�`R�j����O!יbf$:"C��aO�
K=�l�0�����$� �V��'{���Xܨ ��|߰K��*�V��Eo��j~3��;p)��=D|���\�K3��"��ظsls/T6M��{�H/rb�8�ɶ�CP ��G 6����{;+]�����*��
2U�ᠥ�,ݑ�cYO2_4��ř[�V�����y��>���TFp�(Kv~�iĦH���eTc�[>�s����;� �0e\����~����ظ����6����W{���������N���[H�~8�I766�Gٚ�:�_�P1)!�{��b�#�� ��l�7�>.����ogMkއxq�K�Z�ո���Ԋ��A�?!�v=�#b#��Ϭ���G��̅��sU��	�� rPoA���W!'��7>|��i���(/����9���o�=��L���1��2�E��j�hH�yd����pd��Ns�ٔE���p�Ԁ�E�����Tr�<�f�J���h�3��3x%>�xn�h�>�w�6N	"W��2X�C�rl�ARвp��$�k�a��<w���ڈz�44@PK3���$g��U��ڎL!S���q�O01G�B�Dc^x�C�g���	[��%��]���=,�/�2aZo(;���針$diI�=���S�G��r���eH[���p��k_�1�]�0� `kxc_��n�iȫ�&T�^(��P�s�1{x{��HN� g��-!v�X�Z^�>�p_,�ϛ��.a,(K��8KU��(\��6��+0?�=��L�^?'�~�@��g��P����'ǻ���	.;~���6�^4���|���mCe��j#���ޏI����%���S8w���[��c�t�͛�#!�0���d��(��K7D��{�rάl<M�4��{Zɿ���@% F�F�6-.?k�0��p��ٚ�8�²"=@5��7��}���p��Y�4���[=~�@_o ��	؁�q�Ux�z�c]<�A�����;���ض7��~q4s��l,(߲� W=�R�d'Z��=)�cTf]�O��lÕpz;�n~�n?����8˳������o�D�):e
���ײWcN(��d�_,%�ip���b��8����z�*|�LP��%�&m}�q���0���I��')��Ft�Fm.Q��)�3�TH{�D��Cl�:��1�*�g�Y��ؙB[8��-��yL���ϔ��������UB�v�M�o���UN�ÔT6�?�*�r3���)cl��uĸZp)��@ڮo�t���q*��8u�	�� �?h����������%: m���D��fZ"a�l��RQo�PxO�׭�Y1�@t���ϯJ���np�s(��'�Q�s�!���㷙T�w��{l؟��,.96L���Uv��XC��3#3��L(Z��5��iD�>6��ʢ�^Y ��a�PH��v�d�By��]��d�^���S�;�qw��$��>��hJe���u'�䡨�#{r_��<��|g�CQ^3hN�]U^���{�Im�PZ�|������mc�F��l�ޢ�0T�ǈms���@�kK�a[��$�˳�6�>����n��T�#F&�̢ĠH��θ�WѲ$�h�4V��\~���&�_C`q��Х���0���{e��������0����u,���{7�C-t�g�,k���-�%�v��Dd4Ni����&c��Ob.+\�uv�,�8�/�K�^���"]'��p�k�r������G�5�V���i����O}Vxd���൪n���N�[�o� ��� ���-��4�7�V?���h�?��4��orh���lf��L�g(J8tGm����c��IE�'������C�UϷ�^��i���N���LC�ݖ"fS��EG��"�hi�}{E�[�$�2-z[7p �����<��Q,������hB�AQ�B���3�~��}ʸ3o���qxt�$�FM�xM���+G�)�jV%��Ϗ>�4}\����Zw�Q�+UU�ři���@���K��"-ޭ����M�n�:^mz�*�ؾ�bɷ�#x�^�h{4�����B�}/���Jx5�	��������1<F�u*��".B�f���U�F�!�r���}��v>�'}��5:,3��]��$��Лt�M�g��VDb0A��N���5��C��0�L�������H�oBD	zG��;GjG=��t�E���d����o�1�r�:xܧ�!=E��;@��C�-�SV%䕳/;��@\�����SE���jѴ(����Go���޵�P���#Rʎ����QJ9M̶ ��d�ӵ��4)����5����yH����.�ia�t\y�m
�ū���Q~�lDA���!bi:��y;�+t������-�FXZ��aa@�6I��s���E?�/V*�f>g+���X�#�Û(��li�}�$'	V�\���x^]
Έg��gw1��5�Xx�7�<L�Z��@����<�M���c��b�{���m11�g�a�#í�e�Б�$\���7�l;4Ew�U�_��b��¼0�ge���=Q^˃چ=)���[��c��8�,/ќ�,E��x�h�V��39�9i�k��^lr_�f���_w��nɯ�w4*M.���C�iUg�*XA�n��/�z����ǰy�����j����T����rs�zm�5�i3<�Ū�}Z���w)n��-��s�b+�E��?�K&f�7��!��q�
]��D�VE��+|��nj��kC�O<w������Cq#����
���M���y�"�%�K�c� �8�=}�YK(/{;�֠;��0�]�^��Y�һ`w?����zP�%�I�❲/��O�)�=����Po�e�p/���Ғ���r��x������Ȓ�����11�}WB�'� �sYH؁v���
�vp��!��[��B��0��)G@E��~��:ch�K��J`�i�F`� 2E�17e�����#���(M�H�%�؃��0{!o��~G}����x;���a������/Jr���,?�#F�א|�0�w�9m�C�K(�`zz�ɈhTPc�W۪�=Z)�l��R�J@ـ*�{%�x�� �-D�:��Joc?�7�m��_"��.��oٗ5���ﱉ�|q�.١냄�Vߖ�<[ք�/G)\ٟ��;�wM� Y�o�/��/xҘ��9�b��|�#V0ˈܸ'7�z�7*��2X,A�$>#D�A�{�|Z�1�@���Y_�*|_R��}�����m�7���CJr�4�X,N@���S�l Ӡg���G�2~�����=@9�4��Te,V��Pa�l�����<��;$$[�&ՉԨ�jm��&��Q&��U}	�\��2���T����p+y^�h��kM�#��ۜ�4PDB�x�i��6#���E�V>�o�A�I�p���j,l���{퇳���Z�lxH�7*��yc�xu�H�P��&Y��[IZ�%�vX���l�
3zU�X!���Lw�[�xB�dغ��rA%� �>�Aޜ4��]���`&q,�50B2[�/$��B��_N�̑���*�J��!᝷v�O�k���{~���NʹB̃|�S��7���g�9Y���� �x2�=�l������b.�X�� �A�K��{�2w�8$���$�v`����յv��}&.Ou�v��$��� �=.����d�P�]K��V���T�M�Ӛ_���\�����#���`�����x3��
꽇��������\��to�k�s81&�K�kL�	<>�)���������y�mez�2�T_E��s��~�V|E�(�����tIuo�],4�o{�%�w�U���t�𞻅.�%\S�.��:��ŉR���j�D�Q���c����ۅM�SDMj��=����s:�РL
��3;mX1���yc�i{��-S3VD�{�uL�*<��	]vEC�C7b�[����:�m"����q���Yge�:Qqd��qM��m�uv��x�E��No���d �g��9�Ŕ���9Ǝ�^G�Zd?}�X�x��h��c��@>g|m�+�c܊��ry�p��J�P.���w�OM���UZ��+r��	�%kG�RoԒ��ʬ�.�-4I�G� �p�S�hҝ� �~�h��M��,
� !A����,f�FY1��"0��n:���"�x|�&���um&)�mɲ�3ڴ'I,(�<߭�vV�r"��ۧ[F��hm�=欫6*5v�ί��oZHȬg��>��z{}�[d�ː\$i��BC�tȿ�o����u��|��;��?Ǚ=̓4��.�E���D����@� A��_�a,���ִNN����m\<4^S�9��N��V�����vU�kZX���m/lLB����BKI��Lۃɪ��Ѓ�(�Y[탐��@�X<������H+��m� ��c��wu�>�`]��H<�
p�o{��'����S!�Ԋ�W����HV��#d������7E��]&x�\2����G/���L{/qj��(�4ޜU(���#>�<h�L�[ᘤ�� 9�[O�t\w��On`�u̻n�c �����_��W��\�9�o�}~�|*ϳ�ݔ����N��*�11�=jIG�ŭ)i��W��P�x������"����e ��Z��C��@T�Y�K����WCQ1@S�� .��'�]7<�n���B���W�v}��lF��ƙ���/����4�u�L�tc2	����_�t�{O��N"&­�t9G��8�^*��#n�I,�t@�D�w�.�$��M|��������y:�%��xnM.�:?)�.3b���u�v\x�f��8������ш���H��?��
�_՚����}>��Z�'<�UJ�8�b܂��3�����X;H'ƷZ�� �J����`�6M{��ó�"�	<%�b��T�ν���]�y���g��1"W���Թa�Z��\�η!]X���7�oi9`U��M4zq�Q����x�HY�I��ɍ3�r���]���E6��I���t�?�W�:Kk�����)5\��i)����Q�|�p!�H�����8�*���fI�m+
f}h_;`ѐ���^�I�SI�k��݀��t�ڒw�k���C~l)M����]r�^�.�B�{���*=��O�ꅲ߯��~W<G���~f��f���3^��char��bϏ�:���9?9Ĥ��绾�ۉ������f6U��V]�����Sk;U��v|(�I�?�Ur�*ŜR�a��O$��j�#B'P�a.�Q8�0�5�b�Ws݉Ñ�#c}9�1uи�q�o�o��d�iR���5M��A H�nn�s�xgK��=�I?�̦a��8Z�-#��(I!�'a�C?	&[�?����(.����#V�E�R�G�*n�JvP��4�3b�6���>���Jx�U4#��dP�4��q���WmO5�41�R�B���%!!���$��nQ4�W���m`NgT�)��3�3 �gK����LbYy-��/��ީ���mr�Ӻ���P��߷bH���^BYңҒ�TW� π�D ˅�vt��?N{�Z�K����$}S�J�|K�y�jS��1~�C߱y@��u<�(����>�%%�]4N��1��;!
q���G��j|�����KƑ6���b]�3�o���æ���M��63��HЎ������I�WϾ��3c,�*{�#�n�a��`��_�c��3�F��>mxH�pE�]0���� |f�Dy�#�4Ijn��0��WO�Iri�%�?#'���4k�m�9����F�f�����!��J��/]^�������B�#.]PX}&�e˒5uTwA����h�qv�}�#����"�,�N-"J�� �@�9�N�����#�:G���~F9������D*k��1���{�Ә)�w�Jm�b
��QD�P ��6F���.�G���%�Z��� ��q��Z�ȑ��j��ͭ4R�<NA�X����՜�ih��� ���Gp�0�=�C
���eQdDR˅Q����*'�/c]݈���1�"�!���:E/Y��v���~�����a��\%+�ȍn�î4�l�B�q,=jX�=��)&��8e�2��U=�O��@�V1B"��30�^�(�`�6��q�.Z�8��Z#ח�-����ߒ�L)��a�mS�n�X��؏��i1@G�g�y,E5��j��A(�ݓw�Ѷ��C�R���T�I]l������3�4�9��h�� ���=oE:.pv�t�#�z-���+N��]� �@%�����=Ȫ�y��/���Ou�A*�}�>���[�8�v��L��۲��_C�sj*�@1C�/e����]������Qj���1�B��CA��J&�Ht�P�X�z�A��$r�v�)PM
S_���&:4�_�h�>�����8��9��I
z��*���נ���|/����<��9��) (����j�FU<Yj2��Ǿb8K���{ܱ��%��D߆r�h��yvJ%ӣ�)qQ]��y��r�Md��J����s���f����_i�7�{�V�e�vkXH�FQ�"�,�[���ai:}���Cj*ߋ�	�*�6���/J}vO�Wl�C��I�f��|���mX��W�䔹r4�DA�!�B<��t�l�5����\�U�+Ӈ���S��8�ry�����z�_1�L�.�L������֏6�"��)�jl"[�b��>
�xH�~G,Gۑ�cN�b��s+Q0���]v��BE�%Z�gi�bw���E�F����>5
vӣI$�Q���|�a]�>cH��VPr�|:yQ˼Aԯ��$d[#�N�������}�,�:8�pf�a:,�ɾ̋���vHm��2�!��"#�.
mY�·���PR��yY�WA��4?ޏ]��x��""%�g�W��d� .�%��N$VU/L���`�rz[�yR���+.\�tP�S��$�8�l��j�������������#��L~�5	�>��g��ZMOR�N���s�*l$Q���H�H-[M6�L1׈}��U�.���4�}�C�?��]�H�ټ2�E�%��._�X*;U���>`He��yW��,����נJ��+j|��g�_�z$E�?�<X��©A�E~!.���"����i��j7EIn���b�nԚb������3cP��
S!/�yb'��k�ɥ�ޏ�w�P<2��^p�<�#�)�i8sk"�ߧ�3O y|��UD�+u쟡s�B4mE����Z���b�e��>�z�r�@�=w��5��F����A@��ڹ�'��+��vN&���
R�B,oW���i�0���W*q�/.>]du��֓�1;A`����,��Л�1=7�S��T�����}0��啽��t2�«��GͿb؛;#G<0��C���o+�zj�mR\��6@=��M��3���������M��,�+�h�ռ�ƪv�f	0���5�~�u����\�PZ�tD�A���Anx��)Y�gM��C�FZ�Cz�^��*Wk�9͎T-yK��^|0R3bf��@tu�'i(n�R�<e�S��G�Ӡ��]�) �ct��P�y��O�?���aL4�>]X~��VU��e���Q3�1��-�������zC����՟:�/���7R[<h�R�����׹P�a~�s��0�;�f,O"�F�1Np���o� T�αd�}�a��*����@q�%'�Wa��a��� �� ,e�Z=h����^�=|�.�x�#K�!�^��g��R�v��.�K�N��_�����j��h~O�G���-�+|��@w��D7;S�H�*��dJ϶�L��	�T���e�'G=%7���v����5�w�Q:��p�1_�V[�ʕ "�̏�@E���B�Pc�G�'�Ա�?��E�ҩ�OW\�}d�bB�s�����L�c5a����]$8�]����v��,�Z�ǢK!�\�TBX���m�������j�I�A�|�Q�C�.��!�[9���)��Z�nZ}�l��h�,�+�b���v����=� ��|�� �2��W>:��DY5�؅�p%�qffҝp�W�9uPz��oE�ق.�����b%�oZ5�Y����"���� �҉[���ϿI锅��b�s4��ic3���b��_�Ƀ����IKɋ�+29�Ȩ�Fy|�x��#�v��ӄӋj"x(p��P��B{�Q�Ln`���Q4=�Иi��sd��ݞ_���1�)�S4��U�'d����w����(qM���Φ��l�����{���*țr1TO�H��.�۝�
��0ސ˰�z�T�Ф�L�7����v(�}�R�b�6u	n��P	[�����a(V3TB�Cos6��M˪��7e�iS;&��\�i܌ho����l��}T?՝;㽽ƶ���t�I`�_�,=�L_�!"��=�z&�x.�>ڔ�Ԗ2�̓�r�R(˘��p�xAS0�r��R�D�R�	/��ؐ��]��c]$�-_m�ܶ�f��|ub{ք�$+#��7��L�̷�%%�懁 �z*�Z����2�M<�ɿQ�j���?,?��g�h�x��i����i�G�������F����q����D��Y��Yq�Q�i�.ɍ����,^y� ��� ��o��"K���Z�7b�]��4~����+rI�K�<u�Op72��iA����tWQD�b��%{SP*N�H���Y�Y��Mc��K��ຕM^b����볬?w���u��͑�Ta߹�Y�+r�M�O^�B�����[U5�T���+gܟ�im 8�^ve����欎�x�a.I�F�	0V��~�~b����R����n��(=��P��Mߦ�[��C�%S��f�O9����w~���_�%_Eu��5Hnm�6h���� A�k�d�FF�^|��x�F:`	���:Ѷxg�p��-ci r=8ɟ�	�����T�r��y-�w��%1 �W�O�HHu��&�%��5�P�O�W��;��hr�b��v��2w��6?l��hM�o�>>�Ĵ�ft(�?J�47��+�lZ�q�>(��@
)����#"�Js���(�5�V�ɳAa�N��f��;l͙2l~������|C��
Q�S�`N��Dr��hD���}_hRHo9��il�T�翺�F�R0�2g�����,�hV�)�㹫��0.{�hw�	%���/�b<x�s�B�Pp����� Y�&�٫��8n�UU�>n�t�^��Q4#�����r�|��������Ռ�=���jϨ�N5I��u�j�Ox?�1�X��h�66ٮ4���~�`r{ZA����T>���ڰ�QT�F�[�� ����j��R���c�	�1��ܧ�S��d�1w�E}AbM�zk�YY0z�ŗ��~,�,_�(lؐ��Ð_����笑��%9~�x[L_�'���F�J�3��l쁘�0�ng42D���"�������ΛzR'�~��~����6�e�''N��Z��%R��&v����2�`��9�;�Xb�]�LY���8�gD~��&�f�w絮��f�"I��� t���}��
�3��A�g̳a�3m����W�{��q��ͪ%/
�\Ɔ���� �r���3�\T/P�Pz.���-4�G�}#�}�<���)�^�v�1��:Ԡ?ʋqh�on9�ZM@�W��pQ�^�5� &��_Cƫ��z8ے��L��#��T���_��$!��#��2�"N��b�6�(l���s#��vz�D��ғ�B�f���Ǯ�K�m�H=����9��+�������������Y�%�P�dl��!��38a���Wǲ]��j=u؜�!39W� 5?�뙇2_6������ˑ�`����am叝�[�2����ly܀e�l������5�V����� VK;�l@�SJ�R�_:D��Y��O�i890e�S��u��Zq��v��،}{$���uɩ��F��|`E�����m�n6����F��� vUY��7m�u�G)Y@2Gi�5�q���#�.ݐ�����Y��TD��#`��t*�[F�K�4O��O��|ל>a�� 6	��ZW�-�	GS=@`N�����Ě�xBPdhZ���Վ���c��=���ɓ>�}LS}1S��(l@A�%��'�a�����f�-O^��q��r@��e}a������l�Ai�,{�	��t_�L����p�)*z��tB04s���)��	�%�k��?	�ºBD���t�q����G��hV�ٛhv�u�':\�$��Ԇ���NC[G�&k��lU�n.kJr,�	����һ)�X�"�3�u�raö��7B{=�J4���d%���H�И
S�i"�����
��P�o 5��e�o?��T!T�^��h���#�=�̑��ocJ��l�kA�O���-���,l7I�� �0U6�
e����>�|�5�X~�,�j&���/OC�#;=_)�䷉X�����ɖ9�@�����&�=�OG�nv4�Un�"�`��LZ�[r*���)dO�� /�9�=8�u�qLJ�q`�W�yu���O:BL�{F��9i�7�٦�g+e�(�m��k��'��4���T�*w�}A.�X$l_�/>��z�t�Y�W_<a�3�Ń9�����Y�� �Q�����Z-LH\�&�1����4�R��=��1=��ѡ�
����x�U��.-�\����{�dE�����B�������ǿe-n�l��9��j��#!�H���fM�������`���g>��7�����Kt2��o1���O���s.��a�Eç�H���u��(�tA*AY<]��#M�O�#��vMAk�uJ0�9�9�(��n�n)�`��j�s�� ]����o��]����UT4/�����=��bo�?-(���%2]�M��{>�y��SV���o�q�d"��#Y1(����u�&�4�]�����r7x�_${�6F}ƶ$B��·�����z����_}9���4����r�b�/�m��gf|BDy�"��G�q�L��%}E���򦫪���q�$Ԛ%È�Z�Yt���c~A�ۡ_�x���<K%�!<f�+�ph��"<G��c�����^�zC�
��>q㼽�=�uf�=W�s�]�]6G}�~ٺ��t}������� �X((�e_Dfk�m"�R�ha��E)D�*�~T培6;st:$K�rql��CQJ�Iɲ�ٝ�őr����I�1�y̽X0�ǘud����Q`�=v�o2�Q��nU	���%��%���:��J��.������ܧZ
ܳ����2}z-`��.ښ��Rz���X��Z�EGI����6�4J�kȆɤ�_���D�?�!`~Zk,4.��[��>�Þ�^h�7,��ܻ?��6��)���U���
1e�|�%��XkFFI���'	��^�(��x2%���l%�:�޲�h���_�t��'��E�R� �؋���ך@�|�]��pk�Y�7��}�P�,�Tc	�[|6ƯT�˰"�4^[A�A 6ɦ��þR�D���]�LT��������T����FfD�9�\�K�?�qS�(J�|��0O��+TW��v-�K�SbC�'f�;K0l�u�Xu�G2y�k��!�c��(K��f�;Ady�=; �e�7��$'4ݭ� .p��Ct���J�u��G?���wO[f@B���f�#3|Jr����^?�*�z9ѳ�GR��H����.���SB;$4�+0�k�w�������}A�<�f�5o�/T��rʽD�}�X}9#�+�M�>����& ~�k��������J�4s�bQnHv�;C�f�iۅ��8=��?�{4��6�m��L�����s@�;��V&��hC�r���}N��ǩ��Mc};�V�0;-��P�X���e���\���- �u+�������T�Y[��;��I9|?��1�;������ ��=&�qP��@�g.a�z�mg&Jʩ4^�|K� �3�O��2��,gJ��!N���4cF���<P-�6ͳh�r{��3o
`[�骎�%�+�5k�n���Y4��~d�jx��b7�qy�p��kzt�~��2�o�����Si��ҽ�a�z��\� %�f ���z���g
�C:���{f�b�JOҋ ֑��x����uWg7���q�#<9"Ρ���B�꛷|,��Wo0�C�P1��A�����)!>[&Ɩ��^m�ƀ�AC�[~�u.�q�2�#�	0F=^��]Y���#>�&F,���'��'���:����~��C��.�LXÍ�l�i/?s�*�	����S ��J���0K�t}��2���D�p۫}J�5�Tט�Z\�j&!B6�H�ϋ��W�jp����_s��N$݄��΂�R�!u�X�U��(�18�t�5�y_~�4��aAG�|�F|Zu��]��^����=���	�L�k�T\�<��9BNT�G]�SG���Z'�UA�q��T���е��-5uW6^�	�s���w~����G4EL%����+ ϕ$,e/�Z�>��t���m903䑢��(�nAC^�-LЉ+��'r���� �
�U��b�;�ny^�t���6��~մ7�����&��Jx�����?��y+�4g�j��r�F�L:�+r��ǽt@S�_�@�}���g�zN�H �84�!4:����~����k����I ~�RA�x
eƧW7h�R��IV }zJt�[��E>�7uo�ePD8�s�|O����'��v}���˖�ʻ<�^J��݀)G۝ �>;���|U� )'VMF�w�I�(/�?q��!��Y�NB����)�,a%dw�aco#�ʊI��OVns7Q5ó����v(x�u��<7 �W����a��|�܌4��� �(����lѷo$�/���ʃv��"��ɀ���fx&�ڳ}�{/3:�uB��ɒ��`�"��,�T���>X���i3�����E,��#���v��m�jL! |
�Iw^������Mk ��L��3���C9yGE���*�S-)J��L�Sa��?�*�5ɟ��aB�X�������!\jξ�| ,�؝\�@���z�����Nsݻ�W�6���Mr�6˧��g��=
4Rͥ58�����fA,�@����>�2>��"ԫsVm�=o>o��,�^vVQ@����9xo��@�>l�U42|K�E�=QQ^���m'v�Z�	�	r=N�i��h�W�Y�n�޿�m��NJ#���i��e�s%���!����Sje��tb<Ej���	��2��@���*Y#�9~v>$�1�|�o6E�!�=�f��DQ����9C�Cq�`���� ړ��P��1+T�3���$ͅ��v�E�ł+��O������͏ѥ�e1�������>))�YO�� jq�p�ӱ-k��%�]�ͩ��)��!x\h�܎�N6��|�Bߣ;<%:�炽K
�rǃ#ֵ��(�6��1Qg�"a~%+|5�گ���Ü;���#����řnp�tgE�F0[S��6*�@*�6<}�9�a͒��8�͉�'����fw	���;?��#�d'�V�O"�c�'o"�B�i�*JO�C�[�/��n�-�R_����%��?�ß��ț�Ƅ�z�die��%�{`�ӨL=}���c��@�9"����ӷ��#�y��{���Y;��T3� ��g����%�Ò��5��{���a� ����`�T���E# )�=�$� ����&
��@�~}�H��[�!�-oW�5��bV�*�!z8'���'�[��e'68�2�����|����	y�p8c�'�n� sC0/Fx�����B�i�VN�9��]"�,B�a� [��I7�ʀ��9����V=@�[Bw�L�;T������l,^)5ј��ۄ`nb2��d�is8�x��tX��yF��)c��1Z�t��̳����T�~�v���V�C��J+g�do���PX����e���e��V��_���A������_��8�<��F|Eۣ<Ͼq敉6U"[�MP� �N����*��K׀Wwg��p���1�"���㲫,N�O�S�����:{,B8�x0M�R	��n%Z��C�E&��G��7����j��[���B-�wS��5�M>��S
�������+J��7ܨ�Cqu��1�
�Y�l&�C���+;����;c6��g�I ���Q�%Y��,��ALUV�R�	e��G�Ɠ*�۲/����;%$�w�F�!����u��� �N�=�R��g��pg�0$)��6+D�f|E�jhMZ�;J����a�s�W��!�Z�e�Ǿ��!Yb,�08M�\��͘D�L�4�~��@�ڟk�W�|lp��U��e2�Ӗ��P�W���k�_�M8��.���Y�4փ�����@�xQs�!fG0���>ގ���}�{O	i)�w�es1��?��X�6��=��3�\�9�ӵ0�����&FN71�o�t�v������8� ]7V+'�a�`���^31[�pĈ���ٖ]��o�|� �f�e�Z���~��;�N�?�Զ��BE�X�]L�H1�cR,)�8r��-�]���Vs��~�~�%���	Al��O�ߗ����>.l���9���
����qVCB�X�<�9�Q��)7%���&2���KP����:�R0�XA�����XKWR7��(�u��K�b��������|{��u)t��p
�3G<�/��iY]uGq�%$���vRs��s�5��$7[���$C���6�����: �H��̈dC��z��������[fc|�{���<0<Y'��+��#�(KJ�㐵.QaI��ԹH��9�ʫ�`�f���c5]�����Ɏh.�n������~e���8|����Ɓ/�S�
��'�V2��M
��x׈�"�`=��ñ�4"̚��{R��D�H�N�.��&�v�/@|�~ѿ��_��I�\�h�1L�9����6E>�����C�!{���R�����h ��V㱥ɪɱA��9�_��%{:LMy�ޢ�Azь#��Q��5�]9X��D���d>l����Q�4�_~A������QEx�{\�=
��z���L��p{��������P�~Cٕ/HZ�1݋��1��*g�N�r�d���*P�"�خ���˄\���kڒ�*Wk�/�����`/GgI6��%�xI�K�O�D!e�`8�:�e3�A���m������7�f�x�O}2�m�G� .��� y���CK�a3�$Y�__G�}��C�en��i�wX@�����-�F#,}���o�Ɉcq���ݣ$h�vi�ur�^OƩ�	�J��`܎�&�r���eBv�����BC�:�u�j��GXcC`A�q�?�p9u�����8z\��K�H� Ʈsr���b�kL'��3�F"��!$)�s�������
R/9�Ϭ7�p�ol-�i�l��3d�{�9�5븋�nE�"~U��Ǫj_��2�����E���! !�|3��ưyl�b�%�k݋C�C�p'O�:t�%�I�����s���ԣ�6����*���7Xα�*z@I��E���1 �6R)	 lPf^��A��P*'���6���׳yh�1�w��cԍY�!z�U̘:��М٭@j�V�n5�xЦ��{�H�����>��e�F�L��6�Jƭ:�\�X
CZ����Rmo����O'\!���sE�X玾��Z��Ke��w}e�z,��3ʲ�
����	p��P��ox�)��%����xE������s����q�z�� �;�箬W��ɻ{7� 2����iK�Y��u2ڃ#x�N�_}��*��Gؤ���~P��g�9	��VƂ3%���$�6��������G�f�֮��\ i�\Q���QD��*p�>�昤:7��
º`�eaNc%W���`�I�F�[��1�������D�ϩwg(����I�a
��l�H_�?Nf�D
�Wq�XSR�b�?Ze�M��t�G*�\����m�#�M�g�i�>6��\�|w�+�ok���-�8<������6Q���P'h�Z8" ����=�UXJ�:Ԙ �>l}4�V�/�q�LA^�#/rĖ�O�|��D��\��4�4�	u�8��n2n��M�S����ʧ=���N�9@va��X����)���6m���L&>��~ �w�*�\�b/�k΋���RB���`�n��YCrabw��ZPl�7=|CfRq��ǅ?�5�N��.fx�~�kd1�L�کtn�ݮ�vĖ�O�?�}�����K�ep���EE�n�u%�[��P���'�ϘQ�	�r�́g1���(��v7M KP�ή��e�m�����9�&����૊VXs�Ļփ��v�>W�+h��v�=ͯQL�OϺ�9�A�ψ}ٖ�Kj�J�]i%"�=‟����Ǎ�ڞ�؁0�g����H����	�(��͑��
��m��2���'+dHg�`�[��L�9)��brO-M*��	s}��@9�z6"=�􃬅���L�1�ԈO\X]V����P�.�[���Tፔ�;�n�qsm;ʑ:5B)�j>�(Ɔ�p�V�5��:�R��!�b��dُ��AЛ�מ
�0U�>L���T��U����7�Wbq:Q�O@1�H�
Uhm
��;r���aaI�{J�8[ՑYI�>L i7��.�V���3Z�����]������<l�Z�����6%HZ�(�!��6���5�<0�b����0u��߫�Ǝ�}��e%"����A75��)jnC��̃��T���ɑ)�̾'tH�� �r'N��Ėl�<ٰh�#J�Ћ\h�P��!�˰�U���[z����c&�rX����p��Ұ(3<m��f�Ҙx$�:\�5O�i�=\	��y-��^��%-�2%q�I��3���y�ы��x|���$��X�|���	d/W����yv6H�:-�2gƽ���L�FB��ē%��	�˄J};����A�KR?ik�D�v�^��m6hju���^��}�FeH��~0�4���nhM>���'�h�w��
H��N��J$�1�2CDq��l���Cp���^��eWz��^d6y��U��&Pذ���Ъa�X�����j��F/��O���c��B8�A\�y�Yb�M�#�n�Wk�w1�'"|�$��*a�23'�y�{E����1o����&Y������U=�r�=wWI��Iiw�k	��
��i��N�:,�@]��"B�\#7wa��APz�mޯ�c����k3Q�&�X��&��  �Z.4I�|x���t�_o�}�t�u�ە�ٮ����Ɣ7���N}չ71cd��V���x��>&�<ќ��N2�.��E@��9mT�diM�P���ʳ"�m��I�H#V�<��c�<}@Ț��={��N�X��D�	����q�m��Cu�b�!{թ��O�עQ8ܚ�e>1�C}�A�+M��a�Ewy2��%��X ���Z�-hd�\�Ɉqg���;i$y%�!����>�_����g��B_������p�^((���k0�!�{�Kц��v�$\�|�����9vE)7Um�Iʙ�,�����D���S�&�+��-��^���3�V���n�� ��V���(7�e<JG��İ���h����TU4��z
�k=�j�/������a�<�#�|	��/�|�w�C�"a���61#��Z���-��c[p������>�RzuCR�B�0���O����p�O���ޛ~���c���K�'X`����n����I�x��*d�P���g�_�W;�#��tAac5x)V�l�`�d�Q�g�	����^�~�KH3/�q��W?��;G��ͺۿ���ᄷ�Nh��cLĚf��Q�}n�>�hu(Yε��H�T"�or�DI[t�|^���`y��"���J�aY�L7M�Y/�r��U��DGi�,(�����@�J�����L��DT�֐Q��cAdz����S?�y��24k�;�z3~�ر�1<�F8�N����SU�V��Αul{'�{	j2�{)ǩ�F�f�z�Z`�+ȃ�^M�O<�RޠdY?���qm��j���5�۲mA7�+6�2u+���Fl��b�]�)��3@f��af�AW?�E�Xt��"�ԏ;U��K��{<�R������o���ꢐn�wpY:x���11V1� �O�U���礴�� �ZKeR��)��ҽlG �Mz�/�tN�������3ڷ�
WU����Aq�ۓ�>����@8��4h�e(���N�����+����'o�'� (.�}��8��%����_� =0>��0�V���MdD�#�ZF-f3��c�P�NsB���o�<Z��g�N �njt�1��w[A��o"g��L�5��;���1�4�������F��֖�LN(�5�j
|�[�q�P�١���;߆�uƅ�Y�<��֖��Q����;��rk�o�"���n�OQT5��8l�`ژ8c��e��%0c��	+Iݢ>��c��R���$N�n*'j��VT;���h�b)�e�2�f� Yt�#+����|�N��"�iu9^��,g���VT�Zb�fW�	�����ݨ�|�վs�r�d��BCy�\�W�b��ǄX�;F29M%���%MBΥ�p��,8��99C���J�3�����S����7���NIu�zbX��d]*p��C�lz��q���61��@ɜ{ ��Y��Sg�|���ӆ�ź�*$�s��i����2 T]/�b�s�pY����;�����l2��+%d���?��ŕW�'Uؖ�hdA�b��\c�u�;4U���6���=��6�D��7l�Qin��r{�����<����_��@�����;�^���y�{[G�v-���v����ز��bK�s��}�oȳf��/ޚ�e����;M���N�}�jNR�����^ق������S�?��*m<�+�8f>����\j^��k����V���`���� ޣ�r^}x���L�1ɗ|b�3� ޽�^ 5��N���kTkjQ*5����,fCC\y�oM��_����X�Q&����n^��+!���Չ%D_i>��=	l�Ui�<��:(_�KwU�ߐ2t:v}���	�G.P���6QT�����I��䣾4�/���u�.���Ju*I
��%�=
�Í���,���<v�Yl
hV�����n6�L8�ˋS�vQ,���l�!!Tz�	{�;��$-DUs�����S�0m����Q��e���j��%�L8Vno�7T�j����崣�l�9���s����3�z�G���2h����f=�`Ϟ�q�K�Υ���2���dd$�/�s�I捹E�ؠiK� vŉv��^_B��!'��f6��ʍ>}��a'ܕѥNEդq�?هzi4@t�Ռӝ�z߄/o�Pb��"C܀�$Butl��r@��[9���j�!,���$�3����jƎ~qLd��^��Y5�mH@hQ,�[�A�h-j�8 2��B�//���Ew��y;Y�q�����ԯ"��w�q��XWq�g�^Z��,��$~��8��˩��!ç�2�~Aa���3!�m$�/�f�NL�d�R_�����{�)����q,��T@�Hl��RL�C�K[Y�'_I���d"@P�4ʣ|�l��f�uyA�C��	\l1q�]Cuh�Ue�"{�E�����;g��ڎ��-��䙰�Vmb��$��Dx��@i/�B�.?q�e�z�=l7�2�m� v�<Fk�:���>������Ӕ��	�1G��7��.S-S����o��1s֝J_�Xo����	3�UI}��@4���P���*P�p�G<R�߅�Z��MPy��e[�H�W�QU�b����\�������D��P��SMU1~O���e�٢{�H^����;�,���{�OD��_�m�%�4[��aH	i�����4�By]7�]$s�'����	���۳~Q'E��rQ�uϨp$q�����9�p����E����N�a��5iϥG[lC]L���j1ՄU��X�8H1k�T���3�Q/��p�X:Ji����=N��[���ǀ��J�e1Y����aJY�{IM��Yڧh3r�7���i���F7�+�`P�������ý���y���xπi9!�?7�n%�;��5�\K�wo���Q����_A��uZ���ܸ�f7����L&*��)�"jl)������$z�Cȇ������ M��/3��J�7�e H�`pM]l��8�Je������_~����s��k�ۥ�@��/��A�yz�l�A%�/�I#��$aU�/М�#%{�#�֔�ELR��-jF��0%
G��uGđ��3��Ά�-,c�}��UG �9�����(�c|���kg���K����Oc� o��Jm�Z���)���SHZ�H������s���G�/�M��j��S��p`�&ȸ�?һ���	�ΊFY��W��&�~�S��cd��F-=RvS��ny�b��sTR�`J Q�t�N#�8��R�"5�\��`�c%�O)Bc�Gs�-;�3�e\��uܶ�*�m�c�˜�@�f��<�����Uu�ge4
��m���*�J�c�h?��V���wT:���h��t�u�d�h{R/ˠ6��&L�����M'���'-̇��>E$���Z��S��=��QS�I���7�30�Զ�1֕�0�����[��ŭv�}�Z�p�)"c���%�l���ˌn뜭ŧz��w� $����>�-��F1~i�?l������R;�ܗ���ߍh�kd�e�`in�?�v������d�"B"?��uz�R��Ώ��>1��+��*F�d�Tę�T���*Q��YS2ɬ}϶U�{ơ-z�c,�y��6�iF��}'�n�۟2�؈O"�H�b
(h�IG���1[QT�P����T8����@Q�UY���,�6����바�tVG�w�"�,������U	e�?�hde�s��K榕���Z0�JZ���E �k:�膲�EY�D6����Ş.Uo*�`�E��Ԡtc���{�ӕ+8v�p��柰ϥ���G�j����*����)�TjS�m|E���f헑hj,�e��h㷨�&��	7�O�Y�1\��8�{���%���&�I6��#<�a�[g���*n��6D���T"�2{o��{��E'���Yj��MAN��ʄ��B��n�_F�N����ԚM�v��E�efx]������5��/�Ƥ �~�܂bOX�ۈ�b�T��5*����҅m��N����kvL����u�Bf�M��&��z���T���;��ڤ�åÑ��kgd��R�W��"���I.Cý�q�ov\2����l�|!�P%�˭���� [+&3�~��I鈱�>��,h}T.���aϬ�9R�?��W�9JRD�cG� �vη�}^%�3��"�Ur�~�z?��NDgΣ�/d�@��X�"��uq �t�9v6'�
��U�Ͱ�NQR�Gک{�L)w�>����ʒ�am��"�:�
j�N�É"���[T�=} $؞�V���!ѝAi*k�����t��q�	�r���7?]�fO
T��G��̠K��r����Ӿ�A��q�t:K� �a�f6�6�����'-�y7q>�x�λ�|N���&�+p�L�`%�[= ��k$BKcJ%4�n��J݄�5�t�$��H��.iCM�����歕ڂ���p��=V�'ԧ�+�U��!�TV~�):	 !2_�E��T�\�r�P�cr'y��'O��^��U�����X�}O�xW����:cyۭMr�J�s/4��"�2�@�bCڞ&��m�$`J�F�%6����xaq��i)�ج���Ib8l{'�;���h���S��=��ŊX����_�:�A�����_t\4`�X�Ţ4��B,?�+Xp��7Y�w:c�IѺ�a��O�_�����!�j���T�5��8��",���;PK-\&��rw<�VA,���
��&���Q�>e<m��j�TQ��v��'���r=H3���_��m���L-���5���oߩb�O�2vE�QS1��%Mz$����.�`�x���%^W�n  g8hʋ�-���-"��?Լ��>�/��| d��M#�Hr%	����LD*�J����Zg.�\��P�~��tկh�8GO�T6	�I��F#y����⨙�����&d��ɬh���⤬Ɗ���gͿ5����F�7~̓׾gb��b�b������NW��?�����LpSS6�-z�,�Ƣly�
ڮkJ��1��eT�@�Ö��i;-/��p���!�}���~&�u%p�=�:5�F�M[T������4�Ω��o��-.J�Kz���$��G�R�X�:��|�Ϊs����cv��B�P�b٫�-)�6������Ur���KB��ؔ�<boF����#R�~�����NJ�և�9!ul�s[����pgyT_��v�_or56�ڮC}�Q�T43L9s�#g�>��˥='�þIV/�o�|O%�Z<���]�
W�0MI>#�{2Q���f�OJ+�$��eȹ �rbV)|�2��䱐>�	vw���y���]�>�!�:�9�h��՟ߣ$=�AԭC,4K��* ����j���p�_̹t��M��+W�g��ڮ���	�`��l��$�+�1�/o�?$U',��/�v�x�[f��))��9s34R8+�Pt��~sb��mŊ{�M����
\Y�+���X>�4s�#Y��n���	���<̷l	��j���9ʫ�=�<�C<P��(ҶB�=`�	d�����y�3��?K�<�U�t.D��۹`6~4_��ms]�p�Ú�ڮ���[A�f;�����u�&����,����� X�N��D���o�ܟ"�^Pnu�!�~�����vP#wY���߉���`p*��~_0�g0p1����� u��%�p���|i0���ؗ�i������ٶ��%LF��|�a�49����c������fh�Wy����xN��g�Ԛ�$,��ۑ��{��S�[�Y�C���$%yΕ���)����p������*��j!�w�廡�E�@�l������P?H�m�?cf��s7�1�`�W�O:E ���� �ܲ�c��￸`8�~6�P����~���I��zݣ��=x���4ȸ;�޹#'4) �0MN}nf�D�gq&�4E�0K� �[i���@^n�/���zr*j�M���!�������씼�ܵq�.����q�V��۲�H�;�.݆�/�$�=�揼"dDӴtڜ�_v�z��"䈛_�J��G����#D�{d��Fn3zQQЏd��{�`�7�;���Ra�7[�[�?���'Q��<V�:e��Hlע��tC��/��{v�B=xtq�;5R��>E�w�� 顙'�+�� R��Ԡ�7I�FŒ�F7MΩ�
1�Ң��2���ʋ�?P��a6p�h�I}�1zД�*,*b|I�';	1��W�ܧz���&=� �@��[�Dւɦ�z������ԯ9a&�zPVj�p#�C0�T�\��r)��|�iA렺1|�� }�,�!��l\�̧�����O���W�V���:ڲ��m�"!��R�X��������is����<���Þ�3��˓���h}�(�̺l1�Ck�� pӤ������q�fz�����_� s7~���r��ǚ ��ખ'�s	�R�B�c�J�68M�͜�����Qr"���RVi�E��������v�>k���/P�5峘��,��P���VzN݂��?_wҫ3\�n�w�)�V�yV~���\@��-S'>V��>��E��}0=cp��rSVW�u	7�j���H�(�4���N|4귽�f�.�[�W����S���?ޗS�"\���Kѝ�������;�8#l�.`�B)������ՠ����Yi�<�A�\7�-�z�
 Z�d�oi��kt���{P4D�jd��m�3����OUC�яxzυfm'�_eP�]J��Ջ$�^B�g䡫�o���s���/Ws��p��ɥ��Q�F
�v�^8������ �ڒ������}�rK`+���,�q���Ͽ�V���Ĩ�7�Ol3�a��xy3�#��:��#��R�'�n�zĿp�p�d�Fv�1:����/=�{DVTWZ�M++�� .��F�1��:.]�
�Պ�'�Q����*>�G��\ϔ��A׌�iz���/�F�é���e��5��xە]�*���w�k&ʕC���$�l�M(�~��?� @�E��Ԙ�`��1�S���?=��&���#J�)!�����sܶl� ����B�ȃD*�С	&���2�j@��A�AYee@�j�?��Z�*V�|�<�J�BC�I�ju��'`&���0�0�� ���CJ���4��K����\��4Di�`5�zK���,r*r�é��|�v�����kg �X�6ܿݫ�m�p����}G�f��\��&��㧶��m�_�a6�)� ������Y_�� fR����Y���:MC(|�����h�3:1ɳX�Fb�d���_
F�$cÁj��g���}d%%G uo��|T �Y'�J��U�����c��7�+�y�@���E����j@7}�9h��n?$z�Cn����=w���{|��Aݙ���0�&P�|�)��h�x�#����o_�&��H�-)�&h�&x>i�}P���)|j٭�Z!�3�_���E�&uS�qW���_0��r���L�y=��أ><�O0\Q(��Ǐ��\��Y��7���f�%�t��N��m�<4���<_��=[ᜈ���V�#a���.�k���XO�(�c�j�4)4���%��w�-�Ϗk�.�m�Y�M�����b�j�$ebZi���ѰL�D�?-ۙ�J�(E����dpd�;�c�0@�5���_��0y�5K��dlOr��.ꚥz�g��n?���r��	�����>yo�^�"�D�����wݚ$�Ԡ���#��.��X���9�^ED󓋅�ǎ��eT�+ZF�w�_��O�jH�톒�8�Ց�/���m�]����-
��E���`47��t�H@xR���'�����H�zu�v�@�2� `���Ű^�-��R�9�׀����?�R7Vܝ�����X���R�����(�v�"�QW�����8,��������4��=�?��_�Pj���>����_��f�"�tQ;�^!Ջ���v��P-�_�')�Vg�i����:��S~��i��Q��v�.*��MI�Z&�j��uNIEׂN��=����b��n��Qf-X�ə��k�p%o��+;R!T�_O`L�r܋O9=�8;�ů#�PFʫ�k�i%&w%r����U��*ޔ��7X�ޭG���O8���<tE�2�x;O�����U䮦P�ڬ�y,�(�y:�!�~n���t�E-q0b�	�sj���D��s��+�mG�I���2����:�9<cc0��$��2A����=�������_կ���Y��0)rR>-o�m��(���=r	Ϭd�_,n �2��.�s�Hr>h����,��{JҾ^!��ȿ����2��]a!v��'�mP�T��ؐRo�S6.EaSyɆCF�L&��5S\��]��N)��a�=>�9f��g���Lx��f�P������t.W;�8Q{bUݝ��-�B z?N5lC�'��k1��^�B#�0��wl!Q�=��h`I�{^�)$��	6qI���A��ZO8��'��T�(���
!� m��9S�w���A͑�-�����Q/=�o��q�"vh�R�e�NM�
3�))�M�ͭ��i~�(^��F:?f'UQ3���s��]�x�[��S�����lD�Epڟ=yt���=;j8.�������36�fU������w���/�~s��	����e�gLBQ9�6-�60<L�,�O�it8//g�.���^�W����8	�����f���4�'��n��2$�0[���ɀ�ᖍ&S���:W*��.n��F7=U��;��i�A�&�=ا�C;�Z�ŤuYB����fW��V��*��XƧ�����5�Y.]I81Ԫ0Mo����<�j|��g�$A6ԯ�o��N�ֹ>�Ef���-c~.�?[�Zk�NWq���r���Kq%ݎ�3��$VBUha�<)=��%|�t*ޤ;�S�
��́-�a��ư�œ��OB
�LZ'�웙�Fx����Y���᭵���z����b4A�4�?oY���ݠ�Z'�.�do��5$�;ޡ��I5�|X�e�4�m�-�ʖՏ�������"�A69�����c����_���vaC�D�1D�]]�%����ưUM	����	�x�	f�.v.`*{uʩ���m�#�<��	��o�N��Zh�L�X�R|��}S����� � �v[��q-��T%"�@��R���9 �e����b#�ڃ���ܸI��ei�m?�/��N8	�K-֢�� ��-��Y��c����U_+����6���ӓ㐊k�T���X����]�<�Q���a�A0�f�
���g�`��/�wp�����uPi�0q��ə#�\���q��m:өJ	$�͌�f�z,	�Ͳ��F_Kz7F�B��'3�ͳ-g	[��c}]�S��ш��4��:�ʍ;؆Ⱥ�n��0�?�HWz�B�`+\�s2��� ~�oY��z�?�� z��׵}�OX�(fr�����F�K����vb����"
�\�g�jc=O�۰�|�uz�n��mp�1˷/�5�C���3ح�X���^�eج��hր#����3�)�H)���"�"6Z������l����?������� ���9�ǑԐcvJ�wm���F�>�K=p<g�{+X���}�-ފ���"F+}g�ɩ2�xTc�- �s������Qp7W=�V��P]֫���^�%W�	�}Fv�H�����;ǋ�5��(�_y��9�8(5~�;��'zXT�;>�G�7��e-ئ?�7�u좼^_F��]+]���H��n��ab��'����F�[����X�տ���qgj�64�g��V5��/ ��S�u���oT��qIB���}sT\��c��X�V ��=,����4�%��8/�����U�_����v����h7����)kjI�$E���e�y�{bAO�F�y�c-|�Q�&���>�"W��(�9��ٔ��ٮs�����*$ӣ��p5Y\X�$�R����@�}��/���X�x3�Ό�u�u�`E��s�$"ه�@������s5�L���y}Ki�!Bg�� F�Pk\�%�|D{F�hv�v�3Z�&�<`�xi��
�Mw��Ɯ����̈́����Yv,���@����i2z���������9:��%�_�v�V|��b�2��A(C�[tO���G�%���iLΙʼ��6�y���W��+�j�a��[��^�?�z�� 8����Nm��o4|k(A�Z����6Z�[��"AQ���ቝشp��@��2Ν��NA���'���lt	���_e�Q��㷐������t���A%SÚ�L��dkM���F
I�R���d��?��Oe���p��L��K+8�̅�A}�e�c~Ox[p���n����+��U	-h�������el�(�S��T&��(�`T�r�+��$�O������~�`(���m��Av��̓Ӥ�Z*˳ҢbQ��~���v���R�Ku�@Ӛw7T�i���lc+���)����n�����jݏ.�Cc�h]����3�����UE�uI^���Ӱ��7���g=�u�*Q��<��E1���x1%F�})`���� O�1�4z�_:	��,v��-��E����+�ھ_}�h��<$�d�@h,�@��=�,���x����/W7
1��`6�D��{�q>�ۿ/I��Y������uiBF2��"	��d�ژWX����k�����#UL�ɏ��H��+la� ��-�OK;EJM�w�s��M��N�ոz^�O\��h]�g�����l��9>����wJ!�V-�s�hu1�>RR���t�0���ϫ�f7�%�Eh����kou�@�gųI���u���M�{�,!����M���d�SE��4�ٱX(ʄ*���y{�s�3�K6�T�ƫe�v&1�������BMi�~&;4eGB�]*@*p�/T9�΄b��T��7H�_�;EÊK��?��$(�
ġ����oǮ)ְ0�V��#�~(��]���0��'>�����6p$u0s>Ѣ��XfqTT��vG���M�N��dB����ޓ��[h��q�=�\p/�s�(�g��3��(wE1�X����DH�����m��8�I�0�v�u����Tid�"K%KX�-B�zn>䊆f_Ď�n���!�1i�u��[��>�WB6�t^����W���N��S'�_�=�(Z�| ���E ���Σ�uAIR�F�Y��T���"�-���ED#O*!!��F�,�b���8i7t�ۗU J�%���R1�8�����l�V�K�SX�����fЙ��6 ���Ml�~!�l�hter���a�B�d��z�f˖�,A>�� .���q��[k�5��i1�:�=��%�&�ve��JP�g�&X>��8؉��I$`�c����!��>*gX(��h#�;T[�z��1�6��ݛK_K��477�������X%Zx��}�Ԥ��-+���˳6���ѡ)���J��(��d�gØ^���c3�CԞ�E}�dtp+�>��|vڌ�����Ƒݭ%��n��%��s֛>�F�\2a�Y��jm"��LSbR}og��>q���nԴ��Ҫ��y��u�O%^�!���.�6b�����%�٦��ٶE�b.�����
N>XJ�"ׯ"�㇣FX�����8�(�����T"���p�%9�W��A��V{IR�@�G�a�I�K��Hy�Q,cؑ+ᰮx�	��I���%i#��O��E$	���g�84��kȀ��|vX�a5�mkK"�:i�Wy=�bb!��pWqy�A�}M��d�.�YE�Ӽˡc����d��3���c'�x%
fs���.�$ڙC�cFh��;5N��iޜ+��k�n��� ��V-�ڍ�ҿ�� !7���	op2����$�+��= ����J�Z-����WY�&��ں��}���jq��v� ��>�>1�o(�l�P��,�����H���f>��.��~F��V��y���@�%��:�z�h��Z�r��`yS���f7�LN#�HA�Ԇ�r��r���'р��Md\aqr�tɃC0�o�|Uk+���yϑ��x�ua���<��v�j*2qѨb��zi�C��`�% �jC�A5�GDz'E���!ijX�~�����״S��,hjVTkbX7����Y��Srs��11�X��P���p����\��U�����Ɉ-��Ь1b�oa��?R�5<���<��'3h55C�W�gT�n �D0��Յw[v��>2 �� �
�4�P��,b��,�^��z�dpS�-TS&-R�8O�й�jX��Npnإ:5�d�??<��$�M}��>�4�r�m�܊;�s�u�0��̶���Hk�2�i[4�]�}@�"�+e��\�XA~%*G�j���1�ߨ��,~iτ����oQ,�n*����O0$��<�fV5��1�i��v�_ZީaZƌ�~�{���H�!�W���� "� Xu;0�	��g=�*���ie��d1�r�t�b'4z�
%���|"��� I���UV.\�Î�֗V?G7��q����$Yu����E�r=[N	\A�Q���a�B%E�ǃ��M�e��pi�HP�؏�Dc�)�̐�R�