��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�"��S�&G�,3�+ c��s^�w�|�(;Dt��)ԋ�R)	Y O��}_�"��;�Ӊ������^[�Z���
}��Wı��/q�_�n��}���9SƎȫzP�����s.�b�hG2x��[�0�3v��|&���Sb�؇�s@�SǪ��jS�ɿ���R�Hp���.�;���q�/�q��UG��3�z�v�\���y�td�B��q�
�]E��k6$�)Og�-MU%��,k�W_�<F��(-�O�'bw�Yh�O�.��"eZ)E%
���R���~ENY{��;����m�X�n��@� ��i�1Ht��iB?�%��̞=�w�'Msx�"���U �zU��������Nh�D�m޷$�Gme�$���^z{��P �a!{�_�a�*����kD_fO^��2���$��D�)n�C��WU7��|sR���)drlDbW����B��C�+	7���[cHҙ�w��Κe]-�E�A�����7j���C{b�՚���A_&�V��A�O�n�������j|w�r���_7:^7��6N��]B*ž��7�)AA��iW������T �c�������GeF5�h��35��9�1^P=�*��q����\N�k���_fe�2��n�u^�tj:2�S%���ݱ�r�)u� ,�ע�|������^�G����J�3�c,O�=/��9)���"eZ�9h��"�b��2���v�PX�L���u	�:wv�ڢi��D���76zz�~%��t�fq�#�^k�N:/��J�(���=;�!Kpf�g,K�n��ajM}����JB�y�1n>J�Gr\��R훝<�������/�΋��]wAD;��Z_���tv���^oo��������>L� ws��s���J�����)��^�!��=�gҹ���~/}	��i�Md���2qI�}$;�g������ã(�o��s��wR�OM�FݘoW���*#�|�XU�K`���]y'�G	��-�Y�ͷQ�D؈0��i���Z�w��"Qj��j���# 5��5���c���Џ7<���
���ɮ���^F���B�vd��=7�&姾0m���q'�b[��#�IA�ʧ�Z0	�4�	oV�{��$��^�吊R7*n(���r3�[0�_P���YS_'�xm���櫿�ly�.yG�Mϖ�JlwI��l/��$�++Efw�m�t⮺Z4U��K�F9�8�x"eBCN��.񽪽ysUk�"/�M�,�AK�ٍ'�ѩ���2\~!�ӧG��%�!��h�8�T:@C�m�"��ˆꥨ�<dC�ޚ%ZX�������D��p�����]p���RU���*F�[x&.�)�<�$�t���;�Rҟ���{��2�,D��*4[~VaMD]������*�$	��ﮇ�2�L��9���9iuePQ���% �1�`�ϝ7��xI0~�f���%K�?�PPR}Vr���^�|���`N�8:Nx�L*�x�7�s���:���; �y1m�,�Ūe��*yˌ˞ǆ.V�!>��XY!�+�#�
	G|B�k�[@1@&��5楮H���E�v�;T6�_4����E�Ž��+Ԃ�$Dbgya�����U�ӊ�-s��d�E����K���R��3�V��yd6-إ@�6a�'�W�f+�~Na�/X�?�3-�ɛS�� 2�2,�� ��˽٠ˋ�FuޑϿ�E9��̠������aΦY��H�)���<���#p��v�Tja��/Ś�V/�m|��d�'�z��S����?����J,0)4�+QT��??��,����!v{n�G`���'�R�=�c�:x ��uA�J�ȱ��ߧC^ܱ���D0/��Gc2�#�f���!�;M��}{� ���Z���F��dئ�FF��kRe��d����<�����0�S��MJ����+1�C�I��	����!Ih*��ҷ	�
�o� �_�4�3��&E
_jY��&����&�l:4;M����ݯ��Ud�kuL�V<q9�%'�^�y�Ε�r���D\�tgnː��-�����>�b�}��1�Ŏ�
[���WJ��|�xi�Yj>�7�A�B$S}����czKz���K��ŏ�~ηVo�A?�O����˘��Z���3���@��O�63������b���W��y�n	��V�PDy�Go頪 �n-���⃣s@w�2��}�󊵱c�.ڀwd`�Zd��CRK	e���uP���Ao��+jW�K@��jf4`�q�6R�G`�B��CX�W�ӱ�x����Y���~���IJ9[)Z�q�nY�*YC�DY]��PZm�vT
�Z�2�<��)6���Y7����'[����Kr~
%����A�h�:���i������/ڋw�gGO��x���p�i�7��;��(^��]�)�tEru�)�(Ʀa��A�' ��A�&�F��Q�`W��A��c&2�U��;��h�P�D�=��Kbh��l��5*��Օ8�Ͷ/�xh���*�Bԍ�}r�K�]��+��W�~7����C�T��?�Ơ:���Ȼ���s�R&9~SKdO�ٓ�?�����e?��b��r%(fJ%s���+An	��^>�Œ���f�T����2
af鏊Pˤ-�?Xm��V�+pN�s�������w+B��h@�9�`�/�����V���2i>��-��Z�����*2bFE�R���I�dٗ���jqr�̠}"L�ȍ��A�2�&n�2�fm|�[�T�	JX,���㍸�8[�P-�1v=����S�K�S���}���%H\C*Z��&���ж��Z*����Z����Y�o��
zi���)o��"d�!�r��o�gQX�(�(��lڻ��r��]B&OYS�1p��-(�d/�~E�"�~F���n�GOiDd`?#M�w59�Y��#QT�lb?Td���v�g�sꜥΙs��?���e��X˩+���&~٫�@<>n���Q�8, ���l2�c�X;���@���@�g������s����v�aW�"�]��ȡnf���Y�����O���q��qQU���5���1�+�&�V;�y�����B�_���;������&�#Y�7�{���l�� \�L��k��I9aC`�Y�'A���E�\,��2��Q�h�<����甶)Y4)�euu�9���L�k��y��]��JKѪ7B�ܝ9a�~x=6s���f��2���A='P	�[�77՟�����5b�T�kN�.�,��3�]�Q���3�Q��j`v�f�}�>�1;�E���d3=�Y!z���k� :^�=.jN��(R#�ۿ�=@�.Xe�1{����ϕ�2��g��$��z�S��.N�Բ=���Е?=&��q��`k/RI~�N����^��6b�W�֑�p�V�����
�[n�2���-(�%��q1�x-БΨH�1o�& nA����@.Gk����a<�L(M������:$�5�k��a�g����f��9\֦Ԝ������-���P�ٽ�㽐�R��R��i�}�������3�Z �,���KȢ/��Hj����Qk_p5u��υTE��C�""D>D���*0���j!SX���05��F��Om��6:"S�+<9���*S!l.B��k��
�s���z�edk��N2��[��q}��f=izt�뫋����:T�Y��$,x��+]v-��27dp�5)%���Dy�ڻ�1��qs���ۧ���`u��o[��;���xI=4-��UD�P��������7�DT��4�=���0��Y��rzd
&$��T�f�&����J�bxX�̃J��3D9,z��!l~�� ��1��iy���pW��T�o�4�sAy� J���� �o���S0����Pv�!_�NbhS�Y�iK���F�0�L���3�}6���[)1 d���r'Τ^�l*FOi:��
����&�=l�b�<dF������7��_Ħ-�NUxϔ��&��>]�:;Y�_�{4��*`���\l�0w��ç=�7l-�3��nuO&�A��X
�׀i?���E�SN����"1�>��ķ���t�w ���m�S�T{V�+�Hn ����/KDqL�<��7/�6��xo�&H�N~���F���������K�c�!�F��p���CC��kW=�-�F�g=�4�Gذ�O�HL(���_"��Ϭ^ ߧP�.�;{�yh��HU0�h���9@�Bzc�F�],�l +GJ��"���i����d�~��;F�7h���f��{d�����:m���+]��lfB�{0\�T}r�{�5�:���=89�v����`��[5�>˹��`C�W�ݛ'9t�ڥc�*��$�n<��6�� ��*�R�M��`��gljr��H��&M�b�.��0�VV�ȅr&�ס���"�0m��ή���{ �'$(t>;XU��x_��� /{��1���z����X|���$�w��?���;��q��00��Rص��H�uk!ִ*��n��w�V1֦f��� �{	91Kn�r����t��'����X��@	��_b�R;�_�^4�*�Y| �}ȋ����i*�d��n��:�^:���V�+����[aU�F�\���z0p�h�\3�ں���"�IU�}A9O�鑕��q(��b�,c�tQ� ��V�������(#<��	kBE�
Kx��^�HS�HՊ��f�L/�G_����_��p�Ϟ��� G)ի�M�'hܩ���Yn�:�:�'��2�N:ͶRIv@Գ�{٠�q�-|�}!8}hϟ��x�a����a�I�f��<�R	�oDǯԫ���o��@z*r=�6��k�qA��NьOY"
X�Fyq���H{x�8�ʜ6x+��?H��P��ed�φś��Ne��t]p����)�~��fC�/ihn����S<5槛�t�]q���D<܂�R����>��qD�% �GCv�ke�����+��8��Sr]�t�q���������SR�}z?���t�M��6�L�ӡ���F��P;�;t@�l�sl�Fk|�����o]�tԄ��~���Q��&�u].Hj!���s��.� k4��52�5ɺ�xm��φckUZ� ��T��lu�d$ԅ�J��]BO{���%*L�zA�4#Lp�2�g�\zϦ�e�����r�N��M4mM��<t�w{�\�F8���<ڦ��k94RjSh�[\�I��{$D`���0�&�}_j�KLE�����Ѿ]���^�޸�{qe��/Ͷ�V
�:���*/*i�k2�-����I�������������wb��.9#h���
�J]ս��>�u�<����/�D�NDǸ���^�6�j�9<r�}Բ�P7D�K%]� v�J�۴�N]�P����3$��p��,�v�u"Q&�(��"M�1 99��4���¸�E��*q�uj܍I�}���p�����߂kù��Bn�<i&M�����/{� :�TO6y�X�B���x�D6�D��3�_���%3����=��b�f��<��+%Y!	D�N����if�䑸�/�#^��Ӯ��7�kڬl �<��I��r�'p�J�����6�Xh��,�5�1�����������U�A�HL��b��l0p�(��|o�{<��#�)7��h_�WV[{��:��o�����i��|ǵ���Aod�-�a2���B������0���^#d���n��s �p (*���-醱cĮ�$c�� ӽ V�syիݓ�`AB�Jg��Xd�J������糅���σ�\yA�2�(f]'[sԔb���}kv��N��J�l!�\�"� :ɠYlv1�п酀��f�d.32;e�>����*��	���x�
t�M�h1�{�MؖG�aZ���d�0L���U�&��~���l�~�
ޖ�`1��?���#U\QaL�m���s�����ݩh��E濺H+'E��/��1��7���<I�ݴ�=���,�4��F�CC��߱�����+�W,,)��s�y��*0�DR]zE��� �J`����e�be�D�Ԅz��S0�o��;$��Fȥ���*),��r�*Ay��P ]��+h����9/��P���
[��:�%�fz)�mbd�	?`h��W��E~-�(�(����	h���_Ӽ�R�P$_��o�J8W36���!�����=	dM�Q!'��W�� !3�_q�0�� k���EU%�2�Ƨ�i���Rf�Il&0��>�;�`��_�m�Y��e he�\����'�Ȋ2u���-���	���x����v&��� ���VaA@Ӗ�\�q��d�f�vP�e����ζ��@�ĶW|@�	���-R�>�5��-������+�P�[i�9a��_�$�N�9���J/	"Y�a%a�)�J���׸��u,c�G�Lv��=]0��Ӫ�L����S%���,��Y���9���c��k�ϒ��艱�,�����3Xn	�8�j�z`��7�j�Ψ^��};�<̳	�u[½SEv-����:5�H4T�f*���g�.��-�j�\IB�N�>�������R_͟��R�c�
s\h[ZY{��]H��Ј����1'|��b-�8��%߮� ��J+Z�v!�1�C:��73kNa�ǚ
H�#UaW����E�86A[Z5�����a��gX��Dt��MI-&�i^c:.���}��ģn���hĔ�C��\\ �4�����ײ�X��;��wR�t�=� �K�S9��A	���J�+�-Uq��d����x�+�$?�vy/p���
Bzs���Z{=�l&�C��N�u�3vN*_��/�mG�$����҂<�E����mf�|�龗pL	��z�Ú�������AJ��w��И�$�����cf�߁�<���U���`�5X��:�m7g:~mX��e7���ؓ������h@�����>����-1yn.�І�ܟ�<�>��a��Ġr�+<2���\�j�hHȿ�
�2���v��1^6c;�����U�\]h.�Ym��
��s��0����>���
�췟<L��s,�@=!Jނ�Jֱ��\5"Q��m�������α�r��=��`�Jw��2���Q�<�3Z	a�A�/6������sYQ$t�����Nd���9	�&�y������^=qW5iĸ]z[y1O
��O>L�"�]�4T0I�r�}�R&m%x��͋���QE�/eGװf4�.$���/ۘnP���'�Tj��pj:�.��3�o�bo9�OD�]��.�������b�H֥T|k����SF����p�J�LO�(�ʘ'�)��vA�E�o�t׏��y$�`�>{SsX�-�����ʖ�Rr�Aط��>�oW^�T�?=��J4z��,���V�����m�H)m��'v|K��%�5=E�KK>>aZ���2>u�������M��kDe��p���>��b�B[>�v��Tex]7��7Ny�{�򙧨w/����q���w�9@Tf�%��E��"����gZ	�!Q� ��|C�έSu�W0C���۾�m��|&����%����<�R�rR��VDBWN֓'9�s�!��)��U��
g�����1��J�ǃJP�~����v�	�ϯ^�!\�0����	���Yߤ#���/޵!�x�U/�o��6T�bb�[�h/��,B9��x��W���(��^��9�2~Mk�C��
H�i��(�Bf�㰳f0=�37;�ƙ^�����Qlx�4�/r��+���n��m02�S�e���`�/������Q��`s�գ��~<��ZŻ��tt��/���z9�O�OL22X�ZN�E���W�~�kD�o�����e�?�!��3��C�Ҡ�](<G�$a!V��Їx[���&҄��6�e,�r�����>�27�Cl�|,]Η.�4('�DK��b��<Qz!G��� �n'�5]�)�*+�R��?�;�%D�HR���Y�DuX�b�o�`�5@����X/�;6�5��������M������zs����7N�O��]dV
�̼?e���6�[ �[�0�4C����r���Ҹ�1��
e�d1�84�9���^S���wy/�s�RS��ip���(r�q_}�K�mۉ��,�l[�ֵ��Ȱ\��Y�gjx%���B��5����[�7��)"���x�듧R5]-�̆��[&���3��N��,U����}2*)��[Mv!���;�� ��U���<�Y�W���y�8_�	g0�,���|Ie������l�q���o�	����P�=���	�k���*m!����%�><���y�%9=��ux�!��L�XP�o �\v#�1��^������Z�Ow�x��B(,=��Qe����u�i�+GCz�~ �Ij��I�|RTKp��_�N.:��0�[�9-!p}��5�/<.�k[ľN��T��h�\�kJ�-1|(�^�\�JtN�ͨ�e���	i����wCP�^�U�<��| q`�U�gh�M�- d�۫�	�r���-3>���dB!n�'��u���n��ߚ?T2�b�T%��Y��a:v޻��%�!���3�˃1s����=�M��?m�
;77���/M<P���uK[	[�)���;K�'w����3P�PL��L[�~/6��1�A��FCԤ��'�����P[eT��Pӡ09F��4�$y��feZrU��ԣe�ɯ�����h&���+�}�a
�kɴ:1�!�w$�v���H�������[y�:��č,��bӉ��utt.le b�2;:�:�N͎�{h�v�+�uAh&��I���%"g�G������3B2m��96���^�2 
�%7�n0K�B�+ﹻMk���{,"�j߇tUsf�쌠�4h�Ӿ`Ե�O���oٹ�4�E�V)J�|>	�K������^�=�!�1&�����7�b)�U>1�e!�~xS^|w���{�N��ka�_�z�J�0.�/�n�@P���.�j����&��nŎĘ(2i=f֠���h��x'�&3�S�"/�>� xA0'D�����VM��:����c����0�;������1�w"����>��&%qQV���7�+O�B�N?�<<ys�?�+��4ɇsU5�>Tk.��䚓o�k�,"\�U+�l�JV.��ǝ��]?��D5�G�l�n�S�Y��o�X�����@�����[�n�ФnpU$�]��V��@�������K��f�t8[���JA[k��nm iXڋ��2A�DT<�*�I���J��y���LB��j̺	��XC�j����tac��Q=\�s�K����/��W��}߃G.��Q9�v̇�8&����:����-.���E\AM����x�%J����v_[wcpp��k��qE��⎆�zJGԌ'?"	9�&⼵Ȱ�ދ��5K�e�vv���J���|+�7��+��Z�ʂ�[����������KB�@v� �����/����?���[h�����*b@	W��W��!\A��i%لD����=�6�Ԙ�6\�����/M�rO���"�x���Y�B;]��$��% �o*#$�9W<u��}u\ԫ+]I�9��gп�:��;�ah˻�gN����J�I�����y���;.�H�G���R	se#ﺹ*�<�A���n��@2��G��H~�ʷ�~As�h�">���lT�E]?o�W��Xh�9�~���I�vإn�D�}W�?��E�"�97��A�#�������@������d���:Yp�#�e�j'�Kx���4�)��t�kdn��B��������@{�y�����5UZQa�|	��������#���ٸ���1�vN��}��^&b�箊����_�OL��$�}d��,z����U������b�=�u�ʉ_�ky��t~�?O7�Ќ�d������nb<h���?P�ke���'4OW%����*h7�&R?g�G~J����X�K������Ӥ�Gk�nkHPc�_C'bYc��C�<�����,z�)��ʊ3Ç�9H��ye��{nUW+�t��n�>@V%(И2��) �,8�v�[�p]VPŌg�Y&�Z$b�K���I�u[n����a�m"��DϨ@�xc��?�����(v彉�P����.bU����]��2IQR��~�~�3��-��v"�먣���<����P����0ƿE�j?���ꈖ3t��{8��G�|��Ve� 0���x[x)s�
��~��r��/��q'j���/�M� �J���K�	=�]��qg�)���]�7^��N���uk�7�Q�^oɠȸ%>���ѡ�ik�*2��8ۧ�%xb��9��[�޲�P tW��S������I�JG�a咩o9o�2�3�}R���*�r�g�h>��R�m�.Mx��>B8茐��W���c���?�@e�V��S���/����*4K���#,�A�ݎ�h��3�+�S����'�&��խm�t=+��u<�Kʬ.��؍x�ûA	���}�,`�S���2��7j��a��0Uؖ�Nm�;�1G��Ͱ����CW�D�s%ц�\ǈ��UF�N~�ip��11�n��3B�G�7�����m �ÃX͈��y�)�����9�S�����׽��{�1J85����<�o�������÷/��+ǝK�Β��4F_�0����.}�.ė�H{�&N��;l��[��!�Y����� �f[}�x㟹%S]�����O��+Ev������q�u�$q0�cϔ�"{$M�j�<��U'f�?0�N`�+,����Q�?��N����x���0�F�� �V��>t�H)	4��Y�oi�`,_��J��8�2v���n�N^���f� �mB��� �U]�܆����asE"���{��."96�߻����p��2����g3��)��z��w�6����E~AG<�3���/m��t^�eu��?��f¥����0m�*/=l���[ж�7��93�6^�N�L��1<�F�C�E�+}�X��]Wg�=+_��C��0|u��$h��������2Aӽ��(R.�j�)p3�����>H*G����F8��[5�Y�w*4��{O����-�[�����>�����N�w2ݿ��.�7�4s�C�N����m��p?��P��h�ve���6�!a�ct�IY���r�p@Q%-�Z9˗(�Ȅ� ���Kr�c��b�OiKi��O�����d�Is�wI��u̙J�U��۬'s�����0�W�Mb{&�*��P��f��<���b�g"�����;c?_�5�K��<���
��t�^����MS��q�S��!_g;�M��Y�s�m�����(���b�����>Fy�>�V�F�q�w���d8�������}��K� (�	܏qib��b�9�W&!�uZ~C�.
�s !�ڙcօpX�ƒ	�:���� �'9k?�Xdl
/b��x�;ٰ���u��I���I�q�B��*\<$;I�B��$����Lk�w��[��X�uizA�����$�Zt��7�^\��J��a���1#����ュ���K�f�AW���C�Zc�,�w��s���e�l��� ��6Be�
O��ZٷZ��ZȌ�"���d�Z;�
�V��u�OT�����9'�[ʌ�L��m҉�b��&��������hK�S�El_�� �{KraXv�P�nWm^���Ʈ��k�4|�m,l@�ho?D����l���v
b[L׈���GU|&7���;�o��X���)"��(��K�� ����[�*R
͔QD˦��f�x��;��aIaC$H��g�*����⥙��U�aФ3��B�T'F����V���6������P�(Jn>�r���p~#������t\qO��'�E�-�X��Uy<��'�]�k=�Z):�U�*�����/]b�d��g �rR�g3������#z��ym셋?G
(	�W��$QT�cȶ(�]�u�	��f��xgG�"���H֎�A4]��g��O�i������5aH��l����w�r��p����� X����� ʩ�ݗ�7�@�[@��²g�J��s���-ցx�0�&9T&�4@ۨ���ԏ2�nF�	;�o��<�������R�_������ͨR���Q�����ږ���y�Pt��c&{�y���,	 Q�\�X7Z꺼�)��"��L@��d��.�=��Io|���am����2S�g�4�*�`�W���i"��֎���n���0��RG\�*���1cx����|�}�Q*�x׆X�3��wx�PsU5���`��JGq%}�Q\�v+���o��&��#���ډl�Bm�,��቉撾}FQ?��e�~Y�;�_n;���B��I,s��g��uS��3�4O�F)}bd�U�X�d�tn�d�9n943��u�W��N��T��]bΤ���cBpzn�u�~��)T���Dr�>�ŷ�,�g;-Ksď�Zd�2��إa&����xf]��l,ec�����*ͧ�Ӌ,��U��\��B/�cd}��R}/ː�	�kPEA��~կ:�W�����`A��V�����`�K��.�5O�}�)&����FZ��*]�~D~��K�$�uQ`�g�.Օzec�R��+��@�і�%�!����G4(s����K��� �{��{O�Y�f�xr�u0��r��@M3?��jL��� (u��u���T
�J�{�$����_/u↸.��Q6��f����v���Iųp����� ����%����-(]Pϓ�և��\�ܻf�_���l\.�KJkP�M���D�[�R~���O9ܬ<0՗8&?�ҋ� �& ����sVQ��P�rEV	�5��H`�vS�+Ҁ݀Q���"Ѱ�{��C���[5��Ψ���%yC΋�Q�%A'<�[�0���52[���m���^�H�7�����zgFR��hm�m	-��7�t��~���`teX��6��C�WZ�̢6䪖���q��$�z�9�ʚ	�}�����?^r
�׏��s\�S�\��(��7-:[�'���@*No(�qf���s�3�s��H�Q�l,h����W�3�}8��fd�;�
aX����0K��������_@v������o+<_�?�ZJ��c���m48l���g��	G���tX���J����5༪G�n<@_��u��5�Dd�̓�E%�_�����e��/�T�IooMa��9;UWC��4� k{���#�l��R��z�=���{pC��w���u��WO|�֌3�X��R�P�f�{)$�#9+���L&]n�*;�1T0'���bk�Eu��\�=��>�`�Mv[߀+�|�-��A��P��}0Jc���c�f��|��d=���3��O���D��ˢj{R�a��IX1/H����e��׍�B���ٗ`�n~lL�vEI0uOu>��g�<t l��\���m�@����ɒj4�~f�� ��	ɶ;� ����1j�ȝEo��iֱC�ytJ�i�5����Ըr;։�P�k�jwN:_���К��[0Sg����j4�Fb�ܶ>g�9(�3qX$�`�/!��3��HZ2b�����{�_a�)_A���5�b�`��(�mj�x`R��(�J�N!�;9w�h
n�m����a뺲�����%m�e��CAOd�p.���X,�Z��)��ұ]oX$p�8Π��B�6��.��.�V�9�=i_,�sq	�s�RM,Ő��,+��U�]A$�Ľ��D8GsW��&���|�:��T���߭Rv�92�0��}�@h��8hm3Lx�%)<[���)� �;�7-s��눾l\�N�V�ҳ/9*m,��	c��9�*8������
�g�w���~�_ו7
P	�,��k�I�ٯ�l-�)3������ڴ���3��-�}�W��CU������r�t�"6K��P��=%���*&g�АҦ�/h���:���cϕjס���¨�Ag?���LU��R�+10�J�����w������BƘ@{�:���r��`F5�&��=u��h��{G��D#w���T0�Ta�g�a�
Yf����6Ba���\��HF��3ˊ=�
�$�2^82�w
LEo�h��&��zXf���J@�[:>]�J}D{�]SHR�R|��rk����zR���(Pwx5f�/�>�5=Mq���%�u�m31����~�>��v�Kh����m��LqNޑ8B#���i�J e�e��)�>�Wr;�'�%�JW��8=�ze�i(�E����O�v�p��e$�	O
��D���A�G뇖C�km���o����\r؂�+���YD+��-U'Rz���/�5�Ӂl����b���V�����%�z�)\nJN}+=���Kdx�zO�VB�&,~f����X�a�yZF�%���w�����NkpYQ(�(PodA��
������P�{�i��n�z���f�h{�՜Q˕çTK��5�fh��֮͓�L�������X��hǾ�
dUHJWН��V?�E��VZ�_�T��8�4�9#�4�3կ��Frn��Q'tT�8�A'�+����l`Ćs�{Ջ��f^�t�i.�g]3w����$������­��ꏹϾ���� E�-/��B���s0@�(��>;��P��B��܀�g��"�u�\|�uX�5�Fj-�m���e:o�Kr|���k��	�D>V,҃��#/]ғ#ՙg���U�Qٿ�4��,��=��5#�X^�U�
��e�%�@�#�{����|�Hy&�r��u�IL��m(�|��p���U9�v�ڂ�����&vo4ލ���C������NXhx�	�����]����$;~�;K����<�E~�"�?�L"qW��3���}�a_�����Y��_���ΏE\L�]���
||�f�W���Ϛ�V3+�1�%8YД&���i���hc4��d;.Pٮ)�hi�|�M:I
��·ś���^�(Ň�iR4�ap�� ��W�7�1>]���t�6 űr�6���\�#e	��Ԗ��`3�β;�k��2��	�P{�M�';TA�6�k�F2o(j��R^�kd%I?����LD�yŗ�\աjQ��2{��15�ꗖ2��U7f�xDl�f��"��q�q�B��r%Y"P����m�҂֧���'��4̄(�|Xpoᣓ@��L��n���"V�
�=M:˪$�v%�z- t�ȍ
��P���T��-��a�|9���+�y�P*����sW��2�krBD��X�o�[
�ƣ�g��?�]���>ɨЬWlg{�^`٤M�����+\�Hӡ��~��f�#0�C�T�	o���Z�^����ق��xA+&%��o[حjȸ��5Md�8�]�;��B�;L1v#�zkܻ��״�dL�T3k�guU���ZE���N����ic�\C���1�҆��/�)��ʦ�v�̏Y� Bh��-�����1.ٰOd]���.K`@�xx��e�E��e��V�_ȗo�*�<�x�o|.�󫳎rZ��&[&���ܾyB-�>+�4��B/�D,������|�[¢�����r�@W�������bm�,�b���@��q<�׵���Y\��Xu��)"�^���}��f��kg���f�Zw�^�,���7}�x��>��2߄ڳj���Tb��"�7��M��:����f���I���1�<�EF��Z1��\z4 �7꽷�6Z��J���8fؠn��d$�2���3�=�����E⥕{�c�������b�A����h<i����6����H�a�vm޳����W"��.��"��!�jDJ,$5~eox�A��xk	���(d�g�]��k(!է}��M��@f��Q�O#�l�D;�A_eyn�P�C��h�y@=�@,�ˣ���"p�,��Ak$;����	�	���Yv�Kŕ��@�-�����Yׁ!�	{�O�,����KG��~c����������m��G�lC�P�,d�"��pS;:��Y�����S7aNv��gb�C:��XJ�A���"���]!"V�EE>��\���~�7&#�8b�߻��ua~���&�$x�|˕�$bb%�24���"�_\�W&a��n�����ԃ@��=�ӷ�Ձ�;�q�Uy�.�V
0�py�����Y9�Q5�:�_��멲L��M�kʈTQ��m6b`�ͩc�������)
���V�2o�XǦ�.�fmO��{�@�RǏ�ۍ���wh��)��Tǝ����W\��j�s��ϙ�I'��6�N�^ߝ��׺�ģ�n'Le{[�G��8��L���!O�����,��΂n�����Tq>iϐ���uy�ٲ�̤���.�j�aS3�݊יkj�������>&9J�3��z�3~,�0���J��M��X�/!��Q�I۩~��z��z$d��#���C�K�oi��o�c��d^��Yh�Jnut��X���N��"C(��6֜e�g�$��s��q3�[k7�R��/;�F8��'m�q���`lʵ�폻��o�,�V&����y�H���� �|��|�Ƕъ$�\h��mTtՎ��8�Q�Z�~mv�R�ye�1^�d-%�gY���s��Ě�w������1��Xp�$��Ѐ}�g]�"�<�\�×I��.`}��de���36�����*�9Ef'+{�����׉�{'Q%x7�V%���Co	�h���n)/�Q�����!U�fL�U�V٩���������.�:"�_($u�zv2��*���t̂s���T�Ŭ��6�����a��6V#*v��T���m�Y�F�O��ap8R|ޛ�=�]�X	>{���Z���SkCN)i�D��]#�����$�>H�fX(������~�-�*�߭��]<����mx�R����ܲb��t�*ˋ�d�]ӡJhŦk�������`'r�4A���`�۫&��'I����������g��S/��˖xt+Z����~w-o�=�:�?;�'��C��u�����\z�f�'C;�>��1���~ɹS��힘P�}�uܜ�������	�����^������O�t�9J�D������{�5wƇCobqL䍗��#^�b����m'*��O�Ǡ�7��yT��!���$=��+(�%�����f��/�����c��ɇ��ϵ˫U㦈�,��+�EP婆����}�Ti�Y�o}�����'Mn���� <`�1R�@j=7�n{B<U-M�u���#~��1]=�b��/�jY\2�r�3_ �x�ĴQ� ��<������]���7�P�8[�iųИb��`���>g������a� �ʞaAU��-s��[������� ����uß����נ|*�	Q�w���,�,8��j�`+�o���Ɛ��8�7�����L�Ejͥ��$���/���\�x����_��}��Z�y�f,Z�S�.�U������ä�q������!��@��DF%�1X�R�z��@z�C
&YTs�m[�>�OC��AM!W
���?fc^�-_�u&C���|����in�7n������������wLV˔Qp7�(�uЉ(�yieP��T9d [.�K �~o4�0S�*5κ>'h��<���sV��$�Mo�Nq#e]��%$l��]�kn��.?kܝM(@pn��r���e� 	�	ua%k��Sg�(�E�G�������X�m��Fw���M{�Q��s'%
�+�� �hv�(��)���%��O�R�\5XLArӀU�*87O�R����c��l*�P�⬏��'e߆Ao\��@� ���ϽM�LSŽ&D������蘻��՚Q���M������az�YN��܈�A�C�J��2/Q�	�����ȫ�[Cӹt�ܼ�;uR�T��rϰD�~�ν�J�w�*���t��J��&AQ�i���q+���W�Z�&�]gu��襚�	6����9ӧ��m����,J�/[D�J6�4YA��c��i���4���"0ʢQ��-�@^��:T��x-r�}���yX�"�WoϜg����)e���֡V����'f���i�J0���)���H1�/<�	�h�^�$?�+����n�i�M�'T%�0}EF��!6�ǝ��8�R:��� ��&X�kJ�]�M߯�o�� ��ۿ���0���'�]����6�I%�i�R[혊�/�HC7�$�
���1S@N�"f���NY�\Y[��V���iQ|z��<�(Z:���9�^A�o���ak�|	V���v�mJ����M}��V�|T˜D|�����s�?ћ�LL��C�y&߅3���2S%�
�&I��j��6㶔��v2��=����gh��E�&�%�.@[�#��4ۿ)X�l��Z�8�Nw����|�SZ�Tt�/��b+�$돍%�1�e����,�d����+��v��
�U�:L�2����|Ю�Tr�rLG�A������X��p��T��$��!�ڰY ��U��qW�rb����̜�J[ƥ4�Ɛ�ɱ+k5mE*ZY!-&�o��Du����!,	 a��ILЦ�hT��g�ώ��Z��{<���CԘ��͉348w2ײԄ�B��Ӛ���R���XY��=��ؓ0dE�[�Ԥz#�ِ}וR�4aZ1[ ��Nt�d;SI���jcR�+�L�����/�LEb,C��v��}��%A����3���=<_0�J�u�G�N�0�n*�P��س�:���r�/GˍHn��}u3�Y��?=j��(!��o�����W������~�@�'mfL��W�`��O%%)��
��o�Bk�+@8OV:�M�z��t�`��8>�����*�~j��Iu�[T�أr��p1P��ڔI��Y#[7��mM�Mn�R���l����) MCX
ji������A�C��c���-X	�4�-`	i�����I�?�o��F�&��T��Q�s�=���[4
d�������@����{9ٹĈE��]=Ƕ���^��9H����/�����f� 1�=o{eS�,V�,�C5L;�8����g�v[�	Z�I�s��/���I5��W����P`ČOexcA/M�ˑe�4�an٘L��H���_Mt�nM��ţ�C��#\�K��'p���s��lQNټ�W��b��M?قxwȜ~qF���[�>����d\��de�RqQ�A�Ļ��&()��k!eզ{���~��B�Y���T��Y��t/���M�j4�_�W�k	}�^y4$�׍\��p3\�x���M�Z��MMt�woaB�ꩯ�0�Z���#��Iz��]RN���oz'l�$�Ŧs���`���=Vi�A�\Lcܢ��D�yHH�>~ۤ���2��|�r���I�T��g�{E�0��l���ɩ����_��b��Y�b��
Co� P�p,���؋X�~w��<"��$�ᘯ�/�n��pC���w:}��l���0���K��.�`���y�W�=ZI���Jȑi�����/��LV\��	p��3����*4E��XxI�����BW���M��+{��WL΅�'hmZ2���"�[c��a��P˸��(L&�H�e����5oCa:U���v>(�Tb6J��=�}�syY�`����W����G,�9������i�	�p�=������0�QL#��b��UVۀ���ww<T8*�hi��C��4�[؅�!�:�$�`�������/��:ZW���&ɂ��(�Ir� ��53�rp�Dmu_C��>��i�␘��A���]߀���<:R�70����@k �w�)$�
�!h$�m��ӊǪ�>lCrE����-�`���=j��3T2]1;��AO��D��jF�m'r���A_s���d,Z3`ۤp��2��F�:C�fߐ���dF����{/���5gɱ�>��X��xR�y��Y�M��B�Sa�^�Y�ctr��Q+�u��K�%v4��T���}�����v���	R���W��ﵸ�����D����D�Lt�x�������Z���O�M�E�+;�Q�5��_qY��w���������qAAir9!;:��Xv���0���Rr8������7!^P��<������6��p���ʭ40�喇�R��mghd2�P��nU�DD4��x�����mg9�!�5���ǎK\����.���$n_�o����gGA�oH�ډ'];�Z�lP�S]
͉O31��g*ߛA�6����~~�`qPM+������C�E���&���#`��d��txp������Z�2�ɫ	t�8�Փ�!��ist�#Êت���2���m�����NNZ`Րh�����18;�obe��zC�Og�X5�P+
	���A�(�`��*�tP��$5�%�@�0���D�?~�����k���b4��Y7��c�"�����\����5�F�@>�0�ä�~H�H$��l�Z���.x�Xh���3c�86� ;��^$b�'������R������8P�$&ͨ�ąe�����U3���<o��L&Q��m�~��:QX.�ؗ)��<b�ؤD�WY�����+돖%f[�=&�D�CNĐ.�nZ?e�4<1 "���Óͱ��� "F��e0�m���%��a�)�+*���F};�#�����D9�8�1QT$C���tK-���1�;~�'�1�Zj���L��x��D(��&ejt$'��|*���哺$9��;�ͿP,aZ�L�(����E>�Ҡf�'��1������#��f������I-�*Q�3\�� ���Y�E�v��^����Dy��.y��Hbz���,@q�8��hȲ�Ue��4[�ﭐ�`��Ь�h�u���!}��s��$J�C�'�ƨ���CdC��8��X���3���R��41�G*��;4�����сM��c�*m����X%�T��v����G$SW8���w�U���k�q"�U�uKK?Ɉ=1����:r��� ̈́�"��eV=��4g+��]��"�o��]��8A������,T�HM`�6& �>�H<��rS�Q
�R��V��}��ӽ`�S:����RQ�ʦ��6#BbJ�gZ]C=��jfGp|��CUhu���Z/<d�U�է���C�U�� >�gXI��+J:�'�)��D�
�X�z��up��j9�Lք�i� l��"ƹt�m#��N���z���H���N��I�;o� uS�������3��趟��;�!x����ڼ9�?�ֶ�1^P�%˒4j�B�w����)��]I�HA�&�m���$��"q��D�`�8x�M�t���*`����K�H�n�6:���Cj��V̷��vt*X�9��)��HP.�`Y�^�@���T��U��\��Ы�f��Lp�{B��Ǡ[;�/\�*��mz��S:�t+K	E,��;���(#��ݣ���aj��9?�/��꩞\���o(�:S ���N��샒����~�`�w#��D}ϖ�F[�r|�C@��՘�]o�e�ƜU���X�n�<����M;���ᶇ4��H�p����gI\��ќ�}�F�2ce����O�j��o��gM���&�^ph-��)�&N�/��&70�f�Ak+�W+?��ש�]|h����t���ؔ��U6~`�h<� Z�!@������K��%�E���O���qB�R̪T����JJr�g�R��YZ4k	Y����R����#r�,����Ւr,2ϫt�̂��.�����X+��c�n�hU0���~Z	�&Kz�l �L�,�\&�3���R`���~���"��fT�4$.��Ʋ{Y�]x��ءb��3>P��c�ޢ<�.��wO+|�np��k.J�MoW���&�B&lɲ��;�^_�-�!�W�2ەO�z����DO����xO���+X-���ϸ����4l�����B	�)��C��
�O�'�7*8�BƋ���2L,!X��
�U�a�[����%�?t��h�oVZ�3���E}d<P9���2�]An�Ukx���*\c<���	:�tI �c���$��pkP�ou��<��8{B�e����`�`�H�W��'�55�ߊ����eXu]kE8���bO�8��)���ߗ��0k�y�N��D]<7n2��坢yj�/s�A&���e@km����������V��+(u�7�B�B$b.�+�f�{ƱV+���;�����/����
�e�^��\1��
����-u���G����q9��Z# ���݌�z��:T��:<]nby�f���"5�9��'&��e6ɘ,j�ihWcڛ�'y��ޯ��"[�,���� ������}���� �������o-ؔ`6��=Ɍ��/sTS�}g�yr�.f�����w��H��*�U���	���2{����*�u@�g��7�(���Ue��T�
�oV��\xY䧙��P�,-�ń����n�xl�p����&���2>: �>ۻs��� ����p�6 Kn�$g����LQ�-�1H�SJ "�����J���?����c��6s���f���W���%�D�<d�&����QCSa�c�A+)�uW+�C���6<�/�ͷ�.T0 % ���^"��.��!j�X|7�>������Ќ-v��Lj~�&Th���Z�T$�F5�vW L��ݺ� ��ٝZ�o,��w��hN��[<0�߬�F�����u`��}���L�7����~�E�W/�m����X7�?q�S�#ˊ��`a}���{�z&��#W���s�S�}q�;�9g+�X�J�X��]g�9������M��a�tʕ�Ɓ����v� �GZ�7m�0���M�[vn���)�/s�b��ujY�:�A#g�|,�}Н�ʏѩ�&K��Zxa%̬��:�/o�T3w�xb\R�����ɋ�u��`L(C��a-כ7����8��*��r�\�F	��u�#�J��6�y�(��4x�;#Kt�^��-(��РYE*_�^B-�\iit���c�+ރ��D���j�ӵ���P�����߄�XGDa�u������֡�舫�*~uu_|I�����`����A�?itYn�gu @�H����(I�+�$1	\��܌�ی�I���+}��&p�񟂭��t\�o%G��f����% [n�r�"���5i�t�M[�f6�JP���. �#���>r�6��E��eư��5w�hK�O����Fδ$�L�n�Bt����V>7�I�q��)$�3=	����t3�"����+��	�mM�1OH�Vx1��1��횸�]B���z���m�YKڷPP�:M�H���yt�i2�RU��y(�]�d��GB�׮2jD�}`��<��RՕ#f6o6��]�s��k/cZ�m�sx�R4���K�� ۆ8�@e�v�v�k�\�=�/�^��%�e���x3���#�J�ȃ$��V�l19ؤ�1�Ϣ���ijVA�C�<�b+�s$R��>vQ�H"��e�$?��$g�,@�t�7��%7���Zޘ�۩�sΞ�̆�����Z�>�� ��~\;��� 1��9x�x#t�l�iA��P�Y0����L��4����S��Z�����E��b�`TӮF��ւT�ЁK���Z�1HA��{�¹ ��F��l�������9���qC��j���d"�g�q�"�/�]��DY��C�wnj�f�T�f��Ǟ;�嬎�pH��Z~ox�N�G/��N��u���'Q}|�8�����#q�k��V�_8L���_��ەX	aj��C^���Z<<Zd;�~����H�/,/�F� �:�b��	<z|��#BG��I��#w�e���f֐�%2H�[͉�'�Y����m���I~�U�����XvW�ghڤ�f���-�>P�hrW1ݵ�M�eb��������I�b7�H6���r��fm�����wS�|$>>Mz��dP�$i?`���m��BD�R�.�����G���o��?Od�-=@���e���`	�sg��ӼAj�p�f~ȣ>��u8��_V���1ċ��U �jC�e*��׸�=��jz	��U53��(�K���	I<���G����T[.���  u3�,���< 	�	G@Jݎ񎿼��E�,*2=���1E��sq| B�r�RJ=�M��*Q���ˤ��B�����r+�Gp�%?��n�7 $c��n��G,���O���I�s�uj�P����u�ö.�S0v�o�?E׺T��Ug��|�O9�T�Eyf�j�4����/���(h���Q�*��t�6���i�ݐ��x-Z4�~gb�:�#R���y�D�E6wѕj;�K��F��0��-�\�o�����J�^.�����ά)@��ucO�O ��f�]��%
<�m��ŎJ�*��~�ν����
��g�T11���i�$�҄q6�E���$��5�h���Z�ń�t������0��`�->VU�}�@x2�L*���n���)-�C�W�����������6Í���Yn�%�+V�l��yu'	��m����W<9R�H����鎅X�2���Ns�|]`��m���S��؎�Q/�΃3��	��hT����d��n.�a��&i)W5\c�!8�匶�A�1���L�������u]��1��%��r���x#%�5��w2$kP��gȝ��+�}�h>uN{�}�Hh0_��}2z�Ȏ2�v�Iס�,8���_�1~�����K7Gz���I�-��}��	��& XXv��B���Q1�k�ו��l�b��5�{�x�(C��V��5��s%U����o�%��5���w�i�|���8C�	Y8]���Z��a('%q
t�W4h���m�����x���Ou�=8��}�E�xV�M�'2g�8^�XX^ZW�ž;�Ԧ��S��r�<vy�r6<40�����U�)T.X�	Ƞ9`���&=�q�f��t���5�X8ؑ_Ul�l����/���|�����\�yӾ��<E�v��$�n�{t ����wA��:�:�6T�q.X���eO�A�	0H����s8�ء�3��UK�Y.��֓�?�A^ٿ@Q����v���]B+�'��� sڸg$ʜ�4��2��6����;i�z�(-�"Ӣ̭�0����T��~v�4�0�w�u4��9"��E���7L#���\Q�D'K~|�E�rۤ���r�V���0��Ɔ�_u�]�R�Y��)��P�z��1�@���x륶,���ԓ�F~�b�v0��(+�,�Yyn���4��?�X�T"6doM�G�ƹթ�\��|]�D��	��l�E�tZ`M���b��@g�H�&��ܢ^�jz��*ԝ�-6	�Ǎ�n�'��oT��'5����bz-�w�\|��Uk��)V<�f�c��;z��|	"l�v�ʑ�TN���\�@����x�P�@�c��*�7�2�E�-�9R�d҉��Ae 
�(���ϰ�l�k
Gc�X>B�1qlew��o�Lb��c@�O��b�廊#��	*l��8�d>�|��x���p��@j�ь���䕧\ڕ����FV���D�").�v8b����*����,�":�/9��Z(^g��gJ��l}��Px��f�r-a�O�oo��y���b�w9��bò�u�[h0 q;�6z7�`��y���xz_�hn7�H}}�䀮�z>@%�K6	a�JJ���w��a�]�v(4w�M	`��z<�t�d̖�H� � ���pB�7��#��D
q ï����4ll��w|<�У�\0Ã�.��5(����ne�ʴw�l`v�o�}���-D��:�
�Ӿ�-N7`�bC� �.@�Y��m�W���g[��H�l�1�e^Æ��!a��Fw-M}S�)����^�CV�ն��]��Q9�!�����Pm<�Q��4��7U��U��L��ݎ	��f;�� T8���n+��0�D�=AZ i��-�W��ky.3��g��QU�ʴ�IZ�<���~l69�mX��L8ܲ{,\�!٥���R�>�tp�}E��V�V=LD:U�|"8/�(Ol���o;x2�*Rį:�x}я�r�R�F��#�s�k;4,���ej+�*�(�v�	/�o�Fˠ?L�#E�zOߤ��}�¿�e D=�Đ|�&��7�d�����'�a?n�u�҂h�^���+ć�h6 ��'�������p��`���$�L��+Κ�c�����%�	O���x��CX��y���Eĳo���`�տ|4�>�eI^P�I/��W���\�h�#����D/}֩��6�pk�O�����3kS�+45�lX�v̾��vg���[u�F��-c4� %80G!5,�����;4e�28��k���HP��3�ش���_j�����}��|rRm	�K��z���l��"=i���'5u[���%�]]��g3�������WYtǚ��ti�I��Xf�٧���P� C�Ɂ%�V�/������$��;��y�0�@u�p�'�\��!6��Xb�Rd�g��ZK�'0�bܣ�Drصٚ����p:ç1��
�)���(�S�ʳ����A}���1��%Cy;���@h�?\�RΏ��+��%l��
b�{��y�B0_��w���oQ>�%��}�{Z��{@����lpl�7���-RLD����7�A	�:e �bIu���nr���=��^�9e���3������(�R���b����)�'��5�`M�%�Mpgp��k��A<)�w���?���v?Mx�.�[�]X1�?$5P��
�kn��X�u�*O����/�kc[�R���dBn��W�Z0����H����HLj`���0{Y���$��}.�O���m1&d�Y� )� n���k2Bq���Ջ�) |n<�7�B�)D�>~���Q�K�d���ޣ~q���c���Pڢ�����3g�iB[��V��.���-�U��\C��''��N=4%m��$���k�NP���Z�������h�l�:���n@��^�̤��9)��\"
��ڏ��&��B{��x�3�.A����(�s�oz[�7'�o��Ov�ɟ�T^��&W��0�G�a!����v�����"�����r��,�spg#�܆S�LY����.��[��=���{���"և{�3�JPy���Ҭ���O8A��X�]j�AhG�O�ߢ8�f%Q���=.�,SM���t-�P��kh���r�(��ڱ��Q�n�K�s�dv����]��4/�,�����Ӵ����x�ne�Ln/e�f�4f�EeP\��}��r>y��=�ڀm8�M4mQ��A/p������6xS�����}ll܎�`�=Ǟ]�n�{����U��pJ=�â;m'��{��Pp�������&���^�}3: |i���s��"R�L�-:K�I���.��烃�'��;�H�E�s]�D����̆�:%���y��j��oԹ���MH�Olc�.��M�4t�����l(�<�m�x~0���F�} �#k�w�R����aU��@�
rNL�=����%V	�,�Z]bzzE�7�m1�t֖qpᨀ��	]=��� �q�&�\e4���+.�\�Í\�.N��6�p�f}dvZ�A��^c̣�����!���g� E])��9ZK��`�M����)� ���D�ye\��rO����)f	��c/�ɰ�:ɧ���LQ��G(ls#�)��Ɖ�9Y��8����P�&2�,	�VW.����uŢk��Ҧ��D����5�����|Ǡ(T1�HW����z�P=��t�N�yL�墚pׇ\{d:����Q�$��t>ټ�����|�"{���LJ	��ރ8�2��18�2
��K�
���� �R�~�^�(�5��
uIm���Dc)���>k���Kԅj��fO���AV>�ݳ�d��A��_�<�wZ�a��ښ�+*(/o���n��(�
GmR��E�G0o���Ɔؾ�\X-�&v��S{0�+X����6���d����P��چ�6>3���%�$]Ê���z���n�TS����
 x
�v�1�c� l���;�L�����h���t��r����W&�����3���!��E��.m��!�t| ��'n�� �~YG��R�{&#4�K��'mV�o2��3�><�q�*j��	�k%�^~ [']�E�L���Ss�~�k.-��49Ւ��֊���&��*�\��#��J��G�``L	�Ex�����=��>o:�?��b��S���G�=,��'��Gxd�Y]��
�i;�a���� �ufodo"u����h>�;��*sx>r�i��@{f�T]�
 <AoB����,�%��@x���Rm$&!ch�	ћ6x�IB�h��j`\�QF1t4Փ����)�>��ms��P{���Hc�rGv��5}��1s@��]�R>�qH����3�9�@zVԳ��zzB�%gP0m͎B�˵���P��,�J�2�$�[��J����l��?|#�^�8|��ənP?�?�X%%�E�<G
�y'�}�|�S�t�돹��^/�L��'�Y�.�3 �r���rY��M&���X��j57TfʜڛMM�H���>���*�;��U\9�8\��l]�Z:��ඝ˹p?s�C"^��cKg~
#W41u\n~���Խ� �ut���N��5� U'7��J1nN#���� �䲬�ro�>�u!D�&l��ɀ�]g��G$��Oס�"7p����]'/<q��B�	��J,�H8�쭵�\zM�XIq��ղe�ۭԾ	��=K$ W������M�� ��,�Y��GC���_�e���(B���"���;@S#�w�Z@R-L3&�AL����6�r�{��p�C&�U��.�e�Î�R[�%4rGN� 1���(�c!���.��sÊ�1��V�/5tJ�E.��f4O9}�0X�+.c���q��72�B��Z))�+f�B��n��h�ARR�$���݅�.-��'��GҠtQ}�C���0�(tvfR�g�c�'K+G2���nG:Y."����ݫ�ߺ)M4����?^�B��f�����}�-���������[������F*����L��*,���q��7��7��d��x׊��i��>�V�&���&�h���̒t��5� X��s[�Β �%�V�(ylR�w�$�?�*���ܾ����pO ����s��ݡ��?~�ǜ��-�,���+�v�����h93��M��U�2,�N�o�^N֟;���/{Jy'w���vq�A�T��k��:��6�;�9��ڿ@�(�������9j�a�:W���yyn8�̢�H�u��DM]���f|6Ўgla͠,�s8���������C���SH�vO�;ƪغ��p^Mig�(���o_K��"f�{/�`�Q���%��f�9�m@����n���AI���-��٠���U�J&w�Q�k�TROBǰC�i�ER�Pn��Ϻt���lZU�� ���UM���bԆdw��@g
ja�2m�-�ˤ���?d���)Ѹ�^�-vdE+����whF���c�&\y|�|���4!z4�v�W��{P�!�-o��Sq�Bj8"K�T�;��r�~+��z�h��UQ2�	Z]d�_�����_�(_�eF��<3�$�5M����3�q�z}@�*U���wcN��O�=QGf��CW��pv����g�̎^e��s��0JL��Gx{��Qqa:JZ_�h�X�C�ɴ��*d�$�����[�͠�G���Dj	{������Z�Z����EH�՟�O�jܸlv,�B`��a��5�����(r6�8����������o7"A�v�2Hbɶ����хd�^j��8�#�_���c�m��}��(��)����m��z���
&q��͌�GG�͒�$s��V���G�C���
R�:~�×HX^W��uZ��TC,2f��:�Yа׻��8��){��ڮ��9���}��~3:�X�W��ba] Жa���*z3��aA��ǝxVpzN��<8������<�<ZQ�X��'�41�����C�n�5Te�w(��,C�����s�����P&A	��E����e����EGH�"sw���_a��$k�`����?�\ق(�)�V��!�� vg���Xbc3�:.g��	N�C.9�1f�f?�IbiUf@����I��8��`y����Tp卞b�B���$�w�>tl��ߟ��(��G�_�[�)�U�9p��#=f~e�GgXK_���T�{�z5��8FD���i�����r|�.��8B���t�P� 6�[�z5�@���#�z�"90�<aC3�g�,�~��,E������Rھ�T�T��wD��1b��0�����㵁�a!P�G�r˴�!%��`�w�pj����V���Fx��?��,��Ql��M\^���ڹw�ϱ(|��+qc�m����bk�)�������M�=�h�
�E$��=<��hP�Be,���"	۟�Z����h�`�?X��\�r*����,���I��D����3M��#�j��8�z��NC�T�3y�8F��A s'̵��!�8M[��ka���q��a�>�-Hc��?��J��Ɂ�+{)]���$:&𵿦W";�Z:�f!D*jh?26@��L:�'���7���.8�>Bg:�����9���]�0b�҃�T(�cᢳ
-�B%
ѐ�$�5�L���>Jrw�I|Lc��=����I��$�%D\��o'�f�H�X�?{<����� ط�`m�w���j,�C�Sۋ9�)K"�������7 ^�l��+Gp3	+���U� ,�!�M���wa���-w;&�Q��,�nP��X!6>l6�.�C�^B��*1�:��9?VHg� )�Od�j'�TaaȌg�B�tC�%U���4R�e<���-;V�[�`�������LG��v} N�5u�����_�{w���~��V�PU!Ϯ�s��ɲ��o��:L�m����<�bֵ��\�
o���DZ�# X��4ui"�	V���E-u��OɓNT�h}4+��n���{͟� :ܼ���Nv�J}�՗�N�涤 O��ff5`��0IT�/�)�$]�>ս�ٵ�Z[3;F�ժ��^h�'�ldp�=w�u��8����Vπ�tFF�A:=Vz�ԏ�@�j}�+��k0���	�?�}�[�s���;1�.�	�mӽcI]��d�������a�jg�T��(�)�1G�z@�CJwb�W;�H��Q鏒᤟J��S���J&��AMV֞��0΢ѹ�,)?��x��,����x25�Z-]uc2h��!:c�]׋��]�T�fU賡3��62��k�54�A;3m�xL�=fJ�M�*���F�ڀ�o�l~FE�|��ֹL���e]���"�'̔}9��������c-V�2�"A�V�C��5/�x_e"0�1R���l�%��Cs��h#,���j��/��Sŵ��^���)��n�I�`�����2;l��/C=x���C��P�����[X�	Td���r���By�r�J�:�Y`Hí�?�|�P�W�h���� "�������Y�$��@x6`��d��j�-�����~r$�7\�y#B����S�%�6}S)Mk�S)��L���Lw\-����A�wq(��p_~�5A4�������@Z��qth��u��C��koՕ�[(c�S�r���o)B�@�o xw���.��|�K{��P��Lգ�u9�`	J0�m�jSy�GK���π?�<_l�oph���B�;V�%B�͜�ޅ�B��A�4|^0抌�v;,��>g~j�%��>F�H8�^-����]�6����J�<�HO��'m[�rȧ~��u U2���פ��F�9�0	ׯ����*l굣�B�;S��n�%�h�z��Fg��d��,��W��G7�`����H�[}�]_A௅b,>I��@��D 8�n�(��`Y��9��D�^�浺CV"S9��03M-*:�տ�Y�d���>�]�B��Ɉ�X��W!}|�¡��U�u���@�Y�r��Y��B��e�k(������F�5
o�����n��m��C��uS�`�($��R2�c�Z�5���?PkG:|~�G#�LaFE�z�8ELD»�Y��[��
�e�.�����َ�!`�`�)!�W�o'=R�XA���݂1��s"���(��f��ϲ�+V�O��K�� �>
�ں���P|����N���5)��0�+fn� {P��7&�؃�|d�!�p	s�I�l�#HK��Ⱥ�<O�蔅Jmx�� BM�k�o�?Z��By��BE4m�͍�b�g��S,����F��;v�Ի��3��~��:���އ���3S�t�7�?Z��a@ϽH�W�s��Q۝_����ݦ|�w|�4`>Q�x� �
��ҿG(���i�(Lt�eʠ�O������f D�&mm����!���E;���Ax;!X�>��u����>3��q\��C� ��ޭmά�/���KT�h�ɈtN�8��Y���ݔ��)�1���Iht���Ϥ��%����7�@��Wgu��ai��fA�W�`�L�����0W)����2(Ep���F0�2Xdl"4*K;�q}�Y3��}!��q`�}��k�� ����t��~Q��=U��/-��۹�O띠�(���N�	e��b4l��82�
�~����Hq%k�£�"�Xi �y�ڷ]��;��x?N�̵�
X�j����/��n:��YH�	��'�I(��QӉ�
�a��"���$)p��P����K�
�%�<W@|��k��\��/!r�y����î�
��9�&FY#6�Q���I:(k(�>�:�VH"-vAn9�s�x[�� �BiTR�q�K�4�a|w�}"E�}�����Z��u� ��yv����������c��E��	T��������+4iW��~��eR�0 )��*Շʚ��;���(%���p��V�y�P���u���_i�7���q�LK���\;�)��j�N��5O�ǅ��V�*�ш{��i~�*�0���-Z�'������C�-�ND>�B&�զ��L�I�G�=%���0+��򞁆�1c�_�#��oG<���͜?h5��@!x��Hf'Lo5j�M���y�>�P�=H@4i�A/-�R(�։Y�M�g�^!H���*�_�[sG �RmA)��]�]�	}v�x�n�E}�Q�92��ֻ��;��l��T�$>F/i����^�������܀	 -q==#�����e���#v<�`�(��������s��bd�;�ۿsMH�`�r@�(}+
�ƈd���) �! h�J���OiIطX";�Z����c_	q�����׉`�.iϮ���#!Gt.�U����ѪG$)�?��Ġc����H�
��P���=6W�zS��CyS� E2�P(e��P&�Up�z@11מ�'��q1>�Jq4�gP�+w�V�"�~�VF��D��|���<�)PjB�*�*��#���s�6&�� �>���]m��$�
��%�%���x��"k��:�+��ϐ�����
�BRb�?]���{�����Жs�$�
����$���	4d��
�zg��P�5�����H�[%duv����N��{g`8�]�ٟ�7}$Z/��r͞�?��
 �=L�/{6�V�gs�Uc�tU�ڔr@AT(q��R�ٰ�@�S�3�१G��{h}�m��Q��&'S�DK��?�����hޅ<yI_p��jͥ�pz�h�t~��y��I����*2��&����o��P�1?� ��*�
�̪�4"vG��2��FzI�����IU��D�3�R��DY�O�^�/����vL󊉘��z�q#VF#J}�݁�����,�~�d�&q�Y���|l�f�*�f�Z@[�0��}�E�Ff�c\Y��L%�<�*�XI �X
�����^�д�ȋQ���������u��	�w���x�ȵDy�x�1&-~ ��ꃅ-�;:��tcB�B�V5�"�U��])�BU�֖*���������T�%�t�<7��[+fá�Y�k�(��X��S#9�.��]|Jr|�8�O��Vl����.�m��嗸��+�)��E�&ś���h���q��޳�o�����ۣ}!��`�̆	߻�HJ���f�������0-�%�����:��l��a�f
D�I(\�?J�x����O�<��|z�*�������������yBd2�6�I���jO���K�-�Q��O��[?#��M 	e������Biyj����K^R���'�ƶM���ɵ����>
s�42թL��+P�\�]Fcn�NR��$.X������ݮѿ���� J�G� ��	��Vq�J`kxi�O����|��do:�&|E����CB8%H�PA=>���E���	E���PV"�i�Ёǳ��~x�i];�[�l��hTBhQ���9�C�����}�%�;�<�AZPg��I)��8����?��Ke����ZZt��A�}֭w���S�~�1���&���B@k�b�dBQ��^��s&	���׍�d�����
�h�\
`ǝ=���ɸ�o��s&l -�G���$������wk1y�;f�%6&���[��f�4}.E�uͳ�M����1��I���7xXUox�.�SU�p�捯_
����n���xd|�TC0z��zfyۃ�.T���@�����?��O���΅T=��b/4��2
�����aGW+D� �n+���fq� ,p���\)#HX����M~2�I��p��=R��~-�֓�����8c0�?��Ҳl�1��i��L�+|�p��%��\��$ΏBo9�����^`"�Om�<�R�")��uVJ+�	NW��tb��Ќ	��)�nYժS�t�_��o:�<]f�5��S[�<����<��s��c��d ��Ur�5j�N���DV�Ϣ�n� 	���'	H��u`�Mf+�f����"����~�~A�l$�8m��j����� n��k�]5�>�Mb�3�警^\�N��p��6�5.pS�g7nQю��T�EJ@E,���h��I׵�*�˷�u�uu��:��ڝa1�k��?OS;���0��]�3u �3��[��"f�����Em�l�\�0��}[_ȕ2��8����{|�n��n��C�xaa�D�]�)GNt�r�3T̺2���EjM�:&��=ZK�C���٠o=�W8B;��x(y��~�.�-�ЇS�Om��6��!�߫T_�X���=Xޡt�H��#�>rm�hJ\ �Ԗy �V��|��|#�;�]�g��dϳ����'ʕg�sК�^�t�d)	���},P�ͬ���|���%^}�h���4��jM�h�"r:;Q��Ed����')l\�����홍�����o%�*t]Y��Ib^���54]1^�ݚ���A��̨(���R�����
u���Poנ9�,�v�� ����h8:a�=��]�AX	�O��� �K���%w$|~�a�>��Wn�Ϩ۸	�&�o�0��3�&a�磊��I����;t��1��9��M���䣥��,�����Yl��-R���ζ�J���4���	�',�gRl��\�������{p���\�ZD��I>��橙���n�o|�,s#�a�Ҡ���q�d!�]
57��/S�09pQ�1'{�k=L���4Uf�@�6��nH��d�h��Z7>����)Zx�=-`ȭ���������L�oO��y�t�!8A�t��R���	J�5z�?I��
A���>�OиCt��r;�=̠�#h��}��:W�y�pc���c�@�3x�A������n~E<����\��V�*~�y �a��f�K�l��_�@��	�$G��q��A'�T������f�52\�a(��`��ᢡX"=6���m�Ď��_�ڇ�Y�ކC�����8���G\M���Dפ�GI�lp�`��ۦ͓��(�F
2A�$
�A� 2�e*��U�<�ի��ؾ�=;��s]K�l�f����U�p��
�Ї"�A1��v�oV1�Ԛ��0�b7}�
���`p��Ƕ�r�~Rij%^d��;��.��	�Ý�f%�k}
G7��#�]Lk�8ǲo���qT/ �u��K-��7ל���Ґ�ss�l�1V�h�/�R
d��SzH��ч�WV{ ���3Ft��_�,xG��D�E=!�_d�
�j�mL�d\s�b�{��Wl��J����C��3xm���m�lt��	���Fke�����!�"@���B"6������%�����Y���'�5l�^^�գi� ��1[���kƯN'�]�Z)���$�����Y�C�AM���ȃ���@������tK�9	Hǡ��2��e���nE�Fg �PT7�B���4�2:d7j���Y^7��[�K>x�'?���'��6����<�������~CrD/|��~C��y�},��"f�X٪��7/�$*���3�@O�7�������y�O�{#�Qt:�Y��P+���A��T��D�U48_[������(��ro��()9}es&[�3����sq�����E�M%8�ڀG����)���M��7��xi�C��D'��$A�����-���d�:�ݘ6�Z_��6��e�n���)�WU8|U6B���۹��h�ˏ�J�+��O�i�o��ՠ.�.*q[�'�A��:ӨgSr����h��5�?B��6���wvUP���P�ځk�d� p?c���l����`g�/W�<?��s-�Q��G��T?��(c�	�D��RppI�d��2�ۃ`��ѷ�/dݮʩ)�h�.���]���z}���?���{g(Bb�	��(+C�W������Әt��|�qv�@!���~��.��d� :�q����m�n&n٦���{Xa��V�tOm�Z�OR!D�m��b�B����}i�	5��Gc��d4���\S3N��87�9*���h��}FCHϘj����_�Zbߐ�qL���D}�	�T_�ii;��v��V���e���2�������}�0�*�����"���yUT����)J�(/�j�0�}ӻ���w���T�>�pI��s�^ܱ��#ktt�US!]�.�be-����Z��p��؀��> 0C�g�(ć���SI�\0?�s��D����/�򨱵>|�T�~o��|���_(L��:�����.#�d]/ ����*�چ,���j��7(�p<F쀊pr�-?��u�7�s��m�&��T!�6�G76�%5���"ԇ��3ކ��Z*va������4��яt�F=��N���դ$���@�*m�AN�����Q��D���hF��־��4`���Us�.t��f������_����ZN}����r@ǚ���|'����Â��mt +R���]�����R�3�u�«0�ږO�!X�<S8y��6��2�A�@A\�Uכ��H*��H�I`���-���RG����k͘�r8p��|wZ:(�I��][����(��A���� �]h�+�B5˥[�����.�J<��)�A����<�F�3�/��ҳ�d����=�}���<皢S"7n���o�|�xӁ�[{�_�^�ډe�zQ|@M?<L	R��^�v��>_��؎ƣ9&
����LSڳ{��ِ��¿6;�)a�lF1I��F�\�r��'Z���q��#��A=����ӫ�()�D���f�M�KQ�22 ���4�i�C o1�&ۻ�q�3��鸿���DW��3�_&4�����U�0����N/L�ң�v2zq�/�)Ai$�)��}l�U;����N/S�ơ�����.ĸ��ն(N��i��C�<�d�J��Eϱs7�-� 1_78b`���mI����a�|��F\-3�ߥ$Kڞ���**F���T	�!�؝D�2��8��)���$�ɖ2�A�m�B�n؎�����J�+�k����w��D��y8{Wԧ�NA�)Z'��=x��Hj,/�u������V�KD�k~"�@�_�/ dz����)��~뺯e���6X�,�[/�m�y撿4�}*�����p�6�*�Ҏ̡���$�����ܲ��d�^$o�Ը�v�V$ڧm]"��k~d^��2ݧ�o�dQ�f��������.�q`���rG �N��o�/_����]��x<=3/����7�D-y���s���t�)���Tp�`��A�ôC���e宩2k1��0z�.�['Ux�Ď��=�x����p�C�""gK�� ��!xo�4:�d�=�(�A�Z\e�jG���=v�[}����62�8�'�0�����L���k����G��~n��i6�l��v兵[Pވ)~�N�]KR��=a�����l���3�#;�@�eqC;��Z`��[\��U�Ƃt���z�&r���}��9������N0�q���kY7�S�[ ���� ��``�w�9G����du���Ht]���l���VEp�(�&j�3�eQa�Ư��P�l�v���5���r���#�Ա�P�W�R�4l5�Ƭ@ΰ��̅|b��c�0��3���||��v��/��6VLLK��d`�
��9.��H\@I����/^� aTR݉^����]���Gd:P�j��	���H��ǳ�rw�h�t���^�ǝ,��z6x xZE����'#r��Ba�CuKX\�ժD=1e�J|9u(�"����S�J���s�c��:uK��=@���/^k�f�syi�� k$���o�z�3XJ�f�,$'�[5*�r��b�K��Q�Oo��"���H��Oi�vG�Č7M��Y��t:��qa(\&�Y���d遼�Y�#�3s�������##�*��������0�/T%Ɇm-��Y"O q><��_�^�� ���πvVD�k`B�nsE�"�1�S��8tGhR��;6r)6v�/�:�m���3��s.�<,���b�J���`}z�6�F{ܯ�S[yʢ˝�oL���[r
Û}���/����0��g��L�pS��G���}W�(������p$��e�io����t<���eko�r F��6onnؿ���T6��3�<�Mj�V�ثshN��[�V�y������+%
ߧ�a���sR�.s<f�g+f/�t4���	W�̐?���~Vd��ޑb�&i�� �����a��9�ր��S�AQ�%$�"�e�F)��
{�8�re�<��!1�:�S�r.5��\��'K0�Tn���Uy$�={�E��R/�%�������h�{5�͍vo��}CË����oGk��[���X!�9�����̓�bN�m��ND뼕�
t}M_��"W�5I#�D�{��rT��7��0�#Z����^�2}~�3a�L��e��0�Щ�H�Z�5 1K��ؠA�� ��B���O�}���O�K7��f�S� �nb���v�Yx����Z:�j�Su@ӑr��ui�ӌ$�&4��a�2&wilQ��9s�^!k/jデG��[�Cֳw�5�찷�������=�p@0�ά�g�牐Ba�a�P�r���0��c����Ύ�-q�P�d��Vʟ�[�~���s��*� ��kjb�$N���u5w�w�[4_u�CRla����>�*uq4����y�%��
lffk��v�ԑ�l���#�����i��;��x`�]
oo��7O)��љ���vG5�Lq�\�нS;@����'�.p����nm��؇p2Ui�Ʉq�[����n��&(���D��w@f�S�7��K�J=~�]RB�Z�J���5 {[� )��k�V��f�*M��^4���\௟��^(�=�o5�Ha���ھ��s�A��g#X30Y�yV�3
��$�!��ZOc��h�}��a\���6��εa]bJ��ev"�k��X�=pfT�WY1�jOX7�@&��G�0�
���>��������J-E���1�eg�,Z/羇&N˹1C��J��m�M��m���[�ɼ�q���=����?��&Ͷ����-���&Φ���%�u�Ai��^���*���SZ�IDt�g%�m8f5����&��"�^�d+�Ͱ��V�MܽX�˺� T���/�:X-7�_ ����t^��f1�n|�Qov|��w+�.GV������HSH��N���j��Be����Bs���'��
t��K�6����S��J�c�'ˮ t6&��"�gZw�S�Z�#o&p�@����0U�{Y3������Հ.�rB@�($G�@xhF�?~��I��L�9~��b���*��֑�@T�g��W[@ C�&�N��|G�R�(v�K��^����fx��N��ާ�2Zq��s��c��1N(���$
��-dt�h�Q�m�؃)���ж(�|%�?�dW�̣��WW�ݤ�H��w"'/;�*Z�EvW��Q���ЫFfrO��&w��d��	�"�~0�9��Gw��ؽn��ȣ	��.,�ܲY뷜ؼ�M��L��6��	(ɱ�GIVXH�b�s;��`M%�5����{c�v��/�Q��w�nǮ�c�zf;pH������9��q�,��/�X5���n�N����o�ɔ��D�)�9nKe-�Ey�1���VUg����2hfhGJ�U|�!;�C�8v�<��L�����:*�E%�ʫ�j�p=�÷�iHt��4�Y��SP�h��p������q��&�v��O�4ɳ��P4}�m:�=|$'%�9�����N��z�gv����t��g��`��6�ZM,�lB�ƷwH�<|Kd��P���iF��d�/8���U�g��f��U���?�O���P�F%Qo��Nՙ1���'b�\�=��:j�	�Q��L����d��r�iGE���cű�K��l�� �D�*z)�s��:��bS�G��Q��f[�V��!a�I�������zp��cK����������5�Oz�Q�F�x�X�J��;�Ē�h��(t�/����<�/�>õԞ3/^	��)E^�&��I��|�� ?�9�0M|Aڅ�C�Z��e������YY�j(DE^pP�${^u�G��P��Gw�;W��?�~L��{��ZAFPz��j��h����ҏq�YGؙ*����Xi�K�h�"�B��܋4���LN=�*/��{����/jS8�q�+.	���c;�����,��N�E�LBWm��j��W$6R���8/VK���$�$�c����\�q��p�9V߫M�z��	 �C���u=Zu?"�r��r�`�X֮�ם�[��fV2���[ `�b�J:��#I�۸�H6:rG�&�.�j�B�82���X��W�5s�r��a�3���H�˴Q~�S�������kS��S�3��ת9�ĀK���c�<&�h/.R�K�I����PC�T1�L~�;6�)�`7v؍�O��p��x�p''����>���6:	>t��پ����~�d ko��(���<�Ը�N}S:ւYGZ�����F:>�)~8.a@G��@��e֟�F�I+2�U|�����/���� C��J��c:V,!﹅�SGD�<�X�tD�w���9٦Z��V�Gp��}ʕ�<�C@�-�6zz�,�/h#4���yM�z�2��&���\��t�"�]Ay������:�D ��fk
S����9�y�̈́��r)�r�xj��lQZ��9�]�_�W�G�&��Ь��� w�C��S�\ic �c�� f��Q<��"{	(�0'����:wi�x�ӻ*78���PY�fW'܄���*l5���F�0E&�e��x�A����r��w��M�TV��c/�%����.��*�I��Z�6n��[Ƨ��wg�9K5N���+� �HSc�J���Լ^pREM�x� B`J�[�� �1��{R���ҹ
��H��mM���o�暉��V�5nT{y�%5T^V��g��M
����܁���x�� ��h�j���0)4�-O����4���3}v�҃n�k�O6>�KQDz�M�A(%��0q��J]����)/Z��Q1�ZK5�����?��;�,�Z�=�4�]UD��(����
ȏ32#��=_2�X�Z\B��~ ޑ����U�{�4c[f?���r�O����ʳ)@��y�L~#2MR�1����ί�ʕ�yWR,�mJ��m��t��h��grb�����?��������TwAm~ �86չ��O�9Nd:`��rO��u>-q�V�l
u��hf��3��u��w�p�L;|�Y"��-���a�����.�R����6z��Ө��&�l��MR�;�+������T��~�D4��O��y�2�"��`��/Ȣ��]	�m!%y��9�<����"�C;j�$�e�x3�]���c!���t(���K��e�,A�c�k�B��&������;�J�
�JL� ��mL� �kfi�j��ǒ��_�r`��B������3�U�����'Ԗ�P����D\��F)`�VU�֌��r �]<�9�{cC{��x�9Z{�����і���d�֮��.��n}~�$
��X\�*���ƃ�;���".���C{�y�L�ѽ��hf��X��a
	-uJ�G��Fm�SW��������ݒ@�H��E�R�1N6G[Է�r���\�*Ǯ���շO�����o�[	n�)8��J/^���Ɋ:�1�Ps�f�3���@�A?��[��ՇWp&�T��{�Eꌞ'�
���F�b���\3]����ÿV۲W΂��x,˼9j�˳�3�}<𙐮�sN fCrPkf�@t��;���k�aV������5��
ٻ��[psw+O��C �6�����{M>W��i���z��v1�hj�O1�"�+�sge�w�г0u��|�o\�CW!e��a��s��	2��l1�A~�Lc%��68���[�]��s[
-�gڠ�-��]�|ڗ�r0ޱ,OLF�-7�{��2C0Ӫ|���,��ݬV"�k�;���N2��abGF��,�5���]�)��U��;�Wj3��v��02=�>��e͊����t��Q�E�]6e�VH+���R��d��D5[�]�T�d'r��?����4s�=]ﺻn7f25s�j��|F
�KC�����qa=��b���qM����sK�/���c�i�x'c���z8���E�4��D���͘HL�n��e�\���:M���Y2ռ�U� �˝�B������b�E�`Z��Wy��Z}����:��a�h���y��֙#Pf�¬N \'���N#k��&X呹�f.�B�)�SHt »�#ߤ�[�h�UqE���������K�_�[�L��Ï����c_C�h/ ��h�v̾���-������F�oo��=�FhE�����������	�AF~N~���O�\�{���Rк2�4��dM��qZ�����$�ٙ&5��Ҧ�!��+�:,o�����RDAki)�$��كӐC����w�i�.x؂�\�۴bdK|z9
G�.��z�,�9�}R�桸Y~������8�Wq�(�o=�A=Q�o�pZ*�\ȟ�Zڣ�eK�@!�墹�m��F�5f�N�����av�x�g�G>���B��K�9CA��Y5Ѭh�q&O��{��YtQ0�"!*�$�����[*�W����2���"H!�ı�����Z���,ҋ�?*)�	:t��/$ioʋI0�z���f)�`��aWYC��O���a`�G"T�2q����K����"���>f�8�ďm@��
^����Dd��|�A*�x���� E]��UQ�A���������`&�˕��u�
�j���ͦ�+��C/ ���ƾ�*-Đ9li�X8����S��01�?l���7䠯�xuӫ��;q�2aCw��G�/=�g:1�ʯ�&�b}�h�c�O�cKƫ�w'��5��5��X	Ex�P[�v�$u1"
��L��-j��W��j��!8h���ɛ{t-:r��xd-�#-�p�ܔ.����:ǂ*>8�3�&m�
�����ͼ�������ݳ�a�9N�fP/r��ʿΧU�B��B�4�����IzE���Fy�ܲ��~*@7lU��黛�i$4�]�9�,�tc"�F��M����B���b�Qu	���w3$�Y�jL
�h�E�������2i}� �ǭ�\\Y� 7z,�Tu�\/o͓�z2 NL=��M$>@���n��'ל�Π��ʴ���I���>��U#�^���&S)�>i�㲘EWoI��o;�ZA
N�wyxd_E�z�$�dR��Ň:����h�x��T�M`o,��-��M;���=>�j�o�����\�?ѥ;�(�h�$M�HӵuF�t��[��?%d�b��'+��]�;�5  ��|��_�O�>;�Y�P!�U��o n���Ù*>_���w��ZS�Db�L0���c�7�\R�Ң΋�|��1G�������;-+�H���S����jn6�=F����SSH��g�x�KR܍�H�1���,�Q�D�m���gɅ��1�?l;�Cw�=�j��1�ju�2q	�K,��W����-�DL�@ʀ��
'u��Yv�(8�7=��R)��'��dE`䜴W{�3lB��ZJ���q4�.�7U�I^uȘ�W)rbk�����[i�RnE��!�.�Zf��\ݚ�P�U�M�h�a���Y���|A���v�}����t�o�;�ԇ�P�xY��b�yg$�-8�^Ä�K����d������*U2�l. ��+��/[0 �m`�"���6�>
s�@dD�l�8�+u:�РG�m�uN��g���Bc<�)�
4D�$��b� p>Hi�pj��I�!� �-�}��C���WZh��1��R�CuY'�D�,���z���r1��P��kɼ�(� ��8L���8��Q����5�F���_B��4���~����t	EA�,UY���,�8�b cX��$c9	�j@�{�Vϛ��#��b�i;/�'@L%�M�<Q�����,\�H��5{�;}�'Q�������LH�Y\�����{j7�e�K��#��n;�>�Z���.��,�m���+$�b��`��R?Qp��\��l�r�^Lx��zn`f$�h���&~�8*����AD�#X7���|Tc�#���T,�n�b��Y���s��;���Z+�W%��XJ��i���P�=/�͗?'SbE[$"������6���*�yv�|��f�� ⅒ ^wȜL~��rB/�����y�w`������!��C�_R��W�\Ҹ�y�K+;���}� ��ls=��2�I���"�tOw������%#�N��8�O���v��CA�w�r�B�]�zO��p�7f-b���:FWI��A%D������B�zw�p��06|9�q���i���k�ʴ&zK�7hD �L'�:����^��H��\,�z��%������X�Nw(A��=�[23��9'���0m���8j���� ��>�|H���	ص��+�3��'�t��}��E.fuX�?���^��;�uM�u���]�������$ru���9�"�I��7���/���N���?}ʈ�=��aLdG(q}ހ��Ŭs�BxS6�ǅ;jt�@=�ڹ��J��	�*�=�I!PM9��V�
�4ܸ��C��"��ѰJمt���ص�G��I�l���� X[�E鑟�Vj�	c����.߻����562߰m�*�т�Tp��7uX��;}��qZ�b��
ƏU7���>�t��BǮ�/xH�qbY�F��z�PB���
�\fS�x�q��ޤ��o��j����O�c1b�Τ6=9㇁���bK Ѯc�k,��s���MR�F�1�~���	���q� ����P淎O���������3�q��[zt��?�I��`E�$�]a�����|�b�2�v�.9T[�DGU��`�G'�&��`M�y[���	I�B�i�0�Ҽ�����`G�hk����.}dV�Bn��p��K�t/���)�9򷑳X/�,t����-�{���K>�o R�j��+���
a��]�U5�C;���s̈́7qtph ���fz{��n*�����fJ�Xp�f����f���w�~(��L&4�lq̥�W0��~��}D�p�8^M�Њ�xj�����
��6:���,�ê��%�A���F!R:����f��U��D���3���.��������_��N�L߷�-�=�M�#*R���e.�u���zC�8' !=�Ф��xV>4�6�l��{�Mn��4q)�c��e��Ȧ*���"0��.��Ϙ���b����ȓ$)h'�)�YN�߮G�`��m�V�16�� �s�������d�7�r�2��])r�S�9���j���*��KU����x�8WV�ly��|c].|B�ld��u�Ak'Xu�8l�a�uh�	 �}!�iu0��j���b���O��i��R�9nCb0�<CZk]�X�L���a����2d�t2���4$A7�]	��si �K�@�BCY6Zg{�2H�^�6�G�`x��v�tE�"v�.�,�n��9���ţ���YJ�z/�K���� �+�:\$�pOdj��-I�!�s��\���i
nSK��h��LͥQe�P���\rh`,�;^19��!zN�cŭ�Ws �C��ܺc�aR}��p�w����ח~�+��ZK�o���u�5���Dw?T�:�ᵷ�Xƶ�4<���t�;33^�VF�����sXt�a�1��f�G��_! ��V:�	ohkP�w��wQ��������`�\$���jg5d���@���}�پ5�H_(�]B�\�#��r�|׻B�.?�.���ORwj��\�M���W��_AL1�*:rZ �@+��ύz���J��Q2؃I4��?5��_1��fsun	+
JA��<�4K�a��=�Y6�<��z�Έ�gVj��j�w<�Ə|o9]�4��k|��̐��d;�����ܰ�aЇ����ֶQ�q�?<�ʊQ����u�We  w�UT�<��V鱶����q��vDi��*j:��H���١7\̠$A�+��\~4�����v�=}�cHtk2�T�w3���z�s<X�&Ea�o4��G�V�Z0\ڶ�y�̴�a�hQ;��}3*DY.p^j̲m�O=D�l�I �<�s�� �a/g��u�@��� _���S$1�R���}e��=��m����DP��r���-9z���t{I9����evy^?�������P^�6�!�3���Mפ;<qG%�M�ʊ����h��[A
��p/�7�<�е����E>��}��Um�e
hu�\�H
`�ͱ�AM!u�0@%���u頕���4�G�B�d��l{���b���<����x��S�@����ަ��@}a�/UI�o V�\à�dW�7b{��`��'�ZW��0 ?n�L'��v�L1� �[UOo��IE�����yq�z^yX���<t����)�[��&aC�GU�G�|0�"�Z̊�f\�S�F�b�c�+���la�rh�w��qKT������g��*�����5�:�<�d��W�.�C���=_�:J�ٓ��"�U�ӭ�(L78[;]W^h"��8�<j	�@5
z3G�aĭ~/<����h~�_5���\�$�@9K��N	S�գȢ6����&O���U���'y�`k[?����+�i���Q�-����lp�~��L�})ޝo5(�t��˄��_���0�Z�}+,Q�Խ�v�]뫅\�����_��A�$�l$ ��Wq&��9��I�&�]c���ѣ�j��������lJ4|;h:���}9�q���6�`f^'Q�B�ڣ���/��kUщF5 Ą�����%2k��;��|�����[�̓]��7�}��9jyI��TM�5	��J�b�n6P�Y�pK����
ݳ��y����ǡr��`��,J�$Wni����vo��5�L%SX��s����U��Q���z�P�к]�N�dF���MN�?�娧sVT���Ox�HR��a��Ĵ�]�v�nS
���^���7�[E��wE_��<�<֞�� C�\5��C��t[֟fO��!H���iO�sfb��$i6Ψ.��'���#�CZ�s�7ӞA�:ʭ� u\I-�eM��R��o�+�m����ڄ�氁�Ӹ�
$�`�ӻ���~<����D!��g`�������P"��;f�߬t��}�'��j�jr�����`=�q
	߻ k\�FB^Z��R�<�Êj�;�ٲP� �Ýg�P�Np����w�o�T����Pt�P�!�!��&���G��G�0)0s�w^��7�9�}���:�\��g3#q2��R^6σ���Q�$�
y!��BG��[�xP�9pti�ѣKJH��O,}�b�2��q���B���!�H�Ma6]:4�Z�qSD�=2��u����&�:F��3]�y��Z\u`D�T�]���=~ϟM��vi#u��������t<v��~�r},k��ʭ�)��k���>$��c�n{�	ä�)�I"M�2� �=��#��q|3�G�3�7i�3/i��3�f�;G������"Ot�Z�օA� i3ж��n��e��~ӵ�-�ѮY2K�x�� h�,R~�����Ӌ��C�}S�y
$�&�@��5��sۖ���(��s�)���L�d�c�r���E#��@�D�����!�i|�#a�x?X�W�$��"�5�����koZ�h%��>s���\�.D+����6��������
yb�g�v����@Ч;��f��Jc/��wȿv	q5�/2�6}�������K!v�!��pnY���R������������68�u��E��)㧓�%�:�8���oB]�.7�����T(��������xw<n��Ǟ� �����<���Q?�=ڛ��1	�j"'����|#�cvC-aHK��#b�,�K�ag���n5"�|���l�"~��8QP~�x�1y@��3ܱ;ch�I��W2Yh��3���:i����� k����T�p�K�!��͑�b�0��-��r��X�������~��r��J\�㜛�����¤��2�,����S$�(�'��T3UO�%�p���>�d+sOV%5�6��I��h�����J|�-5�7�x؝~C�`��s���*�x�N���%����h1p]�=�_�|�;n���'2%�z�8Yb;�K��Ҭ+if��&��E$�3�ig�N�hR�5�-X	x_A��|�9�0rL���H(P�"5�F�T�t����p��p�d���my�Z�)�����Ue�5��h��=c�-T�8�\���]9Gn'�ŅH��S%:�֊6���t�2�u�rB2�<_��)b�ۀ�I%�*Lx�"V8X!f8\�u���-�֜2x@�'�u��)�r�|&�Xz��UTV7�̦��g3�f�M�0��$R���*����m�!��)d�b��H�#����6w��9�v��N��bXOM	w�{���X'�]��{VM�]�J�8[�5
����"�h��}n �N�LMG�b{�&�F���t]n���7�ּ_��ƕZ9���\�PҤ%'u�.����kS+N���G��7d��I>w9쀉�E[�{�����Q/͡+89�ԥEI���k��nkqa����6��Mn�D$A5=���_j~�	�:��e��<Z���׺�3iv���ы����g5;0��� _�?��s0�����!��UW��$�&����'mr��}�L+
D��T�3ˎ�t��?�&���~�H	h�>5B����n~���>t�䴝���z�娓�`����k��ڊ��/�ЈRt�� �U��n|6��n׆�$l���Y~�ެ�J�	�H,�����6�ߦ���o=� ؼ��{]�m!�W���Ѣ�[�[۟n�������Ht�:�����*���r�;�4��+�!\@�,��}ץ=��3ovI�f�61���L�����4u�$D�fǺ�\��Hkz�����{�F%�[���f�Xܙ}'�3��@X��\�U5��΋C���_�R��uQ�.Ë�1f��?}�y�K_i�@e���-�x��?�̞ u���!���#yȔ��E�u��/�k���k�����3Ї�еr�w�k��+Dx��-�F��ߌ8�R�aӤ7�鑼A�Z(4��ׂk,f��j�AǴ5��^��N�
�n�*lk�
H�7p{'x��p?�ӂ\�FD�������v�z���Ox��p��}�4}4h��^�R���X�ƣ� �Ir�3o}��Rc� s�WG��0�p��¹�7��P������D����>�{[��E��d��� tOQ ��C�3I��v~߆���'Eཫ�u�g�g�@<��pzD�����*�}vy]'�<����z�\.\X�
�Ъ�_l�sٰU[�s�-$��V�'Y���o%fuRR)�i���]�Q90K�̮����hgeYS��ݟ�r�	6g"�X�x��Nz[V�k�G�Ef
W֏��i�>�N�PºF~X?�*.ثa3�M�[�?	��d5ŚF'<S'��;	Fң�>�7�ݾfo��s+��7
��S߅�+U�h6&G����������D��	�X\���j�9��s�<͂�C �L�`��%�L�K��!Y0�<a�!���5��m�)��oB`�&��S��ȸ�ǖS��y�F�~`\[5!�סp��ۓ����
;=�`�gT	2���ZL�������W-g���v�n:����yq�n����0����R�qf�3��=��I�<n��޵���S����S����<ņ�"���y��mJ}�-н�� m(5�����|�o��T�7���{v��A|��)�i
�2��,:��\,)�Vkw�z +�ւ��R�m6�w5� =����,���_Ȱ�p�O���<J#x�_T��.�f��Rn�bVm��_Ai��{p����{�F�1��O���	�*+?�����,�ֶ	ʨ�<��a�y�����S!�L�Uٜ��'D��}�$��I6:9w��a��r��P+9g��y9[�݋"�G�КuMa�s��ԲU?�&�%
�:D�[�r�ٽ^-k���^J���<�sCg�Ób�ys[._�/��Gڹ(�Cڹ`ύA��-3��)�F�w�����m�^u]�~�2�+8��#����:����u>Y�^C�i���z��"DTa�/��m���+ƒ��xXB�G�v)��¦v��=r�~s� EZ⪟��׮B!�ʧC��>�bv��S _�=L��l�<��L(J�9�3�{H���b\�������T�>��I���`�3iOG�Jc��A�_+f$XW��Ճʀg�j;�G��T�/8�4'�����Q6�SR%�Q��L}���,[�e�^|�+=^|�,N��A7+�#�Ty����N�鮴>��Kf�ր�|�r���(��/�jϟ rD&����u��v��@��;G�
g�h�f�����z��e�j�L���J�o�H�s�' �7�-YN�쉄;�_t	�[ʛW�Fg��qS�����DalOmC�$�u�mw��&�V\���G z;r��,��~U[��7x;C-�o�-� ,��݌�q'�.w�����>SU�ݯw�gM�D%�������{_�y�L����,1dN��v�᠈��VN3��@I	�����|&B=���ܱj�(�O�d#�^F�6S�`����֚[d��-�eg���A�<#�Q��!<��ְ�%��(`�R�)ζ�bռ+�{��'��� ���*-��YO��>����v_`-��4K̰����"�n� ��_�H���=y�js��!��N�����a�BGl�QȐ�׀7-� �ʮo8�f�G��E�)���ȁg@��D�j� 02�Q�%�,y��ڳ:�:���)
��|ɾ�x��
ܜ$u��n0�!��������}Eg�s��(����3��p�%��/-,7��e1��ZW���u��-����g��`Չ�|��6x����fJ���S�\���e������d�%�@u��S�2�t����|;��L��qrZ\��@���C5iܤ��I�K�Rez��h�]?�E��_�r���d�%�?�ڈU�W���j��^�ֱ�@�#V�ͣ�2xhIQ,%[򉑞:�0ĵ���Y����B{{�&mZ�Rӽ��Qj����������.n-�4�$�TҌ���L#>LA,��bҚ����~�J�Kv�����C�����Zu v��GO���S�	�T�?��@��X��I�l�29!-u�iK6�>�:D���^+u�9%�	�~$���e�븪��	�;��\���kU�Jٲ�����P�N��Aƶ<�ik<�F ݮĻ�I����Lk���P]�c�v��7gW�sl���yt4���w>lp���J�Nn��y��z�6�,@��Y��	� )z:��544�IE����?��j�l,��GC�Q�����B{�Y�챹�F?ܳl6yC�(��S��+�ud��NDت{+��)�i=�(�
̔�g}0��U]��NH.��{��FAz�9��N�P��c�r=�Zr���|�N�z��`�E`�I��A,` ?�ʁ~�K)���p�x�m�j�A���F�P Ǌ���+�����OZa x�a�'�,�7�,�+�Y�_2ui~ ��y5�v�j95��`��W��,)Z�9Hd;9��Q�R�N{��yF	�=l�77{�cA�s~�a�wi7����z��o��X[�X �G�G�G�v�e��;����|Lҷ���rG���)��hE8�������Ԗ5��a�q^|��Ԭ܏��X���l��}�]Wg���垬�kxd�+N %n@:��l��"B�1%�%��t	���>���{֏�y
�Z�{�����g7�'k��L�lFrP���s̥�=�+��fB�eO�6���5�B�x7qH$�'���4e�n?�r�%���?Ӕ�n���T��OQ|9+?��q�d*��}ψ��=������Q���)}Q,�ku%$��߹����o�	xg������ɛ~�`R�1��j�+��́)o�J�����/�J�����ꜩ����(�Q@\X�;��5�[�5`����T/>�j�uڶV_��|�z:�ǎ��D��tђ�A�sZ}#�?��t��Bd�]�t�|��܎�58�K����>��u����qf1M�ض</�tc�D3@��$P���OA.εfo�k�i���k3a�ZnR�<��)5�pu%V�G��D�=w�R�o�-��0P���b\&��Z߰�>��O�k/e�+�K���L����.L���m��� ����4���ɥ��Z�XVK�^��lH����?^�e�\�A��#�l1�ƲI����\f���i]0M�����������#����آ겖_*s>���C�@4	"Uo^$�M*!Ȟ�p�� ����j�
�VA�B���������˖��z��H��;N�{7��R��$ᘯj�/o�Ƭ+,�7\�6B��]���9��U+?�	�8��U�X8�R�>�����O�� 2«���|�9Q���Ca~�B���ؘ7�u��u\���c@�����ul�=W�(�O�3�r�;V�M�<���8'�k��V�0f��\�@�憈����Hyx�$�Պ�|����(`o���_1�eP� @tK]$���|\�#%/,?i^;���;5�b�+Wi�⾈�hu�bA;�*�����4D�*�ա ���*)�+R�.nN�z
%a���^*J*�:}��5��c�s}��w�u�CT�����'�LG_u9T�e�u#:E��؅�
�d8?)�Σ΅>Ё��\�="�&tNy�הfNbc�]&��k�>�h��-�kP�J�Q����}fSW�(��M�r#ȴ�TTZaJp��(�˝�������nb�~�n"�Y���x�/4������� �|��$Fc"��)A.,�q�_��K:$;�N,��S��:�R�M����'mp�
�C�v�yPќ8%����G�m�������*?�q�w��F�N��I�'��a�e�zg�9N&���`���/���	�wRC%����;6]fR��W�_�G�
j8���=�*͟F�SR3��ٻN�eH�G�LM'r�fي	k]�*G����5Vb�Z���ٹz(G����y�Z�3��g囡��"��A�
Z��c�`���w�=o����ƥ�.�W�ܧ*ٗ�d"~���
��6'T���9�4/k�;���/�����"`��$����Ж /��
�%z��0�cW�����A�o�`򍓤&��5܏�	��f����sʶ>��Tk�Z:+��T����8��P��gC9Y�AG�䮃0L���r���~"ԉ�O^b�!�!�J��h�޴	�^�G~�E�cjB��)=М68��/�r�-��'�]�v/�U���:���d�]�焐$�&�
L����.e�Ӥ||/U�=)��x��ղ�)����t��&̍�W�9)$���{4�|���pU� �e懫#�v �i`ȉ�]��PXHڂ�ӡrQ��T::�!J��jR$�ҁ�Z�"f�"���&�"�
(yFwRO8�6�Gd�=˛�~�[1����)��5�-���2�"�ͺ�T�E5���G�i���:]��)��u]|�M�}a|�&`�`�ř3�����|מ�)��Eې}��Z=�	t�� �2r�Bs����o��E�Rw<��>n� �F��k_0gB�+�c\�˹�iL�p`z�:%l1�0������J�!=q3�:�7a����?j<�����s=@#B�P�ց:%�[݊�OE���qHb1;ҴmI�XC���VINipj�j�<Y/8L��'�z}?������~7������]�Ѩw!7��r/�?#�ȨWZcTLŦ'+�93���_,i�E5�/���nb��^#b���׬X��,q$)}g�3�G�.�!o��3Ox��3��09����\b���dfj��d㘀���	5T�m���WA\ll���F�F����?>{E�\��̬���KB}�qL����ѩQ���r�? �%��H�q�6]�� �6�7�Fy�����Y�m�P�.��\�%�j�y,�$�#ְ���3k���3���|4����x��Rw��t����W�bX�^�h��W��ῦ���h�/��ƀ6 y�bkU�i��i�i���ZzX5����N�b0����M$SZ�H�����;ɪ�2��� ��c�O'!�2�_��)�)��z�+f���m����������D�<�C�@Ǜ֒��4�>i8/��;(��K�I���պ-|���eFuH��z��cm����3�
D[zˡ��>�Tqr����x#=�i���nz�ъ��̞l�8�����7v��~���Z�ۯz�6�D	u�罙�W��9�`}Z|r!Id+��Uw虷��O�h+���*L��я�H�b�h�M	��{��M�g���*?C��'tN�kd1¼ƅt�u��A�lNS�y%�zr/��)�=�}����VYr7�Gw�N����}�o�����&��Q���'�0�Z����=� �g"��x�@fEMy����מ��,�jbk�w�?si%v{�[G���«��@5ɫ�Ŷv�s�Sp���Шmi%���5Ss�<W�$R�4A4���S!��(���QVg�0R8��}כ��(y H�t��;�wo�O�
J���	~�<^�������Y&�g��A�b�������}�hۭ:/sXX�v�s��V��[�X5�;�|���c;�*�%��C~�ݟ�H�j��nJ��ˈ����ҥ��Y�R]�$�j��s�P% gi�&�9T�)a��3�;ڛ-Ab�c�׮X�(,�� 
������C�4|�ƛ���*BЏoJ�����7�wb���5#��"��@�Ih�M���{�j�&+Hl�Š������H$�\��b9��.ʓ�6잓7��t��!H#�6��{�^�|��\wG>缾�E�m��7���C�6�����U����	�/Ap�>D�e��)CT���pܽ�d�׻�;+���'�N(��,�M����<4%O%TԇS�g���2|r� �N��}�_�\\~潢H�ܦ�cn�P�i4D&y��z�6��-�Ⳁ��/��m� (-���Xޑ��Eɕ����H��������L:���[�f$��������1���+:~7�s��P�@�N��[Vo �����)_A�}O;L���[�������K���?��8�Ç6��E�/;W��X2���чr������.P)ӆF\^����Cj�^5z��'-ѷAf��$��/!MH��=q&��;�>eZ�g�Go`��}З�p�K≏���u�ڴ�ڥ�m�����R���b�W�uÄE�$4���o�F�q^�[�lu�V���Wd��4 �Ƒ]AZ]�̿�W��g�Ő/w �j��6���fW2`����h�O1>���I�.��0�ʵ>�d�-t��i8b�����;�L�����U�����@�	C|`����3���R�ݣ����\�Z\��Vc
����� -����C;���D�s��_���w�V��7�g�濱t�^h��E�&V�U�}6'bb�g�]6 ���M9^榥f��QZZ���J�����#�l�Д�ʚ7ǲ�$�5G�"��y�����8*yz�M�M0�5�h��ќD�q ����^���k^N�\�z�%V�ψU�܃%,Z>G%;����5��z�^�۰�T	\͂
�eJs*�����μ�Q�f��ݕ���E�	)�\ӰNA��h��TLV��Z�20Ǫ�8J��a��ȅɚ�������e������<]�5)`���j�T��|32��:��7RK��t���`o�c5Q���/�Q��Li�n�P�A����Oc�8B���H]E-����S�\4�9Mk�h��I!I嫠+0r�E�#�_M���t*��������p���'{F�F�����NKF-���k����hM��A9iz�p|�N-{���4-!2�A-�:3�b�-1 YQ�f,l��KG3@]����S�=�\���遱oY��ٴFM�u���/u'd�,�H�@97�YjZ&e�&�[�|���:���o�δ��ԃ6�װ@SY�����t�	ԫ;To+(tܶ~Ak�e̈�EJ���o�5��������e���Y��U��N�*�vȱ��y�]�Cz;�t��z��TdҘ�ƕ�9�v'w���l�U�.*�Ѯ��ʚ|>��8�%G'R'��2�z]$��u�_y~��[�\�ӻ"$D�?)�(�fTP�7{�O<ow�T�����| �$�f�C�g9�e�e��^̨H�� �7�����A�gte���;��%@`i�z!T
	aF{j1��^���p�q�{���r3ɮ�L��T	�����[9,%�Z5�m�W�����0�t�����_���r�L5�7�kq��b~I��qνN��Uii5ݷ�����@�}��{B�����7ݝ�| �R�����D��Ys�L�T�PY��?{�$z��=�׿�O)�L/�]^�I�[�����X����כ���䋌����Pxv5�p�IΊߌV�x=R�(`ƥ3m�NE&	�Y~������;O��2�4�9����t��~yFf6V1|�zPۭ�	����VO�3��/W�H�۷ꇗ��h�gb�������6(f?'���7mkX�`�_9�������Ce�Θ�)��ºNO:������~����{Zڐ覎A�/��m��'Ô~���<(��IP�E*���2M;-S�aăl���C�P�.�p��9�	|��I1��h`��� ���	�0�Jl��#oa ��u^�擧��H=4���z�#/�q2G�iv$ɸ�p���B�Gӏ9\��������ɕ��Yv� mf��,�a���H�__#zjy [�)�8r��H�D�E�����E�t��`�y�A���b�y��6��$=�)���q�V+Ϭ��Io���w���z�_�)�7P��&�U2%�Ǿ�1Y�;��_^��<�ͬHrd����y�lJ�:"�y��Û�%��R�ˏ�G=��?$����Up�[%�2�դ]X��Ǎ9��:��˞�2L{ ��G�W��N6�7rF���œh����¤��1z(Q��م�W��� H������S�����Q�GB�ډ��]ߧ���+Mx�Oh+-�x��Ÿ�0���K*�$Qt��x^���}]�(��?�䍲[�F��������Y/u�HL�e�*�P�Q�f���iI	a{�|i�\)�G����M�R��	&�f��\��6Z�� ����ps��:��D��l��/���y����H/���*�|Q?�ͦ �)?�{��K	h��,�j���s�o�S��k¸t|W��ZN�ư�̲���wp�m^r��nX5,s������lyL�{�O��i��!�Q��^ۆ��,�F�-���o��:s!8��J�W]�����҄Tre͂i�]�kl)w�@d1�rjM��~i��{yQ�V.���o����i���f���8c�ޅ��P+��?C3! j>f���ě�J��IW~/}�q���[o"��]���'�78�`����7P�Q�lp`���Hwq��4Z��u�ݑ�":�'|�)FG��E[����
mjr��O�LG9}-�-�_&=g=�E'�Z������T-v�:>r�X.Cl��D�(�T}H��4�eT�*%.R�� P�}�U���؈����pA�Kqi|�l��οU!F�*����w��X�J�8���"Xi|D�VNv�HGވ���+���{��1)��҆�kWNa'�K�K���Bw�zᇸ(h�a>�&�(ҤQ�oZc���d��#����v�n#��C��?�M���	@̩H�.�amN���g�H�j��xh�r�3���w�Oa��L�������Ɉ��<5k&��*�v��T2s/��}xB����\[s������v�4@렇�EH�������`?�PMp���Uѭ�I�˷4��Ta}�'W�)�/<n6`9���\�=oG|����"��x~��$�\I�0�w�&iGe�AF��l���X�3+�Ǒ��'��_���{�p�Ì:UD��_����#�^��d��R�A�;|+�lQ�iV���%��A�66^��a��(B�x�� ?Â5��;x��ڂ���.gd��<~��X�ȓ}��a�)K5�KO7�Lb��_��+��C;��	�^�c�w�0(����[��]��Hp�I,"Js�����Z �X��r��2</m��?���8�� ��M����@N�;ʧ�î��cJ��^�F8F9�!҈��k �_JV�_�s �����jD��1O�N*��	�a�Z��pўyCF3�����<hF`���s���)֐��jг���<��Uk��!' ���M�ז�3vԞ^ғ���{��F�$����u�8�yB �ɔ�-�$�PI(��9���i��Ŀ.��s���^p�E��8)jN�zY�}'9�{�{$q�J�\�qs�s:��4>�:G�:w�n>�V}�@*0L�=uAr��� k���W%�=xS������%QA����/���Mk⬈��w{�y���=5~����b�vb�1�[WW51��2%����q?[�$)/>!u��{���V�^�g$�ƨ�r�#�x=\��0��.���1K��z�4b�o�
�'8D'����I6�@�e<�@��o���
e�R��˖�N�4G�X�B)MA�X���%_q5�11ni}�q�cZ��q��|��j���ڙ�U�� �7���<�G��8'�5�yE�ך�ڐ�������Q�i�Q�О�V��F���{� ���U��/���qy�Wr�0��p��`5���r�g��=��I���r^���8#�yk�Nv�\CȜ&�cc�� �u�z<p�	�Y�8�v��dH��(�30�iN8�K$�Y��*o����(���+��}Q����q�T�c��W�6�t_x�8z������@Z�c֓ePb<�p�fJy�זVU�G�����������X��0��?��2H��=/���O(*FV�c�vT����Ur�h�������&0����W$���3�NK�4r�nGT�*R2�c��s����\|ޕy0��ˑ&������u�˟d<:F�x�<��	��ޟ�Q;�U67�G<ye5+Hy���5��� 9�����.��1LP����-h>=:����F> �-oeMw���M��.��n��n1(O����n"n{��^�8'���[�'�]�QgKP�;1e���*]�:b�z�w8 -��K��̓�Y�;�܂�YA�f��ҴX�G�n7ZZ<<P���e �����PF�@��G�h�~77~�[o $�]ݴ��M��ipOJ���?;�� '��QX�{���tY.�#�)����C�2�ҞJEk9Bz�*B�Ρ%͵׊D+�I��[���_����8�&�R��Ců]�W���"���CrrTc"b8��>IAb�eh(����u)6�>EY��H5F�݌Eyz�d�.�I,$+Q� cx4O=5fS��~��)H����\��Ğ����g7owG��{����ַ�Ff���l$�d�A��H���lD�

���Vȡ���%hR�4��هS,��|��K3����*3�;�Mr�Ģ`U��N�W������\�_�/��\�]iW�B�(��ހ��|�����k7���[��Ml���(cQ����;����1���@4X:#�E]&�Yջ�3ʦ��E�Ϣ�����x�כ�a�a�Qh-9z���D&�(����}t$�Gl=��;�d���a����緱_�`��&�|�A�u;q��a�w+�mg�ĳ���[� �"�;ͯ0�䲱�-���C��@�g��m��#�
܊�8)�h�ع�I��l ���'t��O6��}<7����moT��ib�b��f�􌡎P���d�:ެ�h���H-��fթ�h�oz�$��M�P�s��e�A�G��
JO�%�T-�_���6�Y�n�_�)�����p�Ux�z?C}%�3\�J`�9T\�����:6�]t]��8Hz�w�v�W�ܝ �+��!���`(��՗�"蒱��������6Ϫ~�t��5�R�$$��6,���T����)c�zx!,����@�Hف	��+�� �.���ÿʁ�5�x��ua���߱:OӅ��5õ��]i�]�����_�HH����h}���~P���K�/��A�S��/�n�4�:p�<��a��of��ٹʚ�==����ư�0��ħ�/^��.�V���ϸ�zL�Eq$�^�oR5�<��(�ux���аL��.�Tn^[x%�לmKF�N�7
E��N�[:�b���FpS��ۋ�t��gC5��Ig���e,�b�4�u)4�8H��L���^?����&Zk�`eʀ �ܐ�o�{�|R��oB�� �R�?�;q���'X'�I���j��Bƫ1h�oZv�ƣ���|�s�$�u�W��?9��_4^�V��㮁2������6�Ztb�m�dl<�Կ{��[�4e@��sN[���j�;xb;�����|H����8%��P��3j"�.��
{�0������DHD�wl���b��	?7e�5��R,���|�¯XX���	�����d`SpY�r;�����	g��Z���7�i�\	���� ��QV������;�RӔ\B
�H�=�H����r��1�}ֽ��v{����{�L�q�cR���X��>��X���D�uqڮmx;������`Ӆ�����T���Y����VU0H�,<�%�1F�0���:����Ս�~bBc�t�D3K�^����0���]��C!UM���;�ĭo�h�h�DȪ]���dUJݠ+��Ae��Ql鬼9�tk�ho!���{�����n�`�0��3���/Z��}�I�l����6��w���2#�E��X���U��B��ICIӺRf��M��@��=�Q�w��$'��lʞ�+�j`Y���N:������I�v`ҡ�h�O©�߿�#�֗>l��\�#{���=.�cJ�O  �[�D!I�$(���"�}h-��	��5M�JV��ӯU���$�l/V��Ֆ-"���Z���jQ��`&Zk+U��\��R��P�eKBށht�ܗ�gD���H��� %-c,[ӄ{f�q8�(fE������Y����B)�l�L���KJVG;_�@��T�vRKX�׍i�#��� ��g
BxR�Ғ��,
�7|�%J��R	9��/�_�*V2&���+kVL�R��t6�A�xB�?J��O?�s��>�A��[s��q����z!(l��E8�F���.y�J`�9|�T�Wm��f���k<E�%��������PXƌ���5L�����}�x�hgh�#�p.�l��n=4 S��	!��T ��҂j� ������X�T�u��)r@�66/�,���� ��֓�"�yRZ���Y{(�փ;!T`�f��3y��q�m�(�+2{�@����?d@�����1O3� ��y�� �.vpO����x9�ʯ����7ۛ4�r����C�0�}F�b;��~-��gW^��v��4\�,П{du|(49����InW�3�7eH�{=��,���!X��gc�,��|!ns��>����*�J�Z5�FN��!��0б�K*sYi#Q3(�WF{�(`�\G�|tq�e�ڈ�:m�#���E��r���8:4��Wz�GšUB��K=v�g�#@��F������/V@l��.��t>�	�����V��VH]83�Q#�#��]�/74��8�eQ�Ĭ���sU�A!TH�UhKX�.M�:�*�.	��;�=.Ͱ"N�P[8v٣Ӛ�������x�E���!�K�}0��m��>O?�B˫Mz)��ax�����0{-2��b�Z�4�@�K���F7��C�`�ΐk$�>����p�q�"��QT�Y���]
+�iv݄�
���S7��Wrr��kP�\ M"��m��_]m����RU��!&��ڱ��N�h��Y>�ױ�
̙�rË���Mە�~x���x���n�^��7۲u�#o�����WO���d�G��+���:�B���=���4�b����dYhܷ��[}�Ob,J�  ��h43@�����	�$���d��筑S*h"�f��3�t�<�-,�G���?5� OԠ�|Şq.x͊'7g<�,�Ȝ���Y�>*\�� �i|/1����n����̚���4�$-k/��5V�:�m�G�T"�ģ"���
�^+	�/��Pd�RT�[c��ƪ���0�kُ�ٔ���V����O�:�WmF�S������k��>\�
U��4�1\�Q�>W��vTy�d�EKe��Y�^�R��b7�Q�K�Ahg��s�&� �{7�>!"R�u\~r��˿�K'�a�>9+OO�_��͋��wx@�>��z�wy���"B�)賟+BGK-_H�	�3%Y�:�!W���'Z��i�|)�4����G�ǝ�c�A����}̮?�Z1�$`ҷ��]л#�H�`L{��(l�gɇ_�h������h>��z&F'�xȵ�YXo���ul��6�`�~e~��p7�ipb�����t�`�ْ$�+��p��u�"dN��[6U��
�c�-w'��/k�ryϠ�2��g�"p-�_Z
�N٤4�H�1�i}��eט��z���������H1���7�v�ӆ��X�%��Bg?��n��D*���fx�,��R�e�xPY~CAK_B���/�>5�5�Abg}Kߒ=��z�X\�ES�0�I��Vrgc��� ��;ZTn�0>�/z'D]���[Q)�Q��c�����5<���ng!��� �����)n3����	��ۮDYt��%Tn�1��e���.!S��4���]d����y!���{V���{V7�{"uLc�U[D}�m{��ݔ_ػ�J�"͑��`���1F� �깼�_D+�2�1�w.�?�0 a�X(�)@�B6�^-�՚�j}t����a��l�3i�Х�n�y�g�+��@nI�Ն�=��q�w64��:�;����d����'�y�=�u��7\>�5���������:�D�#c�d��pR�If�:�N��3	��Y>v�qwa��ɇ�#f����˂���J��=.��f����߱��b�1_��I�[�����ȵ`���Mц�]h�$���5�����.�(�D@��3��)���0q*5��2¤���2������E�.�C��,�猽ye-ەc�Ռ�ԐJ:�Cx��mO��d�ϱ	�癘r�V��������X��^�(o�v4y��V�f��@4��X�I�X&̕�R\@�X@_T�S[��<��Ѣi��̜�j�nc2Y��8��0RO� ��r���1��wr��F��6�o�]�X�=F.���"�=�0]C�'�[/��v_�p�kO�cZ�I"}��ʄKx��4�:F=��'TPg�����R�=z�+��~fvA��c�D%�D������W�ĥIx�A�a���V�2��5ӺJGO����2����.
U�C����l@���aW��3c�S�d[�S�f��\�u����D������"��3��4�D���-�hο�����q�&�-x���Ϙ��2N
HE�k�;~?�M2:t�V��I�1�f�c�0���6������Y���|Ȋ�sR��D�:�a2�h�}QN�o5|__Px���A��t�ހ�Y��B4ҁ�CF��i�Xp�#K�J�9+p���&a���Ý<�.������B�3Q�8x2�*�� ��T!p�פ�^�Xj�S��9DΛm��\[��;������S1p���$[�.@��R]�0�o��C�o��i�|M����s`*�������0�LAF� &E�/��Ψ:ݴ�,�����5z�|��,1HPז�L�U%�P�W!��mr(mt�,�y�k�<XV�Ï�4-g ��ߐE9!�t̹���j��Bd�9.��+í)ꆶc��"�ɀ�}��*�:�m��5��]�3Ĵ�l4�3�OA^4���D^�q���3��Ir��0�X%[�	[<DA���Q$������!C��@!�5��R�R�<M�N�
�O�C�ʁE���R�6��΢9:u��P��������pK9É�g���V^��e�}�%���'Wk`�:֜3�&�c��)`��;C�;ė]�ʦ*�1m�Ttq<4reT�4�Y�痻)�k'�d�=�V��"�&��\������60 )��� !�"��S�)��ͅըa/0������"����?-jΧ��(=��g�V0dh��sjED��Z�Ԯ��ݧ�JCnU���@� p� �*i�n�VnBg뉓K��4�g�Ydd��$�4��{@ˬg�wo!�M_$,�)�<�9$lV��HС��1����~�f�@DB��y��tZ�:m��-��]���]���"!�������A�^:��).���μc��{�Y�1��7	L�b6�셰d2�����)r��b�yҤ�״Z�+5����"�D.�bn��?Ե �c��´���Ҵ_��o�-R�O��f�Q�`Y��'�[�{M�������!ia�����h����\>�6�>��Τ�H�)��^�¡���<Q4��]&>6�CNz�xu{X��p�6	5:��y�h�>��ϖ����9&2���'7��Z�7�
4B
)������]
�
PiYx��b��Y��Bp�6�.%j��x�RIJ��L���}��w�W>>��p��ߑSc�eW��g܇ݖq�~$�[1 ��9��_O<:���me܆������^��Z����:`-���h��d8WU�;;h�xf�뼕t���q�M��֌0&�-a��q�ߧ����X��Ø�+k���ۑ�}G~p�! �\Bcv���B�o��݌^��q���^ミ�
��iU�H�:@O{���O$�_�d���F?�"�w2�@W����h$/��}\��` j��Y*�����Ʉ�qo�����W�_E|a����ҁj�F����򷲛�5֝O���$|�i����91��Ck�z��	�bϋ1pВ�����x��a���RmI�lj�	z��Z?�>e����a���w��nfg�R��6"i�Q�q��G_P�]�@�3�r���L�Jz�r���|Qq���dN=4�UdIb��<��L���?r7�Wlb�s�d,u�pnl��w:[�&tMT3�#V,�z�e�
��8�Z���^��A�=Sf��	�U8�;5ˏ�l�^{؃h}z�zY,P�2����4Wu�Х�pS#�o��{s4�.Q4, ��9�.��y�����'kL�U7�Nh�3��IX�����iu;��V��|#���I���o�{8Ø�WWK�&��G�ljM���:�f��m���<�%Ag� ��n%׽W;��F���^��~�|�ޱ.:R�S��X�&M�f�̰mH��rA�t�6������1�J��#�=���od��M���L�JYC�pt8�"���:��NP�s;�Z�Z:6у��X&c��w7�u*q�����J�Xo)a��+I�&1�|�!��r{�򛑢�{��x:՗���7��4C�d�-%P��'���%;��(a�R7����������8�b�Zo���Za���N��á��e��n�k�X�
�YQ:����P&��+'��v͚�\�V�`�"Pv��hy�lE����'��{d���ب�b*�����+�̸X�p.Ô��.��}�	��Y_JSg���p�F2��ً�T0|Y�f�T�����y�6�i0�c�$g���C��.�������6�F)��'��4�{2�<hh ����q@U�{ @*Rˌ��h�KX�~A&���u�$TQ����:/�"7��w���Df���ői�Y2X�i_݁tB��5�ɲ(���Z^���L����$mR�� E�3H�@��El�-H��3��F��	�~��#����#�A A�v� Џ�����:R�Zؠ!f�w��]�w�S9�^ՙ{�&�c
z�>k�r<@rq��?�ļ�n>D�?\��=ċ�@N��P<pZt��C�8M�2�E��|���+Z"�ݠ#^՚�+*q5�~&B��,GK���%���%}��=�D��|��"�=����Xy�`��<Y�Dl����S�Q�����ͅc�� V�-ud�h�f��;aqU�uԑ��_	��D��#��<��Ѭ����>�\� �zpb�%:I�DSbo�A3z<�P�@�R?N�8�}���v�R�w��x+M˪�F��Rt�e�FDR����%�����ǽ�N�Jo�YOL�.uRa&�.�Ʃ�P�qt��x�JpA�U��0����e�F}��t�\�/1�{2~�vR8���f�J�2H&��j��9ii��ȡ�NAs��63������b�F&�"�A�2�Z�$缾�3�НKj��;=k�����e3�Ow~�A�����/�f�iV+})'�,����&.��	X��I��8g�����-�s�T&+�6'�б��!u�7���+)�?jg��\���Q��4�������+���{�zg�B>f������3���勎���v�Do_;�jO�B��� ��y�|��oX�3�yt�����[�Z���/�N#o���l�.�0�7���[�p�Z�.�Kڸ1 �6�!�n>\�m��R�F�Y�_.�c���헲�.���\�+�H�䠴��%Kk6�rUeY��>;�����s:���?+�l9�DWΗ^��--�W�?�*R)$� ��X� đ�U��듊{�:�g�5W`A�z0)%�-e�Go���+n���5 '�)�[Bk�D@�6������� �U�R��?����/&6e�y�`a��45��KA~�}z���9�U��ۄH��S%[�:���UtB��/����-��`A����N#B�:G٨=����M���L���@�¨��Gc�Z>T�9�>��w���&�?��	���-�l���Ƃ�i�N�t�a��1���4;ЗjRӱK��y-n�c���*L �X@�%�"fWز��8�O���<��gj?��J��9�Z4j���15.�Ȱ��Ϣ��貊q�����s�9�l�I7��Tu8��K[<m�?��߻��ta�ZhH"�"��9�pQ0���B`�j���f��oA��@�Y´��S�T��K�~�r5�	?I;n���MB���{a���v����et2���s�}/F�a)�@J���
��EAj�	�b���A�2:���8j�>���F��X��S&��&��3ڪ]/�t���A�&g�5��E�7���=^�u�\��q���԰���T������%�	2/�Iͽya�u�J[�f`�9myW	'�~�GR誚�hz���zPj����s�\�,ƫ	:poe}��F6�"��֙.�+�?ʷ����?����|���[Qr�������D�3�|��1�XC��7���4������V�\��Ā#r�ǵ�H
��ǐ��D��T>�=�X�7�M��u^�:�@��lx3�<K���bA�~�^� ?[�6n��c��m���2[�P�
�^�z�j����e"l~y�tiʼ�H"E�&�mK^�k�E�X�u/�ݪ���o�I
�5q${���j�������ъ�A�����B�R!ST�[�i��4c�����7rss|8���U��֗����.����:'b�|S���1h���+5qkm�W� =}c?�	FI0�J�N$���E�,84đ7��R�@�`nj�|e�uF8m�F�sq����]@�� =cq��6�T���*���q���4)���Agݜ����\^�~$��#}�M<F�l��oxW[�.wk��bǊ�	��	�����n+A3c�Pxa��>׏��G��j+x\W���&�`����0������UA�L�H���E]	﹑�I׎�i�[D����_����n�b,�k��*\�̂%i���)!��&L|��s�����@�|���+!D�[ #@���`��r0�}���ɔ�j��k©D�V���C9��`��[���A����F/6`������Y��_��+�O����N��&۽����g�+��	AD�=9��1{���L���f#;K�i��]�B(�/�`�(�u�{��k$a� ���IpQP��E|�#,��I*\aԞ8�p�#:tM�]��l#�$S&���=�$`$C�YO���I9 GG*tы��r߱�"P^1OMc$L����JG�B��4́��ח~k��g����Yl�=��ZV<��E�$��g��3���(���3 �2�cw|3����6w���|<Zן�ֆ&xQo�N��1��A[�ܔ\+�f*A�q�:�	t�?��OT�a����(C��ǱT1�����il��|\�����x*�����{4e5ֳٖss:��/�V' wN|�?L��,���\�QK���/ry!�ezkp�&���|���� qZ=�rG�����L���PH0�-W��������\�b�����ҧ�~g�C<�����Y�3��A���fkҷ> '���b<��|t�Ñ85�ߟ�A���F*�<��/�X?d�ة�O=���'d�����[<�/����鐟�� >�3��
4��h#y]�E��m�a;�4��7݌��ԅu͆v�y,=:��Ӆ������F�S:d�N��E�	�MD8�&�~!oH�;Sx�+�U�e�������e�g��1S�b�e�-i�;�����P�ҫ薍rV8Mq���邝��]�ǲL����?4I���7J�<m������H��;��o�Cܧ���:7��]$r]�pF�����A.Zx��[��CSa8^�*���bL���-��J��D������c3��K���#����8��LG�S�ș��G�~9�ŉ��s�
�O��ŉ�i�Y�����vJ֏�nth��Wq�j��A,�v����1sR�0sG}D��f����Bmb���OrL��|Nu��.��,�u��ݵ��:��k/d�g�+�KN�tc��6�d%5"bTo���Z^�K��R��i�\���o3s�L{�1UC�wp�#e�>�q�VA�zH��;�� (�Tb$g��r+J s�����ʀ��(ּ�>��]?����6�gmQ Z7!J�'�O�����-�I�+]�$*�bH����S;�@�&$�ބˈ+Y�s%Ě�J��C0v>t	���5j�Q�{$�ĵ4G��!GX�M]j���,��n�����l���M��@Nm�e���MC��p��e�r8�A����u9�����D���y�(�3���� u���&^T?-YQZ9��7x��7>]�qk��nzv��3���k
��=V>��i��GP�ULlU&Jx� ���"�%?չ)��<�
en�bv���ÛАLjϊ��ۯ�7���y���:���-Q�tU ���QG}���M�^�h)�^"\��-���gbz3�%AP���]������st� R�N��'�%;��6n��[O�L����2�I�4'�~D/�'-�:bY� H����䌲�D%����jl%��?۠�T�9jC����aB)γj�$	%W�E*��F���D%�bpҘ�Q.Ңn�c��|,k�!ț�w�B;�*��;[��9i�`��(���1��k�����x�Ƙ��$�:�n��2��_����eΚ��"W���K�b#���3�k�+�v�vVn?���m� D����j�-�����"<��	uI�i��vs�n�z浬�⻆r��)�:��Q(Gw���:CJ�ݹ�^�����1U�6i-l��qҳF_`�ٰ�3;���}i���(Iq���'���@LZ7ڷ���_�5��:j��[�勹����i�؛X��V�Lh2�+�S3����ݕ�=���I�V6�����uM��:04y�0��^�\sL�*�fi�;]�I��4FQesIDLؗ�XTpj����,��у�xG�����̤[�9Q��P��D����m�T^�"��j�:I&��@��l���B�����Y>�im�L_����� ��ϕ�-'���%��-`��d��ol�%��o���{/;�ʞ����
�z��t�i�[�'��$O �������1X��F�/H�8��?L,n��˪5=� ��D?U[)E���Tȱ��:g4#,�tl
����������9�0�$�9���Z���0�����b_�������]��7cXI��	��Y���\�|���>
����ū�as�Ź�W�ӿ�;H�&����)��|���V9��\edt+��\.4A_H��Jk��M�z�~��Uh�U�-�M�Є8�z���N`7 �|m��rD b
��,��]L��,�ڳ�X�/�&˕�{�f'ސ�&Xo"|�0ԧ4+#�U|�uw�?��,As��iU�ԀJ����L2�k����*9�ٜ�F[��l����U�%YD������j�|�H�{1O�n�7\�o���\ɤ��Z�g��9�ڻ�y�,�/�=�� �-����u%�UU=�\z��3����q�lVeĥ(�������Z|��c-j-�
�ġ��Gwb�%��x��<W��Y0���}f����?��'k���z�꠨�9<�w@\�d��������ٕ�#ۼ��T*�aܽ{lß��F�(x�2��:/��8p�/ev�����̀$܈&�Y�ˊ�h��!�D^���[1̐���fF_��X�d���kR��$�ɜXأ�j�]�{��#�y"�_H��II�^�>D_��(�񛉧 �,�����$4���)��յ��8�i���W��D�����TQ��W��V��oV���=ֿ�Ǉ��,��U�ݩ j-~=�DSx�O�#-�O�]]�d�y�F-A%�!��Gb� ��k�"������9r���T���;P�4W�Z�~�!�ׄ�x��asZI�q�t��X��	KXE��ޤ�E�c�n�W�g5Ӽ���P�ZN�|s^��)��f�)ڋ�VÖ��Q��ҷ6��<0*#,�H��3�1s�S�6����F�S>o�1)�D�}��p���� )�  �c�d�c�pA��Ya|����`?2}�"�$�W9_� f��C�R�c���d�$�'*Uq7l��Fʕ�W�Q�{�O���wz��<��	p���\dN��Q�~	����+��td{P�o� ���C+�26mI.����r��_F��T�9_ �=�����t�7�c,R��ԟ��w��!�F���.Lv&4��2��U|�ѺT�0��$�������"M ����=��D�oG��+W�	�_�A�"۱�_
-���m�Ḗ;ٶ����R-�%,];W�ʀy��7)�����aSR���~KO��5�A��ȁfřĐU��������2�y�E%Ἃ� �r���uö�@�����k�MK�}�?��^8��I�q�_p�����d�u��iƣn%M{��,��H��Mu��ġ9�P��_-t'�T�q��ʳ%�ޙ��FnI��c���k���!�/н��e���ܐwVY�b}�)|6;k��睷T�)��[]G�!XB\�S47��A���S��N�tz(�����9�I���� ���������F�K�;��>�Wxh�]���� $@�BuD�I�������^I��}�ע��T��L�X���M�q���h������Ҏ>�Kz�@aCS���E��rp1�Z���@8�+(��.�C��݀80~�_��;�^������欉)8�k�Ee�@+bT��;N��ŀ�����؊�C�*C���h�\�����f஢����]�D��(6r5��?����Na����Y�]�bPK̴�3Hq��r�-?5[2n��'R�������XxH�_,2�<O�����M�/LGRoG��>�PQ� �~�������j}؜QFb���N�J��I_W����f|i;j�y��v��+w���H�?Y��J��LT��(����x��$v�Ƣ��&���.��lV5����i�`Q[�̨����n�W-�qR���q
��������ڨ#���Ʌ���`��q���-�Jp#�+d�mE����gX/w�;�CfB9�C.
�ѧ�0�b Kc�j�+zS�n���)��9�w��k�C�y[}�K�3�����=k�'��  ����~RY�d5�@�1W�d?��yNj9+�qk��t�+���ye8&�Q��tW�(�k��V�~�X}�#����X�F��{�ed�:ASK���a�B�К�a)tL�~!��4���M`%�-�FB�U�H�v�*�'�"�^�k'��E�::+���G�>X5�&���N@��e��;��U��Es�� ��v?˥~&�K��&���x=]������ʃ*�S%��e�9��(�u��H��Dܴ�SU���J��w�TMZ5�x��J���D85���1��}q�~��y�F*$k��pzO,�F	I=��<�멈��0��u�B�6��nC�Xs~��������֑�C:�^���������6��97�"g���%0�S�.�sV�D����+������݇�>q3D�a�=>f�<ic�F���\�B�6_z�\}�M����|g>׾}����{���?�
�� �,�Q�Y�;պ����I��h�W����咮f�X��I��_i�|��N��]lr6�|�ILp������r#��r�7l���0t�������� W�2GP�(^X�z���x1N���
��]�Zz��E���*Q�B{�ak~{�G������"����h�=�A[������}��XQǭKה�Wz~+�MVu� �������h�������3����̰��{�=����W9Y���L��t��r����eޫ�S�=�4��e�_B^"� "���=�X��b�s\�!c������y ?��u���
���[���;�1�1�y/t>�38T�^��Ƹ>�d�%��C���,/�.L+q�Яe]�:�+,�8��M�L:�c}?J���,s	�2�I@W�p*�����J��(,�Xhe��3��c@��|A7��V��%�"�����
m⻠Q|D�PSU���h91��x�o���ـˠ�� Vj�Q�DA��=u�����D3Rˏkɉ&�"�����j��z���?��y����}����tBt�I���kb_j弹��(˳� :� ����vI��B]무hK�������:�ը~
ee&G�� �a����9��ĩ�;m6�
�ӡL0�e�D
��� 7�_��մ0'�I@0��z7�����|�(!?�%�_�߁@��R�e�d�ݞU
/F6�o+qL���08�%�%rI�9�s,�q�`ɬ�>)�O�S�JXt�����ŧ��v21���t���;���#���� �B4���l�d������7	�8^��ә��'
d�p�8��Yhy^Ӛ�e�:."�k���?���EO�3�+�V)��+N%�`�m�E�(~R$3���*q�˶�Ы�)�Q�=Ե͒�'�>v'����� �~��*�~����ӿ7�	�0A���������/���Spj�h|u�U����JlW� d�0��awh�4ɾ�C�i��HV��	�h�(%�$b�p7 ����I��[��(��w��	Q٥���@ބ��&0�o����k?\�	��2�b0���je�D�T�u�U����uȘZt�F����������h�A�O`D��i��ţ?������c4����\bF4��&\���'��#�b�#��Ǳ�$�Pc�\U�7����K�3�0��Q�ϛU:W�ݻW{ta:�%�<L*��d�͏2�:g��we�ơ-P}3�m"W�n���V��s�Ddx�?�����=�NI*Im�O���b).��9���\%������ۛ}`��L�bO���J#��:�|�x�䄤�s�
<~���_��~0��'I,Z���B%�����,��d?�.����I,�Q�+� � 0$'X]8h�#Ӥiū�P�/m����X�!�ݶ�#�yC��
�O�/.b^�)���qm{D@�'}i �H����� �4�W�7�U��=�޵J<���z�W�%r��Ȼ�Z���~���D*�,���fv���mY�|�w$��G$�����Y�7��]����fd���D��3�5��k�X�X�镉�Q���������_+��U���t_��z��B�i��Kp�ЕÃM4t 0�o��@Wގ��:!C�p�T��쁯4��נq���f�0�q"f��|�Įjh�$��������,G���p�[�%�?  �{������k�t�&ȋ4��Qq�
�°�������+��v<�����D����rY���{����7e��-m*S�%�-P|!�*�oS���C]�W��pA/&�
�w��TwaǓ��6��I�O��E�f̚�w�����4�����
�ֵq�( ���ݐ-A��e'���)�UM&�+*~d7��Ej|�䖠R���h� ���Xd,?E[[Q�����׿�0��o��V��r��T�!�Ś{Z`G�05~?z��i����l8~,�j�y{����{�Y�)r^���}/�IG�霦��֭�a��Z{sZq����"�j�N���"�D)a(}2\�y���{+=I.Ħ�$��Y�Qr��|��*�ű"�����~Я��O9�j�K���к/y�k��"�Y���,���fP]#�l�6ر���=H�P2��W�z�A)�r�z�IV9i��uX�=1ZR��g���2Z�s�!��~R��?�⒱�L�i�P�7] ����G�a��oΣ��"���G���H����
�~�����s��e��J�"��G���'��r��:��+�0w��U2��A���;j�#������(�v��BRR��x��o"D�M-���_&fV���ʶ3�
� �֜}^�/;����8Yg�1��\�%S�g�#Mkʆr�y�>���jLd���б�{�нl�D�R�"�uU�#�SWU-x�A�DlH��o>"�:U�z��ʝl�de|,R�h�4�
6�I.?ɀ�U��[���Q)UL�м:�I�9ዙ�䤰 ��c�ߗ�^����D�(S���yqJ������;��)�z��E�vd��n�J,H�{��%�-hz\G��2����
�K�_�D%�8ݠ	X��|@l>��?�a:(��wC����=��99�3S�f�������yz�%�m�����dH�s+��n���s�_��.@fjZ�C���zj��K�VL=�9��F�m���W��i��㙫ީ��`������1�c�%�� S���G\+'��ڂ�$��}/���g��l#r���Q��:�4*��W�?���H@۰9d4mip�0&@�����;�!�`��$^��s]���=��O:�����O]Z�I�<p��^�@Jc�Q�e݌�����=@޻d	��}�����a믿�N�V��_�E��s�p�pp�>�b�?�	g5��.R�I�wl��vOc]�>Ȓ�L�ek�w��hf�*PO�|�H:���>�𛹡P������#�`��Ǳ�ʙ��m��I����H ^f�����(����֐�z��Aתl+�GP�~W��F==]���V�@�O�ڦq�xo�
�:.�j�ƆM#�Mbg!#�A����tI�T��:�.k���ө����](�V�A�b�	E��X����* ��|�=��u�4+�x��gDS������[?oJ��߶}!Z�rsϴ'ῆ�k��6����/�y��w��(�8):�\���rÔ��MU�X�~����{��n-&���Da�$d�=���iݝLH$8���W����	�W�7@�c%��YSkY.Y�c��ϡcU#o�f�ѷ�g�<��f����M��
�d�ٮ��I����>JB8!Fy��ʓ�U�:��)�����q�I\��E	��� ���n�/YW�[
���+���j�	G��*�NI�֏�QW�th]4�"��`�"��/#�nF����2J�ׯ�S�E�R?1�b'F<˫�2�#���"�� �y�5�yWS��iŖ�0��@���a��2\MZ{��4�B3��9�
�y]@2��<ߟ��� -($�(��y�ڀ �[�����L�,�����@�ޮ��&�oБ�p��H,`m�a��r��N�Aϗ?�iD�a/r�'�O���x�����P:�#�׈v�P�+��j~�$@`�1<��&/�Eх��>?���e����;o%uO�R��ZpiO՛=1s!S�T=N"�8">ŷp�-~&~-Pt:-2��7�]y��ˎ��6�7��Ջ!rDв@Vh��Iof�7�>��o�@e���[�&�|0�(&(��KR�n�?9�-�(�\R� F�:f�S�
c�c����%����gPz���54qk�T�!:'���^G�9��)�uC�
K�����'o��2�Á�ֱ���`��X��\Kl�LJ��OVY��e�����0�4q���3%u�T�]�l5��")i�8{;��!��	��b̲"NA?����4(��Q��e���8:o3Tp�?w�pT&kV��IvR#��:�E=�`�O�/g��¼�
)�#(I�`Ւ��k��ȇ�i^��������SFw��ʣ"�r#�B�X<��elO&�P�~+B�k���o��켞��<�g�T�!�%���+�gj^.w|[C�D�E9Δ��%XI|�՚L���=���q�e,=�G������nx~x�[�Ѕ��������!�Mo�8��������fwݰW[S�k�G��ej,yM�f�ABN�Gk��z�����	�[^�4�	=g�
����C��Mn�c����n�-+j��ꖳQ��Ks: ]I�Oʧn�$><��S�8�Ϝd���zONUNW8��a��:�`���(��� 5D1�[� �o���O���¡dTX��U��3!f6��կ���{2H+#�	��|�,�¿��Y%�/�'@�3.�#�.� �.[�//3f��j��M!��˧	��\�0:�/sĞ��UoP*�3=����ι
6���2�g����3��6�L� r=�^��<�/����;�.�3n�)��~qSU��U������մɓ6���M�_�F����e��$z{���)X��Ig��}8[$��!9���?q����Ю�.n�N����%t!����Z�K�>Na�_����8Z@^ ����O���;Q��#4��,�oɎT����	�c���"(�iJ����=>|C��|�݁ &�V����Yvj^�c���m��4�ѹ��+�-й�_�P���r8�q���m�2C���rLc�I�ǧ�I;�t~(�-�P4�wl8��\x��te����2֯Y`���w޺��W3<��%�es���)䘾��J���aQf\�2�1@��\]#�I%<��zI�>���4�9��ֹٟ3Խ�Rk��˓�*��0��f��{|2v�Wb$ϔ�u�Y}g�Ại���<� c���F���[K/#��~ �9Tf�^�~���[������)���Q��i�^;m�g�����2�[E/��.{()��:�]�O�}P�EO���[{���O	�S���X޿R6e��v��C��1AǛ�d�բ=̇�� /(��+�������gP�>���U���H1��!��k�˳}���!�_-S�ߥl���3\�w�KH��{:����7����_2�Q
~fp�;��%�f����H_я�%��k�o1)H�p��>p&�V�SS\���؏�K\�
����.��HS(��j����DB�Љ��OtP��;*������8�٢�n�g��%1���_���7&+�d���F9+� J7��F����F����$Wȝ[N~ol;��
'`cy�m��޴6���rS�!MEzC�t��h3r�_7�E�u�#�4��f
�>򐬀�1
2�,H��4~�.v�PV8��E
�5a+��l��`��Q����Uw�HڮԚE�H���4�i[9���X�bc�&l5"g#q+[yf�X����_��t1�d��W� ���Z��$�ʇ�����8��k��2�95%�{� ���x���~��Z#������Rɘ��oD�ᙈM�OJ�0�!Z�V�	0��cD�Y=<ei(D{�n*"y�����+�eyW�S}.�U��L�f��j�Vb�jLm��1�@MDz��~d�v������B^�y/�:Ɲ?w<br��vE�y��*�,5iQ�����W�FH��٫M]���FAh��/�%�ch�S����Ex!��)-Vv»����Xa�������_��ԑ=F�H�x��Hw���{|ͯ��H�O�8pK���_�̀+��/r�|�_8N��Aj-7�59Xϓ/9h\�;]�@�E�+���
�GP����,)Ⲏ�
 �\�[�q,������顦
�n�e\sH25��E�!��}����vѧ��V�w��+��U�����),1���p�b�$��>�۷���wǞ�r0���+X�C��b.1{#o��g�&4����z�u�i� s�?7��6(��3�J,��e�:eXe�g-/cw�di�U[�LJG�xX����9�el�Si6H�*���ȟ�D�POi+�OC`�In��Ҋ@�^F?	�v;�|�J�:�u�p����k��)�(����PUC扼p��p�~�U��q���vb� �m���ä��1�Bժ�4����{q+jȍ��|8eJ�N��'�gb�S�)=Z�v弌�������[ƔD�3������dp��C0- I��A�}�U��d8#����D�ɵ����e��P������c�,�8!ܔL�~J;R���D�c�^��J:��kc`Zקʲ%n�Z�3����2�� מ"%v�����ψ�����3��^k�/|w)�A�_�~��0����6��:*l��0�9,;�}aP_�<�XxH�L��|�OC�øb�H	E�ƐgB �k����!tu�N�J8�u~���:��O�W&ɀ�ܲ�|��Tk��b�b�P�U�"Y���w4�|�M&��Vg2����%7G�GH�_3�[t��K���!�Iyŧ�c���J3���#B;PDV���R_^,<+M����t<�x�O����9w�&*�]_������A�&�@z�mU�i�Ԏ��JB-f�4���B��r�aF���M/���5o��������K��4Y6'p����A��@+O�z���)�l
IR�p4g��Ҽ��V(����,�̡i����1��0�>܋��=��ՋB�G��໶V+£H6��m�Hb�V���/ �r�-�8�aڌ�"M}�Ƙ��$�1�����b���5�?-��n�4~ß䞡�z��~�r))&t�ND�WzYi�(�3/�	.gc�W~�i�b%G6̓�(T�U��B���G	�_�׀�(��޸��T�`��$_'"q!�>�a�ݛ�t�F�6��+��Ӑ��QXۈ���gyS}�Hj��\�ş	���:И�(aV���O�7Hś���������v��	".�i�
�VW�k��S�S�}��1E�^n�1�n��yڽ9�4��ᒀ+����j�aEq���e�hwh\a�PtH�8���z@v��jW�\��g�G�"-���zP�bK���*�d��9"v`�PDո������� ��LqDԆu2$�����*������=:�|d3����[R4b�	�%�uʹ�4��� �I*�q�nq���}B۵}��z��ԵLu6z<M2�	̴��H8kp�`#NO]k
:qi�-Z�B-b�{s���"4��g��'~:��U�)Ӥ� �C] �Np�ZXyl�|��g�2�{�(H���[1���J�\��8�Y�dI��(&Z�T��P�9������/
�Rv!_3y!��"~���p�f�Z�{G[>׈�A[$���d�W��DyM��u��WNhin�@��=��J|�N0gN%v{j7���31��9���XRPɢJ��}T�I�/1	��`ĦF�:?�e����[�T�c�E�"��b7���z^�v����0{�1TW�D������h>az��gu�� Ԕ!N<�����e�L�J�l
c1,�ڕ���9bP����M�|"Ƈ��G�M���ʓKb}����������>��T@��;滾|�Fy���zM��IȾ�_�_��[Q��/���b0��zC��$�� 򰵺W��tV p��.��1d ��<n�fԟ��QaY�|�`�s��o^�i�l���0~�s,B�����0���p�F��X�qC��.|�"��d�-���]���Vox	��5/ ���G�����*����l�[��E#<��Y��i���Q�e��z�j��Z�M8��ĵ-��%L��M��8�r�0�/���O�^��K�V���5��"��Q���|�e媪W��>J�-$��Uջk��ZO��c+�%{�Ʉ2�����M9�x�m�f5cJ�Ϫ�7;v��++6x��S��D(�v%�M��s�F0TG���T����5I���}W�&zߟ�$���5��n�`%���/�����$ً�X*,;�F��r9���������i~�<"�����
{�G�������p��5^n�-�`����*R"�c�:�n=��X`�,�oIic�0�|~K������hl�UWQE�G>A�;�9�2�v�h�LϏTO�"�幨�� ����L/��*��J��J*�8��SP��]�r#����^����& ��=����y��Ԉ��j�k�y�/2���q�²O�<җ��ɊF������L	[,׹~e�����'���4-�Kz)��#$����S����N���g���a�VF�B�r��:X�s�m�_Ve� ��g��父:�onBW�f�� \�X/a���&r+����!9t���ӳm�s��E�Π-��Ƅ���pT�Sk\.C9#�@bԋ�����Q����+��"G�D�a��&�������\mŇvS��]O՛�|T��m�ފ�~��-MW÷;iFԷf�K9i�<+���Yi=%4}�˵�J�aQ�o'X�/�_�Ek�]�!Dp���������q4;���Y/w�W>����3݇,�,��q�yh��Cmp��ɰy'�Zj��+I�Z���������A-���B}�P��� CnP~ P�J��y-ۧ�=�py����:x���p�/:Īc�-�YZ�g�A܋u[;�'�����ZޟYE2ȵ���TN�6�"h�k�fh�����Jl�E}kP�ٽ�&���Pݦ���̋�Y?O�fO���?s���jK�j�I�w�1VŬ���4��q�dt�&3�e��	<"N��b�	�J x,�QW�MS������i��68�J1�1Yge2a.��7����2vQp�x/~� }��(�f�Z�(���*'.c���/��_��3�';£�i�^A"����Lr�x��$Әi���3�����	��PUc�-����`�tk��-���5��/��8�����Em4��VB�Y�GA���}�ӫ�C8�h��1�1���rʎ%s8#��n{a85j�#5�4Sin�}Q�#����ȫѠ����e��*��4]qv�ِ�:OV����s�zU���P���x.�M`rP_�N{� Qײֈ�������[Z�*J�/��f�bȃ0*�6�Gk�W�]~�W��*��a7�ƐtPߠ ������|B3;�q�vR����C�k��
�r�^���p�+�p��?å��1��^�Y��1�4!����A%����!;���(|2,�E-	��#N��ND��̌K�93�t���C�a̭q���r�ݑ��bh%��}���el�1M����ޞc�{�tj�\a���Cm@a������I��,Z��YK8�%R�r���v�5���$��WM혧G�i��5u���}��ɲ*�rw���ݪ�Ŋy*�L� �ӹ�o�Mc�u}�Ͻp��P�A�݆�ԛ�b�>S��d�T��ȀĖk����yK�Ϯ$.m��+�8�O}����)��6�rz�B-�jJ��Cԋ�RT�Aljɦ���ڿ�T|zA�]��TpY�[�ߑ{<���B���xo��d�ȼ��;v5}����}d��4�'J}��U�uCX�#U�Z�N*�p�B��r�-�s3����z	���ԈP�;螏V�p���p�_�M�0U+84�
Al�+���
Ϯ�B�,�M�'gT����o[J4y��0�b�3�+���J^��5�G(GtIp\�,J[�S!�P��pk�8.�\'8N�Y��ٓ�o�<E�%d|$ً^��
?^H�X�ᓩ+
�]U�Z��;���U�,8���F�M�1�6��+�����I����A��0u3����\���Ό��	�f�XP�����uW;gIZ�l��@P�;`~/���� �F_#uE��9��w��+6��J�L|mMy}�������;Ϸ�#o2a`�³l���uo y'Z�W2��#p��/�$��	��ӋF����b���7��R��,���;�#R�J�x	��uVI��O����7J}����B2	�K.ϝV�	
 OE��>19�C�Dԃ�̦�+�$#�|��_6b�k5B%�{:�}�ȴ�'RC�T��.��PT�@�I'ڏ��ˠ�.��"!'/<��'�qԓw�Bitp�4H�\)�����FRP3�d�����U����{�pW �y&�%�]�YX��b���mwj,<���M[�nρ�Ne^q�C��Y\��̌�Ou�:�Z�g!ڈT�}N�4s�6�g�ɦ�f=C'*h��+6���8��<��Y���|��ݵο\��g6w��z���E���-zde���=ߪV�䜆B��"���`u�{�@'<���o�@�;$�|NXq����Vm��/+�g>��wv���Û��H@~+IeG^����W��y��D>�/8K%�b|Z���������s����yWXI�{��*i�� �{��=���x���E4�u2u��m�]vE�RqL�
�M	Ͽ7
k��Q��\��B�	�G�w�`�J�GY"�A�ddJ��do���hC�4/��>�Z�	�F07�0U]��p��^�P�x3���R�"N8��||
p����k&��n �C0�A�)�E����VZ�pz�Ԫ��
�T�
���^��U�3 �'��¶$vf�<]�-�rDW\��gi��(�8��u$r @j6㟥C�x���&	_�zV�C:R;�\�m�	�Ȁ8���}����S%���$�ﳟ��ݦ"ZzziA�t~W�*���zqT�P׸��J8�~6�#;2 �cI
���d�ؖ�.�UC������$�Af#�)Oo",������({}��a��W~��kI�T�7 �"� ���c����F�K6�b������ý��� ���UP�j�r���Q�>�Q���A�# O*��^@�U��M��9��
w�p��������#�JL��G�'XS]�_��0b�m"#�70M�_����a�$�S��� �����^#�'g�cPΈd��{U�ѺkF�!��z�u�O�Z,ԎM��p{iD��R���ZC�zUЍ�V|����C��UE��`���6"j.�6[s�?�(�/���s�3�BƮ
��s��&�k�JL��ݾt/��"v�$1&_�dFQҒ��+Q-Ӆ�X�hYfZ�H�m���nFÜ��D�N�5��u��~W�%~�{"�Q]|[��?K���AҔ�N�:���� P�M\1~Q�B_w�2=Y�%]1}��]���0J��A(�a�\�I����3���B`:�g�c��v�����0'���}�E9J\��^��?��G� ڄ���_���f���hR���w߮<7����Yq;��
�-�lA0��c�6�����5�(6�6��ei����م��2v��I�{[�k�2(�ȡj�>���ٽ� ���0WK]=іM�ǣ6��zPܖ{���>s�6�>/�VorCQ��9��2؊�������S�!#�Y���^��Vu��̓�Q'?��� �y�`N{ZwG��^ȼ�C�$ "޵㝜8�tM�3G�?���_V����/Ԟ� Ck�ثX�=qm������mq�A���l�Tfu�f�^�Յ(t��Y^�b�	@Q�$���x,5na��<!��?wyxUd.�v<.Wh��a���a���F�9F�l�aυ�v�Pi$�Z�˒��64�#l�b�Ռ���b�?��&6N�"f�������T}�yD���?�~#�j�*����z�|DV����vQ$Mx7��B����2g����8��4%�|ߍ�;�8d戺<Ul+f��0)�o=�ݟɖcY�s�G��$�w@J*��N]3O8�]��\�l�$?�!w��n�Y.)����@��d��`uZ�;v��3�bc�̂�:s�]'�z�B��J��8J��e�B��lJ,���?#�: 5�E�[̽��q��S����s͜�7�>�M����]k�F�a�CivGL{�/8auH���^��/o�ds`�ө�;=��< Z��T$��s2���,�v�+�錝��'��2�ա|S:��UrH�[1º?��=zW����g+C]���_ZHR֕�Й���uX��=G։�A�04���W�R�ӯⶏpR�X'D�F��tٲ��y�Ms"*u�v���b��@D7ZQ�©��rh=a�F��'[�µt�y�*�f����oǭ�{�F۟| :�0%Lߞ��U�ه0)Q&��bƀ���iL�E���9��,-�y:P�Թ:�o��6�����\D��^���z"�����-rO�ɛ��ع�������'և�
�(�$`0�UI�'c�T�WOU�s����1�wU�W�`�D��bhP��HuCMNKl�M�#�GRJP�����	�S;O��b�ݛ���v��=F�=�����x�g>�v��w_�P)cc��
��(�/f}V�M,��=;�M�����D���2�d�q�*st| �m�c�j���j�[�>������{�4T�<�æ������&)c�m��'KE#����(:���VX�����i��̫v�J� J��f>�J����}i>1{�}<�A�-�&z�W.�>�f���t��q�Ϻ��_yM^*�9�v	�j�a���M�>��P���b���е���L]Ig��E¼I�)�"�K�ED�+MfL��k'�����muP�OAu���ȱᯒ�Ykۼ�����Ž}K�tL)�������P���v�L�g�=n(F�X�(6�Զ ���4�&�<���<�a*���hb�N#Y�B��z����/�i���|����>J[���|m��uv�N��-O��	Jl�Zt8��I
��/[r���]�J�ڎ�ܙ*�1��iP(l]�_��|��p��.��h�|��������q�4	���ha|<Zų�1,d2�A/�e�x:s;9���E�7hq�$�*�ܫ�Ѹ�9��C-�z��F�by��X������)��ں����Z2���w�|	wH���-�~�'�XP��c��ޜ_�X>g�%;��c9��H$���V}X��
��7��F��"I�|5^�8uhLc�P���>߀��eX�m�-��ɖ��d������K��t����`��qZ��T�2X4��	,��G�W-n���.�����7.�U�kV�c	0�e�ݮ���t2�%��B�:�~P�l��ٴ�?k�����P(�8���p��î�A��GD���um@��I�;�Fx3eT��C.�n�zֲة�t�f�vKJ\x�ů-�ϙ�X���;��ɰ�y��>by
�%]SphZU��r�����w�ķg$�ҙ�2�M�C�8՗�5�\��T���� �
ì�ڲ��~��Fŷ$=���5����S�#�j�E1�PU �V���S����3�攲\�[j���)�;���9/��{��u���x'ґ0+���3aUznh�-I~�����|'c�0�:|r�آ�W�7��y	����)0R�d�8�C��ڷ��=�n�॒=�;Pfm�ޝl�r���8�#\��e��e<�kl��vu/�eS:HT�9�!��y�c�wX��T/���e�%r�l�,e%M�<d�<����-Sku�	w���p(k�=��&��S���>�
�����!z�d�wo�wE�"��[�����k�� �����Ǯ-h933_b�4jI�o:Ox� �y�+�b�vv��P.��T��R�iY�
��c0A����O1�gEQ���@�h:�0.m�e=SS�f{G}���OQm˖�Q~�S��k�u�J⩎��'O\ItPz�������Ȯ��#xF���Ώ��R�b<�g�$ƣy�U��i�M�`��3��	�I�a����3�����d�/��'�FsK�ia�9�1�-4�5��P�״Kx�R[���H7dx+��wdG�:�J[I���q�������3J�aw��m6���}+�50Ec�Ƈ�3�kh:��Uh���%��3Bݺ^���f���
�0�6���9���X��)��"��]�����9#���R�&����H-�����Q&�"?A�)5r@������J��B9���Ds��f�p%���9���q.���5_�,��m>se��7�H�}/��?\u<!v40d0)1��������A��_�(�""B��f�X&����Ǌ����Z�����Ӥ=���gǪ��~W��ʩ5�js�g���\\����))��e��T�jUEJPu�f,/ +�r�� �p���1��*/���H���C"�	y�C7A��V�)�!8�#4��_iQH"�Pi�jy��Q�^�����` ��o���V��ɚ��dj�S,��}"��=P�����ע�e�����Wyq�I �~=Ͳ�Q�}���e?I��Hgt�W��J�<0��H���C�Ca����N
�Q��W�YVb��h�>l���U����D�������K��|�A���	m��dD{����
x���"�z�3�1#�>�j�Z��:�ش����,��լ�o�~*�X�����:5���{f�L�4s��d���<�+��Yď!�0��~�(��J�z���澆D�ٳ��e�����`�D�譠�pJ{�g뀍>^�QW���dF%��fCl�����j��KR�+F��D�ҙwy]��c�2̐)8K6{��^����;K��?�ϐ�2̏Z@�����q�IM0%q�-���$��]D�����Ɨ���T/��)$��ʴ��2쩴���D�)��ؓ���{7�붃�S��7�=+��|/Ոu�,�Z`�k(~��Ƿ�4r��X	�ٙ�J\�S�"�Z���×���t�"�1!��4�&����z�6�����sN͐࣫�=��1ΰ�F���ZYˁ)?���7��U^l`�M�+w)QU���ǘt�
.�gD�I$g3g�L��6�ŤBiU1�O���<VU��vL�r�����کg�బ�-��Ҏ���z��?�[5�n���alqL1^��pg��K���t� a%5>Z��zv#�k�X�O��iqB��8�.OK����~_�+�v���L�7���\�6����i6B��Gd+�3X�'�ϣ�L,���V�����FX�u��r���S`�������+Sd�9��Z�l��(�`p�xbG	��<�Z��k��ِ)ś�^�]��,�{����0U��(�Q V����WG67<�� �?��ϓGO����ݲ��$z򻃘��Cn!�B����Kcw1�h�Z�n�'�0B������E2Vj��4)Z�0 {Q�@z�USr�g��B�׏��C�q fJ�|�Vk�=�Q0��	r��z__��u!��ӯ]]��2v\M�B˳iO�����̨i_P���}������@��2�שbKϧh�u<�pO9>��T�G���E'̼%�?�"
�����i���3����l��!��`�2u�h��UFe�3��g�e�M L�ILY�㖒��-�0��J�ȍ�f�ub�Í tc�hfp�a֬��K�1*,U�< �a�&�i���"�F�����,���m�QC*���%����a�}�<M��Q��(.�����Q	0�9n�*��0Ǔ�5Ԏ
�h]�X��~�^�O٢��o�qW�:���I� �{�X�-3N��ED�B�d��}���OH2��Ny\UM���?�#��4�%��(X2v����!ܕ�\���h*H��	L��2'7`��S������M+�@e�dSU�����y)�n�T �c�֫}ש>er�QB,t�Z #����4��d�lך���Ӵ|�⮮����$ՙ�p�v��NAt�IG�T�j;4ؤ�
Zk�<�c&~ңIp�DM@q��;���uP>�`L �]��H��C�~U��"+a��$<����k��pGX��~%`�@����B��.�c8�� ]'bG�2F�ޓq�;�en�M�D�Jk�ſ��3!�6ö�{b��� �����Tl�p�t�D��~��g��,B���q-hh��>�+��G�.��^���7?�/�5�XS�_�4K����޾��C��bfj|�OM~m�$��9/(��,�C�z+׫�~��.��p��E�[��*��Wu(AQ��[��sόW�E�T���J�-O֮V�����bŀX�luc�1W�z�v����N4��!~9�f��D��sԑefs��OP���xW��(g���݀�HՑ��/�+.�9�5�Ga��9��X�_q`3��Nh�~Y>����C۔+M�%����۳��b���������R��<r�S��c!R�v�˨��u&����{�T��V"fPx�Z�C"^��L�;꬐��/��T[I�3ЌdnꎉҾ�p�cq�:��_aku`�X�4��cR�y5f��(�2��z������S�{6��o��o�}<ꏥex��\��o�'��2e�Z�cS;!��c!$��~QQA���H藗��5	Eʗ;��ī�QR!1jΒ��a>���^���s*��,�z
j��8�̉u�5�+_[��9m2�~~�e�*��zCϗ�+:q��j�r��m17�o_T�BBo��mv}ި����ؓ��<�Y�F��%�(m�3��u�=�G���Ȧ!{�z�t�IϺ3�_$���3g�P��a'��@V�1<u�17ɄUh+5Gӂ�6�� ;���d�؅��(��zeɍZ[]����;�ۣ5��8
o��+B������qw�nidKځi\yvL,�~g��v�c7�^C�B �߽6s]h�n��`���[hƜ�wpP\~����M��g���jɇ���e����9S1���W�> ۾Ř�k��Ʇ�0`��ř��.�^����l�pЖ�>>����ͩo��5����Ӟ����y���M��a��+�;HH��t�8�r��o�_��[�U����������E���enn�>r�u��d���u�a��zec���X��|�˲+�fx�ZC��3�������><Z��ꮅdRJu�h���u�]���������L�B%P�S�zc��@���櫄��E@}a3�����`F\�����!���`b��n�ZG�<��I٩�Qg�� ���ڬ��m�D%{x��I��Q�h��N��H8hi-&��� .���d�f�A����mWAĔr/4B�Kc.a�}`�2̦F��,�� >��X��
���1��~s�h-7B����ڤa#���=n.:��c��a���E�qZ��d�K.�K	n�b�bŃ���U
?�X$�q	|u-JHQ(��&o�g�t���S��<)�ґ�_�������q����7�Y[��~	�b.#�	�e�z�J��K�i(��+K���e5[3����
�~��v$tڃ��2�d�|V+Ź�L;b�=2�!�w�m6�߼g��ɀ8+��b�'-�R�Ȳybn�֨�(Y��eL�nxz@=>��>R����)���"�{�+����9h��6M�M����g�ԓ�f�'�PW���{ :g��<r7
�$V��g��K��P�{6���bm
�4����t]���j���u$%��AY\�AY�u�,����jc��j��O̤��m������P*�s�]L����S&��$�c�$X��Ѩi�����n�k��h�c�h��C��l$n,�,�T��CFY<<���l�\�.�jOi8G����r�*s��	�˺W6'��/\���im��ksHe�Lދ�wb��������t�|}ߢ�3}��^��!(�B�q,ɖt�I��8Z�]��y�<57@��
#�͋��8��kY�ͫV���;��ՠO�u)>��$�푯��N�ق�u�d��MX��A����(z&=p�-�8@⛍��Qomę�n8$��ĸ�b�P,G�&��1���#���a|'��dL�ѳ��UPؗPb#Tng��+�d���f�~	�+���s�Y��)�g�6�5j����ި_�����������tR��V����7�ו�z��7�$6�7��"MK5;���M&�b<Bߍ8��FI���xa��L���A@\�v�.&��9���ݬB��uù',�<y�9�Hݚ����A5N/1��A^[L��H�Jf/x��#�7 �y�&��La�9-{�<����.���/��� ��e��<�ϓ�$qe��ok����sUz(
H�^��?2 AS|��(���4=ǲO�r�f����0\	"��F3��<�<ޖ:�I��_e~a�q*o�ek7G@���$מ��[�tv���e	�7�H"��õs6��M>��x��;1Ocu�A�q�L?�ۥ��T�}�f])({d��؝/1��bʖk���u�d���T,���d�|=3n�ߍ+䉮 �~�𷾞A��Ft_{�ӽ=���O���8����n�'���)�ͣI���0�s7�$3Jz8.sb�>t��O$f�N����-.��њ�%#�h��O���y���,��ڶ>�����x!�3�V/�
8���ҝ$�;����5_���O{! �Ml3U��2��B�㫽 ��L�1�G�<�Ŋ�:�h�&`�7n?9��5 �/��L��A�1yA\*9��X�6��=f�����9 ��/�ͻ�:X>���Z���_�����vg)Qio������I�Cp6�w�4�����~�gg��}3!��_�m��Z�m��<Pj�L���<��a���솝\�]_o3�����+j��>�4��9�G��m���qu�)�SN�SJ��q=�_A��IT�q�7G�P��]~-$r���� T �����;0��?����ʰ�8w�A�K�,VŸ��IbX_9� Y&{&zM���e�mp$H��9[I�w���u�|�A>V�/Й�ۯG��2UM,|��4\�h�RN�~�c�ێ�W�{Z�2��ut @��XH�,6�Y�ػA�@�M�L�H���ʦ\���#V�O�3nw����}ҡ�-2狏���#��/s�f�(�)@��f�������S1��H�uO{�6���oP�ZJvQ���`ϳ���ԆFkm���@���\��X�	)���{�,^�ޟv�[�؈�Z�Iѻ��%��R���%�
θW*�p���g���"Pɥ��M�[K'j�U���o=S=�:�̚���V���5�b��je�I����}�Y��!��0ȯƦ�;OJ6/SU�����b�4*P%{���3���O-�q:���(��ӊ>A����F�ɏ�ϖ��+�&U3_������'�cWߙ��hU�덴��B�����>���S���ܺ�vJ�@�6E�E�81E��w�K���N��|�h_@��K�./� �ٺ0���_��iͮ��&=��`@d�?�P,S˽`(XK����5���A��gBy�(	�y�
\C�o��('��r�����S>��m��g�~ ��E�i��\�����!�������| ��%�. �[���ϳ����oQIn������@��ʙ���`F`Zɞ�j�A��z�Ǥ�ըN/DI��n��,k���o�}�������mb�Ì��#�u�z��w�K6cwl5ڵ�,:����&�C�}�Xյ��J�"MW�N=�]le�v�����L-sr-�m�v�#i��B���ˢ�X>�ǅ�!�MZ��{v�����u;�\��P���x����Z
���~�쭉�h�毐y�����3����qϘ:�i��Q�����U�߹��xį}ލUn��� {P��C�ά�wgA���J��:��c����h�o9�S ��@�N�	�*�f?1�N�\WXu�
㻃�WB��	���O�1��y���@����L��V?D�N�ƭSi��9R�1C'�T�*H��ϥ2�/����/�XREg���'��}�J��y���r&������O�z���(/Rk�ak^�"�{���Cqo��)�FbMWhM�K���]Z}��-�0.�w�\�s�NP�K��Ũ�lFK1�p1��UpPF�ƭ�8��i��^�(+����cv���&ķ�����U@�{����1bm�g�þUKM���f�],���O�w;�
.��;%�28�1�"��i��*�6���ܡE1nU��-��y�DY�L#1�n�ۙG=LK2{����NJ����.� ���ݼ��o���&7G� 8�;�.���>�P�J�Z%�O���6PH�5��W
�^CoD���� ��!3��Eê4����,����(��J;�J���D�f�M�QT�r���kP\o�ԣ|�xq-�7�@}�5���H�sK�Z��b���g�:��G٭�.h ����"z�LIMu�#��ܦ��p5����nB+M=����>�5$}8R��L�H䀐�w����@�ȳ4iJ ��.�W�^�����Ak#
H��<N"�t�>IM�;�Yy�goF���fYO�e�7�4�!S�S��.(���㲷��s�s7Z91�5�\m9ꎩH��}L�s�K�#Jũ�����(�p��(�܋ԟ�ɚ$�6�FC���_��b丅�i
�=ѭ�F>�i��KU���������yj@�| )m�����w����+��2�W.�0��� n��Bb<��M��w��;���e6���m�o`��s����Q=�ئ�j�n��CjZ��)nkN����3R�0�7$��Rd\��a�v�B��IjUNۦ�m�IC�,F�J���`ҏ���4��l�ǝ��9OgU�D�n�zN����� �*�P�O^��0S7�Q�^aԙ�͜ɇ��EÜ,�s��$)7��S~�"���&����>"p����[��u�Y�T��m�5�똦�+j��4��@O�4�^���T|�b�]��9�ƣҳNl<!�	�'�S�=]n��)Hp�	
�W�=�DJ	Q�I��!;�@4�$ ��^�2������󠍵�a�3�f��{��3���0o�s�;��v����:�TϺ�7Tp`>Erlj���S�-~a+S][rἯ:�L�5�m����V=�5��qKn|:	b��N�%���+�n������2�H�4l���CZu��r�E�����UPU�-�+Ǎn�ƃ�q�GCd�}�
��C��,�Ӌ:K�o;Qt�Ђ���j�ɫ֤�B�?�~�|3����Ȧ����L��H>�L��t���~�H�il��X��g@��e���0r�a�f書�
��|��A!���	�r G�*�b���K�>5r+�	lz�J�!-#4	{����rw�(~<k+G����'uX~����*������F�W�g.�
�y��Oꈬ�?ۋS�P#;u�yM��k.)c?�U��.H>�B�);y���a�ˢ }�K���|%1kCgv�ǐ��:�
��o�}P"����xi�~��'���%�cU���ņw��-+���긩a�O\�ch��Ƴc�c�lS�yy��`��ly�� z|�*㮳���/yO!�'RG�wEPu$(]=��P�B�����GD�-J�5���M��������_����-��ß������d0B����CaU�g@ ��^?,��<p�3���h��ߺ��a�χ����`~�2�	�ć�]�hMG��P
@Y�&P�R�]G��O\Y�aT�{'��n���r��P����
\#�q��>'Y�wm��߭ӛh����LޜB��^֒`fh[U�P$�z�Z����[��:"�X���åH�?>�cr�A"~�����
�
�Ώh�M��պ� :��KbW�{�k)
T�����<�5���H�~!j�\�3:[#���0[��q�^p�;�#N���B�|O�,5�<5!��6�-r�5���=:W�F��0~tim�$��63�D��E}t��s�Xܶ��r�gX ��EF"g��+8���� �-���O�;�6�R7�J
񭔺�(�H�\fw'�7Z&�	��@J��� 0�wqy���o�U{�CW�D�(��"
y,<A�6���6���t�;��e�nw���։��Nf����ɔ�ĵ��r��#a<��i9�8ٿ:^Q6��y��s@�c�r�U7����LO�Gf6�����
��<��.�z��x_���=��k����-�]�f�8�7�*�'ϥLg�#1���{��G�`D�Zl1Y�̭]\c�����~}-^����2F�fxS��Fc��ڮ���J���ź�X�A�ư ��:�D�B���G���xw����v�*���պl
|�x-�D�<V���L����:肏��|��´瑩m�[�<�����*�m�\�i0�/���jC���u���ڔ��N8I���Z�:��ȾF�y&�'����Ѹ���5O~�����J�:�{�n�N/ʍ�_���^�B'��"�TR�����x:��5��b	l$�w��P�x������$#̵�v�d\~ٻak�����O�G]WF�~?[���ޣ�n�B�#�w��� �JW��#��v���+V�L ����W[e��mU��:��O�\m<a�?��jud�"�*ℤ@�h�Pe��s��F<���V�??�w�D��d!�o���#���{XY-�NH�0�C�.;4a�A�"}8Z
�T6�-K�N�V�an�}{��q -K������J�@��1(�~\��I���K/bEȻ�ʭ��yC|�#���Y�\����IS>���٨�gW�T�Ϻl?���-bQjhZd�yE�Y�5Y�U]�=zXK��V��q'�B|���zp�^u��(�N�D*��nIȾH4�%�hgB��g�7����� ٝ3ame���m��/h(��ɍL�i �aZ|���HR�_���d~"gqn� �f^����	���� ��M^5��	��!d���b-����Lr��ɬ'TK��ڔ����xS;���Dz	� {W/�C3�#�C��DQk&m�q��������/5�S5a` �
�?���q2���h�T�Y�1ӏ����V�K�Xd�Ӳ�[ލ�A����}n�Q��9��\
��j�r��lV��)�9�E�b4�XbѴ�%�8�d�cpt@��E.V�*�L\������w�_��q`T7?Z={Q���������V:NvJZ�H�/�4������:��Ʒi���셁倆��n|,G�1��G��ewS�IR��1�풯g܍𤽎�����ˁ��¯�wG�W�B��b��
��W��	PP{��is<HDβ���ԯ�3�x��I'��szOu�I׹P&r���m�EN�}�i|A�bo0�l�s���x_C�6�ٚX~��s�H��ޢ�@%�JZl�)��0+A��~���Z&��!>��
�����0kd�/D��<�׃��m�ϱ�����B(#v��wT�u���9b�{l
����"@��0�;��9�_=�L�R?�}����RY��.*�p�Z�
�>ғ��G�?:��5vs���,	��ʉ���U�=y�^�*�D����C�rv�]H�.�_|�֚jgjn!�HD�*�j��L��E}my!����/bm�}]/ן
��i�P����H���5��NKd>�:�=��L�O+qA�a���]�B�[ ��J�Wг����_:�NV�hbg����R͈7�d2��*e4��g��epQ>H��U�a�Bo�,k͝QE�B�y�!��%�\"��$P`�I>;�$㕇���D��k���~� &�m!���c�avF���(:y��d���È^�xx.�s��5PXЫѴX}!�������V���'zf?�v�S`U��?�Е�?���x�a0�	,fI���qQ-��QhST'�AZ�L*�}��&y��x��,�Qk{�W��(9� e=�\"F��Iiפ�((�?ЅH���e�	K/���J�E��EeS�f�7���!&�Di�K�T��Cz8xI�V����n+�����\~a�����;�Aaɓ�״m���Y(!O���y}��]u<�5K���O�<�u9ZB��>9�����Ǎ^6�8�Ru7�� 7u��AX+4"{���.xJ��w�]C+Aɻ] �JE�{n]M#9�-��"��a3qDU�[�hR��Ƥ���E1 52k�Z���
�gk��&i*w�������T���R�T/������@�~�w��Gu�ԏ���Zm�b�*d�X��v$M�՗���� �z%���DRﻥ���ыV���_I1�3耐�*j��̇)J��'phJo��:��:��dk�x�*QO�'d�f�|},)��f=�kT�e6-� o�[���.�D���L2AF�@^��Yr���6�X,;��5����w3��,Ut�a�LC�~/a���i"��.��H�-a}��ʛE-B0j���}B��};���#z-\t�y3�:2�
��A��%m����A��'��d}�˂G2���E�$�)�K���LAM����Z���;L����_��݋N�g*��?5ٵ�kIAM9����[Mmؓ��e���9r��K��ϧw U�&n���b:+$�s8$%�&6[��-�C�ڶ �W��lH3���W�j�-�wh�k���h�\�Tk�\��=3B��|;�BE��Qސ>W��F�`eO��]�iQ+��e�}�����@*�.w`���N�!�n�?��Aʍ��.G�t��QH��y"���q����� �(_CR�^#�!C̈́�j���$�݁���8�!+���@U�{7�����.�&#���*�=2v�\�,w���q�V��9�8i�IGH��A�]!��X�ԉl�nC�.��Ĉ#�dfX�]w�\$����7&3v�k�vS�����Ⱦ,�z1ε6i8{�>^���y������r	�CX�]�٬��\�c5�,��Qq�U��\�O_6�_a�����YDw�e�l��$p��:�E(g.h�9p�	�ϛ���	ͪ�O�l����_x�B���@��j+G6{[HQp���@u�����r5u�D�5��;Hgʒ�x�ˠӦEATƍP3By�Od�&��3�A~��/�j&g�m�b��!!}�(�4��%g	_A�{�����ygSաr�WQNQW;X�OX���<�x9	;u%dmiM~�u-@!*��g�����/�.�'�[z�Y���Et��+�\�Y��s��/�*e��OV�:����{$�I=��K;!�����O��"�Ku⧔�A�^
-L-Zt>��^j�:� ;��Yg2QXX�.]eRA��0���4��K�et��;$�)�=���=�C�E$���׮���b��W�)U�p�F�0��H��R��j-� ��������*�L S��LU+�q�O�19��FS/_�����5�il�����ֆ�,��'���`��BaŚ�8
�~�]��ݒ@L�<TQ��;{�d��QFk+�t��)%�$3]^:�&�f����HQ���h�)V�I�<
I=4da��ۥ��&SA�-�\� ����K�b���pf�Vu�+�b�s
�7b׺���=R6dc}�?�|�X������Gҙ�����|�B��s2����to���^ڄ:�� 7TB�[X��c�B�\�����3��j���m�Aw��v�G��[�B�_���%�T�0`c���)�W�������J\���5U�*�-_Ǣ@m�����{� �/l�>(�����,�Շ�����m�V��*�~��^��W�����5�W�û� 35Y��oJ�H�������dV�ŷ����������E���~�U�����6��)(N;@�/Y0�}a`���3�P^
���EO��_qH����|�Y���SO� �'���lh��J5m�^�á�i���������{\	n�t�C�*��E�4�%O,)5�ݟ��2�(ir"*�J-�=h��YP�2�W=C��Ê%��J�"��PO�N�SjUw��23��H��.�(k`��|����6���}k�X\^��w��e(i��gS�Y��K�!ԓ�&E�E����σd�-M7��sZ�|��x�]���L��v���f�<�����F`9���cW1=��7��	��W85��>�ׄ'���"4�m(���Y�{�6	c��ljyi-�p�tr�T(���6*�Ws���(˪��A(͵U�;�;�6/Aԏz�`�Q�eC��Y���Z�^��u��g��J?)v�Td�T�sGU�G/�@{.��5ݷS�vH����H6Ypw->T������L��J��K�����[�3�ڻi��K�
�,�`�<�Տª47�@6x~�&W&��`���~%�P;�}������@M�����iɨ9z�X�P�{rX���:�Z�J���Oa͟q�B�&_%\����=#�F�:����i�H@I��U� �r�n��ڰ��폓�]="O���
߬Gq7��>�@�g��M�8��� ��Z�ߣ��ߝO���s�T#���FpRY���7��M\:-<R��\|�ܟ���V���`�N�\�8�Tȯ��;Ѓ*�i�
�#q����)�I�c��p�����s:�+��,��oƈ��?}��	�ͮ�([�������7������^�o�-U!	��Q��:�]�%;���o�ʫH��o`~�ƶlIt�LOjJ����{L�y������hI��Y�e�m�^GS�.Xw�չa3�<x�+�+|��`G�Oҿ�I���V�9L�lq�i�N����cO�
W
�VW8��{g�ؕ�l�_̞�e;Im���)}H�ZZ\L�sz��C���V�����n��%[���7(�Z�A!��g���X1��1�
��{��D����ҺGDk�/N+��>.A ��y�Z�Ӣ��R������A�I�����D<
R��wϚ�+:H�	.�xFY��/1�Ѩ���Cgx�����|�����s �dOS��r٪h��_�+�Gmcq'�1}�)'z�t��K��&N��/��5���]b$�*�RfGmjմ�WsxcZ]7*1H�u�ԩ�m0���#��ɽA��&�^_J.|�%o�V���
U��M�`Ǚ�X\����yK'��|o�ҩ�x�zM!N���Z�E����i�a6�2���XS��T92T��5,S��S}�X�a�?[{pa ��}��a��&|���9g&�Q�A>y�%}�����$J~Ôh�P_˕�s#QN�� 5�h7�2TC�#�I6�Z ����B.�yi��8]u/�Rui^c t���򙩗;r츍)�ⳤ��\#�|�@o���ٹTic��a��wf�Q��
u���K��3�G��g��FVkJؕ$������J�}�uĎ���DY���u+��~2�W��������X����y�,��X��H�I�tx�a��U�&`���M���@�k���1f���!k����YҮC�ˣR�[}C��v9��WN���4xn4D�KW�����=�v�Í?��燩�l�S��h�*'�G�5�^��9�x��P�m�G���[�QE��D�=Q'��G��r���H��5jڞ�]�5*TĂ�Y�;7�����4ض���iI���? �w+<?qϒ��%^�<����7qd?A.օѲs���[����Ǩ�t��`D��(���K��Z�|�Z�:�O��ܫ�*�i������s���9!$J]�w0��_�,#�eɃh�)�eq�	�|%�ZQ��Qߋr&Z�5�	�q�w�^ݓ�D�F��&�����y�V�1!f����9��gWҩ1�@�xsc���q��W��^���8�����j�A�Lm&d�NIl���|ٟ�{�\�c�"C E?��~ٮ�dEV�`[��Jg����I�A�)Y�>L#e��̓��d�	���@7h���֖�9xs~�|@9�3�$!jd�ÓT��t�����ěr��_���9�a�[��l�~o=ѠQ�n+*4q����b�ll��P
���׵�>�$(�c���c ��nv���K���́r�מV���Q8M2�I¬V�mMl*d͂XK���oy�WR�_ ��k�eJE�����[�N� ������{��Q�?y>p#l�O����}f�J�^n?�F�%�T���+f]:��O��tL)�x_L����.�Y�p9ȋ�n��'�H^7Ń�L���iZ	�A�yIu� ^�ͱ��M��$�����[���6�:�U�L�m���L�ɻK�S�^:�͉ma�V�l+��Z{ �����I�(��Nѓ�^a��[�UX	�{���LE�`vE�:Q�$@Ͷ1=E�=v�$(�p�ܲ���_r�f�O�/�el�ϒ̪!aw,��y��^�@#e�	 �����)���G��+O�O�l�m8H٧d V'sxW=%�i����Ԡ��[R�)	u�8yVg?dq|���i?Gh��eTW�?Z�Zq&N���`�T���"�\��
�b����<�佟Cc�)��D4 3�R+��U�����;H��p���;^H{<�v�5����P�)�B2v�l��Q���:p��5�r�M�7dj�����g�n�,lfd�bs����7HCpQn0����9��C�{VX+�3;�U��$P��4��Φ��w{�cD��'T!Z�Xx��b),�ˊ� I6� TXJ53P.������f�9��0v��C��̰�R�]���oX��k���Dil+42F8P�[��C�*?	�F�Y\B1&k1�"RE���ǥ��m�v�����ϻ����.�=y�j�.^t �d}��u��|�TM�,�ORiZQ���"��r���������q���"������L�O,`w���k�i~UB[��͕��T�Sk�&jqz���Z����ע%l�cvj��y��������V�h*�gvSa\+i&��o�Tw8(�Ջ�*X�T��0N5.�<[k��IP���5���-�϶�|�$���.�����M�k�a����C�5*,�c��.0����gy���I��	�ves���k,�:�PV�Զ�-*��;����0�C��a|�H����y\��C��K�z� !�9����i"�3�3lXo�⤥����l	��K��,���vU��N�lOL��?��u��ٔh�gD�m׽|�"t�)�O������/<�J�)r �S�^��
M�ک���`��H]c�U�J�����i�9-����S�t���1 ����N�(�O�Q�"5�1��Yo�N�P���Ĭ�V���m>2�TE��6�:����yE�E�j�de�:���5��B-�4�kI0�=1"��ʺzۛ�<�=��>�ӝ���W��.�m\�奛y�
�%�q m�a�0��%ϭ?����~����X=�r�x�����$�%o��]��t+��n�*�e�܃(N�%�揄���G0�%O<�y���+	N~�; �;ai-��Ql����b��)�~C����{�)ꆞW7a��r_��%��e�����"�Qɲmݮ��a���#�>��3��G�3���N�m@C��	�o�D�C�?�JjpR��X�G�.eg��l���G0��r���iKEu=^sVܪ똛�(�M	��Mҗ6t����Hl�g_�Um27�s�j]�l�#�Ń��Uy&����>u辗����ާjskn�lM/��s���	-��L�$}���ܠ��G溪�U=ǳC�~e?��ok~���t`Tu)��_����3�����Z�=<W��iSc�I�J!�fd����5*�X*l���	��Ȃ��ܳ7�0 �� |�*�v�y��D��;P�N�Цi���lQ�-6-U�ab�O^߄�%r����>*r��s�"�n����8})�K,y�`�=���@�7u�����2"=��
W���D
�D�?}�&���� s�nk����LW�1Z ]HT�o�0��# �]��l�O;*�mz�5�
t���ԗ>�Cl��he �Hb#�+�Y
vˇ28#Y�mo�����Qu[��A4��'�y�MY�by�A���f=�)s�@��;S�D,{�
ℭ�sh�W����nrjy5���g��$;F�+O,��-�~�����ϲ�ѹwf�1T��c��t+�=VAĞ�c�x�� �e��@q�:-!H����CIT"M�͵�c��P�!ЗI�_��Gwp�K���uAȷ]d0�XX��]Ɗ��z�-�'�{A$i�?��5r��s�j$��x��3�Vt5㋺�����x`���8�����4փ��"'Mұ�7�h�Ws�ܪ���]�Cm8�L����|���ȥ�o=�i�����7�6�LUu��E�2���@�|e���B��_�sP�B���@U�\g�Ƌ��&讙����WLF\ׄ�?�Cy?��t��Q_��8�h�'��^c�V��H�|���7�3g�R}�~��5�:t��cun��8"� �K��?��O� 񂅤 �����Z���s(�����hO6� ^�"�t���Y2�c����V�'�B��nVr6����m3n��Og(��oY��5��'���߲�Ѧ>�W[�Fu�L-ؕ&���,|bN:u�
�Qˎ ��u�FbA�M�:|��3<XS���J*F9���DP��@�$�iȭ��֞}-���2� �"ߟQk�S�1�u��xe��ߦ:��9~ ���9���1�-�>6E-F�5�'��^V�Ie��<�����������q�v�]��Y3a��4��/�J������{��lL	?c�6ŵ�����\�N}�d���55�p��p��^/ةiGF����c��j�D��H�"0�?\�@N~���jVq��g(.�Pݨ�4aj~}�W~n5����<柚3��T�m*q����9�^ʨ_��U��8�x*(�-&y$s�A�-���J����A;W�@RVjFh_��Y�>�$E�L���/����w+)^Y�u5��Zx���}fT�3�^�#�O��q��M�M��I��/Z�y^J<-�EV]piY:|*�p۹n
b��K���8�>t�N��N�Ypi�(����hGCF;��a,�ЩjrC	=G>˷I|�b=��� ������� PFǂ��-N��#3��Jo�	t&��2��ˊt�o���	!�©n*��)��2�F�K��� �G�q1��Y呈u���tG��qE�7��^u��m,���ɔ��MI�Y�4X�H���������wt�K&���sc��jHW�jy�\Q^ p6�ls^ޥx~qP���RI���b�mg�m��]�K)��n)&�+9�KJ(�iay���i�*�o h=�K�V���  ��v	�H�A>8}�]'.�8KoNh�3��bV�d��Q�O�ڛ�;���)��;J�s�ZO��}�C!�`�#;m�u^�dz�Vc�1�:�<@(��M�p��DW�AP��������m��r�`�97!m>/X��y�uVn�]^#jI > �F؈9~ľ<�a�U���3$PC�;��7�En�6
#�-JF=^՞�J��f���g��Qm�]w2��_ �9��96��w7�4d�\�	�A�R����N+�;4lPm0Š�]�tú^*����T�8_�,6ܝ��R2���*h���П�0-*����.r�:�S��$�>�M{�M��&��W����6@Uj.��k��ėcӤ0��	!zXL���WW��c-VI騕\�XI��$�iwn�h2
pK�����Uj/k�H,�Y��������Y<�1��BT��l��ak���p
�7*	��,pK�njxo��+;�J�*�� ݈�iAW��9�H��(K�,E'����Ƿ��F|�,�vl�0'�w%��
�^O�*�8��B?��rRl��(�m\#w5�7Ý�P�~ �9ŤL ���~L�#H�ϮN�W��"���î�&O�k���ɏu�,	����>k��!�[k�����E��ЌNJ� %G�v���F�d15�u�&Uz�=$��|0�!�)�)�0{	�y:�%� ��)|���m�ĪX�Z��k�F�z����:)��E�5���7 ݂�{�zk[��Sji�d�Φ���+��/�����r��A�;]Ӧ��ѝ��w���B[W���3��C�P�3;�T�Mi$�b��SBrS5�B���� �Xkw|TUD��?��Z�g}P�����1����>_ �PS�g(��Y?�2�FcUY���m-�X�2�C�pK���9A&��Qm��$>j����-�kW5w���z#��LM{L�H����L��y`�6X���|��Y���+�����e@/�:�x,vj���f���?f�٫|v�%�]�=&o�9��֡�k�`���F����bX��D9�!k�7�xn2_�\���td�F�9 ���]�H��)h��Pdpv+^Ugd���m�rO��D�@�1�(Z��	��a��a���d\���5�����\ c��J�$�6tYB�����u�~���L�H�%����)�Ӓ�=��IE�П,���o]����֛����ٹ	k�&
*�0�m��-GRl>��_$�V���'�-W����%]\�u�qMA�7 Q\G��X���@D���.�����&A�q11��&Hù��X���	�m{��i�#)'V��f�.\��@�>����-H��t_{�ʒ���R/�4���T ^��Q�"��&m�KwF��f~Nt��pUAw�Ϛh�œE�?��`���5g[����F����!�`�&��G1�E��s���0�*6?�����fÃw��Z�
:����^kv�oy��&[�����`D�l�ˑ� ��b�7�>ĩdym�|�P�'�z��هZ1�ܔ�p���@u�|+��>; ����~��~�[U(�9��T���A�ݐ�Em�:W�����y1✹�t
��J$�tH�
������o�u
�/=hz!��j[���g��$l�y�pu8o"�<�=[�,c��NhvZ�w6���t�� Nϻ���w���&�jC/5�e�&�z��k�r�C`D��-D
�WOM��z[�f���Ppw9Z��/�
�!h���J�ɕ���m�g�5;�Pd>������}��ND�gd�- ���R{�I�ȹ� X3֍�����+��z2�\`����S�ɽHB�S3�<�'�P���鈈y����M��*Ő���;LD�6�l^y�$2Bb}Ĺ�9{���\d��ͯj4�`��\0"i���<��f�s��C'R���C>�fw�%(����s!��Q����7�t�4�o}�۝g|���gP�r�f�����3�-$ਤw��,�K����+,,�O߇N�܀A�p�6�
��`�Mx�����#X�A
��s�j�0��Y��==Nv-�dF�a��6�!.s2i�-��:)u=J�]'���U�v�e������c����H�z3����~R{��䗳��9 ����{�0�Yo��,��2y"l��)ֽ���-�Bw�*B����#���J�G���q�Ah��ǜ]qk�i�a,w���=������5u��^)4�[�vN���Z�WX^E,����,��=�����i�v��ѓ�f����3D�L�I�x�#�`��d-W�ٜ�9Q��R���8�e�*�&��@��2�1]�4�ʤ����}�w�u�]:�o����ϑh���#��d�6|ww/���ʱa"��cs�RԐ����$�X�+f�Y^��X+����G�N3S�[��;����3�8�O������-J�'R�ӽ:=��	�j��*X^2�:�zO��J�m��wӾDL��WM�uՎl{s�:���|��%F���}9��=��|{��e�o�]�B��$]qA>ظ:��p�h�|y�ާ/܏��X��N�H����xy������'M�ys��UA��	F�V�5HO�)1� ��?���٫a�P��ίޠW+c�H���>\��P~г�y ~6���������a�W�RLcM��<��gj�:��R���$�����xݣy;�,ÛE�\�l��
+�	]�*��i�=xOD�0�.���r�x�D��zQ> ��ɮ��YQ6���'�hz�l��T�kh�g�\^���im�>�V��38Ԩ!���