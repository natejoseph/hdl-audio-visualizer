��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�9 �jAl, ﬷wT�����*�u�sbH�v�%Ih�h�M�f�K�I��G�����TM�d}y�����/���X�J�x�u�He�Aq�/-`/Ϧ��_!Ͷ��k�n��ޒ�0C����b=��Ha^��V�I^� R���JD8��/S$�����y�,8�/yaO�`��!VJ�m`��<Џ���T�]�7Kki7��ʖ�B��������o�@�q�2&:2�T�q�T�!Gl��kT�u�ʓ�q`%�����mT�9�RA��F��s�?���]���m#ʰ���P������r�/���>?�Wտ+<�m���3��?���b��(v{�3��г�*���V4�"j�8��w����Oc�������&U~_DԕBf�����w�S+��e�����3SdG�)=`L_ȁB_�i�T�{��)��`ęb،7��Y�wݑh���L��g�JL��r��=��-6
$�hR�
�Qee�ΣM��#���kT�D+�t�-�~
�I��H(���
�v�$`0���apqm���^�n�4<2�%��͸*�0;����^��ߨ�$� �*�061y�MUj���L���o�&�1��TI�-J��;�@4�2M ��89MCB�ʰ�H;|*ȅ��]�����>
��z6:#�/;���V�㟥$�X���f`��;�]�)ez���z�n.	
ZU6�̮g�Z�0�l�/��唄6�����KXD���)���5���q?��&�OX��^D۟,p�D`��������'=Wh�"j>c%�BS�S^�Nj
�g�wD)*f��L�LC�I:�K���_'K�B��!4�ŷ|�8O�10=mUFN��A��$ڹ ��j`��!Kr8�@�Kz`��V�
<u�4؁��l��p����5}jp���ޓ�c���р�n�ՏJ�� ��o�N��5KjbAc�:t�q��������W޳�ǌQ+��Km����<f���NŖ�h%��*yǁSYE�jpi���l�֢(}���:B,��$�\�I��@A5� �g�)F��F`�!n,C���K@�";��DG�x[��u�({Vi�xM3c!`Ei߫�yҰ�(�zp���G�S����ٶ�̳�qo޵�D_NF�2��׽L�L�Ҥ�B>/��� ��ۓ$g����Cu����~�ՇQ%��m����>����S�6�
4����Q�H�V].tޙ�櫧5�b�U2ʎ�20���Ã�u�R=.�����'~���HQBxu������� �	�{��旯X��G�e�']A�M6ɸ�ʸ�Rڜ�4-^N����I�>~r+��z�0��#�}�p�����Ս�T��lێ�KL��}��4���L���\%�@D�Á5Mp�@� �H�xx�h?vB��`�p��m�+g& �&'��mCu����4�f�b%�Pk[af��K�m��3{���}q �4W�
v�D!����>����#N\ࡶ{L�2Q�_�D�x�d0�á�m�HiE�ѡ3��߶v���&�6"����������F"3M~��V�����f�Fl��)�h%�CMh-�J�v��,�g��D�M��h�p׹ܾ��1�(R7f�%��XM�7d-Yg�cPm��T;���"9���޴\+FIb=N�%s{��Zm���|'ꅕd8�
:��\5��}�Bֈt�l`lBTp�u��#�l������ ���ÉJ#�W��_s��r��J���W�C���6v۵xrkE\�D��D�d��C��lѡ=u0٦��F]C������x/�.��i�\�����}��г��a�=��ia�]���Q�T����*璽��6��c\l_�l��"WӲ��c��ҥ�>B�2|�7��tE�?�Z�4�q1�A�Bղ�F�~?g�ҌM�7�/mr��S�����l��g��Z�U�Js�d�0J���L�N�ϫU�� 'V���e���?b����Ӿ�̫r�>˒����Y4G���~�e��E-��:�93�L4疸�7[�Դ?��O��G��25���F���*ِz�����F��ن�,�������֪.���t���Z'D�3{��E��(f�k��<!k�r0'&�)��4��;E�m�ɉ��F;Է1][51;F���(��7�a�O4߫��P�	���H����${$~��R!��Y.��ފ?��-И�G�I��rߔ�μ���@+�c�<��,����5-l���9y�gpߜ*�Ѯ 5�^=ӓWb���ٓ
y�\p��&�n�Y~
�Ѭ*��A��*�
"־�I��=�fD�p"��ah`���Qi�f��U�~��OocƼ_AyX��HCI<�,ַ�b�n;���W2��%�ra'^n�I�Mo���-Қ6'��Dq�$�sU�oc���y�z��P��W�#F���\y��c��@���ؙU/����A�T-���#O|`9��G�Xk��7x���w��}B��;���&�����lyAE��f)���x�:���Qs�PSF�����\A�W=�BHI��,E��Z?!�?��1����>��E=k��wh��ԥU�v�u�P��'��2iO,�i����?��Ӳq�	���<]�o@i$ڔFB��s�ڸ1|�.�;��AcƎh�C��GB�"���O�(m�=�Z�>��r2��7s�k.e��د�;������#쥐+����!yE��8��iZ�5�"^Cz����ɟ��Ee\�\U�\[AMTk���);4 .�����[�.�����5`��(�ww3��k��N�i�EqG�M`CS+|_0����8k�%����^+I�8��#���O��n�Ơ���LOu���@���og�OF4��)r�U����7H�:�28-7x"wA(�;�c]��	���m;�M�'�KDzV D'�g1NY�g���<|�jw�g�PV����u踋�o�OY1�����8$�L�y�PO^Z���X�&�g�0Ov!�z�Ώ�o#�h�×YajpXS�N�.�7;-b7<~���w4��H��A�`���W]�.r������xO���sP������LX@6,&o��s��s���(�������O��<l��B�&�W'�ޫ��p`���]�n��:�,ikS� /7[&�������E��g�#�f!�z���w�ƃ7cc��"��a�I��J���9�9y=����W!a6�.�q/��u�${u�֟�]xa�����=�;�z/����?��Gur7���'q�'�̲̻}���ϡ�j�a�'f��X�=	4WaC�����_K��p���`B�,/����jXv��J����O�^��ܚ8��r8}�66�O闦ը��j��V����<�q�w�YE��f�:ܝG��ܚ2��T�ey<��_e?i|G��iDȚ!��o����q
N��d҉=�:��	B5k+VX��f;�x�ᚂ�H����2=h���9����?�r��A$G�����š~����䎞���|ǁ��xR��JĪ�#\v�	�"�-S4.���%��n�_��J�5"��"c��Bb�[V�x���kW;ulS\^�@���)�Sp0F�z���C��t����D\U1�Äa��╦�Q�i]�
�c���~՚�w�b�RV:<P��L�jV�SZ�C����s͚�'@�l�F52�^�5A��"d_��q��J8�Dhh���-sST��d٪��4ƥ�>¥�(T�,���~i�5%�t��3�/�w-��r*kK�����ɓ���)�
�16H��N�e����2�h�RrKɜo8�}�F��?<ݼ@�d��9���)29~�O������ �`�$�Π��o8Ñ�1[�9+f{��}X�j�(u�W.�=ͽ:����"�6�.��� �K/��C�cK��ǆ�T��[���q'N^�RUN��Կ�JNmj�1�ޕg&���}�ѯ�$����dٜ�K/�CQ�P���OpJG��ľ�T���ܛ�)DCC�4�K��>�V������<�
���¹i�|6#M=܇�!S���$�f#���h��Ɔ^fM���b����*`-��g�'?gܷN�}�\�`_Um8~��ϡ�2s���wԎ�I��4�t���5� 7���!����i >rҪT/��_d�Q��}�B�b;���&V��	k+�mt���ҴR�ؐ�Sk?�]�`�9�A�f�J4��t{}c�ؼ�6�?�n9r�<���^���FN���6%.�b	����ojd�W�|r*yr�h@b��W2��'��;&��04��%������������x��U�x�^۫Q�[��D�~���	_�Q����"�oq�s!Ò���[6p4��������m�i��¤��F�h_gk5$��?�V��\5,��d����$��;��JAt�0Xc�f�@�pf.e��ԣ�[��o-#}�)@K+�(�!�M�o������M��h�G�of]��K�}"�*�����@,{6L 	�Ps��h���k��4v�G_�QJ�,#V1�;UZ��Y	 4�Q7$Tc*�C��?��J�|"_�[@����l7��\s�����V<���3��@" 9j�h��i�7����Ʈ�7�%��[uU\��GPl��A�x�p\^���{n|��L|^L��G�/p=E�ag0���t_�~�N�=�R���Շ��ol���c�nz%6l��Bt���]�H�w�!�_�1�r6~70l�^�6��r��Z��}�W�?<�L���;���4� }7i��]E�*�DO!��ax�k�n'�7�G�Oay���m����@�ϛ��$${��p�9�u��"�Sm	��UV�x&���n�C�eɼڢ㌄0��#��NB0���R'������ #�-ܧ8�Z�6��x����Y��%���ֆ�26?���r��}���l�N�Gy��eˋ�� ��p+����)�C����c���#�<o��������4y��9�-H��Wi�gmœ�^/1(5�	�n�S��Q)r�GɊ��o�:�]�� oI�`<����f���i\�v�?���d�m�ѣoi;ej#r�&�$A*��~��>6�F��P�"OGR�͸K^ܼǿ�WGNC�UIs���Qٽ���s�6�&�~�R�Fܦ�lJ���H���KS�1��0��+�&����AӸ2_Dt�D�O��2Iކ�4�ym��-�'a�a9�~a��c����/�U������3�֚SMS��v�,��в,���:����vGU0t�ƴ�U�9y��U���pK�A�,����ϋT���?9�D�.]�f*3,���~��Y�W��sA/&��j�O]��0"����M�Jt�b�5��B��)�۶�׋���Fz/�ܑQ(ZL����/�5�L�^���R8}6�g�����qXU˅K�\>|ID��¢mt����9_���
5Z��$�-�#�˵��א�W�UKaRy��u�$���yƾ�F?�v�Xm�~%	�-�
�����cg���T�o0î�8�3#�ː��"K��s���**�c"I���`����ec����I,�"��˝���Y"%���]`��F�B�693� FQ	�mzK6\�j�8��T���8�ѓD�D)��}]��!̡�f�MFC�mi7�DB/�m$��&�����
=4�i]��_8MX��g�F��')M?20��u@P��_IR���zm����9J���/z�.!�^��t r��yv\X�	g7�R��J7�������:Pb[b-X��>kE�2[�o��Z�[>��Bu����/r5���o�1����x0$�p/�ER�3�����ƙ���N�`�G:6o��ۓ]�gR0��Я�,�_��I�� �1�w�w���hQ	T֩���un]�{��h��@4	w�Oa�}�IJعI�0��Ƴ���Is��H4��xont9����	d���3��s�:2�G=���,v\o�P�9|:D�Ȅ4�h�#o�p�Q��ĕ@I�r��	H��~ϠL�xj�Ku��,�;5$�f{��*��@/s=7�g���S�Q�'�E�I�7�e|86a`|��1��}�ȗ_~_]Q�6#+K�nGC���Pfa�p���uп���q{a��l�������;��<� ]���#D.o:b3�A����L��N��K#������t�C���ٯ��2⵳
�܏�v���|�&x��Oi�)����������@Y.6�nf9�ɜ��
@ά�͇ۘyxm'J"�$�*�B4�V4/X���4�âJ_ ��:J��<{���ե�/��#�@Ћ`���s��Z���Y�n?��ĥ�vk�
F�i���j��V�_{����t���jJ�^�9�G�����2�O���iEw��\0��6�{���M��8���_��t���"�k��@)�#2ۭ7
�}z1n�T�Ng�^[�R�!'#�v�(��MF�24f۹�PvL �S����Bgk���s}�o|G��n/dt5�U��i�'��w�*L��o�!�o���/U�	m����8�ƃ�dFI\h�" _��I��k��w��3�2pЯy�k��$��e�F�Q,C7Kp��`ɞ�Ϻ�르+^��:ȁ]��?*-5XKKy��G�s�?(�)��P�c>H31c�Sdָej�\&�GO-R��r��0���R�B����P/tڡښ
ԯ�΍u5�]X(����(�[��b�w��Cew���z���#��D�~G���c�'�}������(s\�txqĶ؅�v�昽�k�/�L���6l�BIto�2�Uy�<�"��h��1�����m���"����PR���#S����|ڦ�$fH�(W����q���a��=yąނ	4ƀU�H�f��]e����&���0N��&�ߐ�*�C2���^a�(���v�x�U&(����e�LH"Y���[g��҄���OpʞV`3��;�� N�Ӧj���u��t�h�e�@[Ho3]{�`%&ś��Svi��r��
��0*ȁĵ��Ctyl�� ?�G�rK'�Q�c��X���2R�~�:�ZzX�1,O�Qs6F�11�uؖQ��bv��3!7��۟��v��� d��:G��o���ӭ�	9��-kc_��5z��磬f-ŵ�*˔�7��=�&i�ǁP5�ڳ����`��3����L�4���)CD%O�E�,:.ƫ�a�n��i�σ��ҿ7�	s�*�p���H܀�ru�Hi_�T�,�h���ۊy�����LP=+@�&���&ط���=��v�(�w˷Ze����yK�4���q�~��u���Tܕ�~c���w(����iC����\{�����0�������������)7	{��0�3�dͳ%b���Yz̤�����'����>����DS}�l���M, j���:S*9�s�K
�P�Ύ��9zM�ݸ��#H�<pQ�>=��3���'��p�ISɫ���-BGj�,yQm�mj��s�
_�a;�PɴIZsȄ�["nI�2ԊHrU��1e�7����d�:����_ܦ�$�S���F[?%��V�0q��Zc]�.a`�M7{S��J�t-�� b��)��Yl��sF���8�a����B>����P;��^?��OY&3�P�"-O���7��@����ZCe��_i��v#=�Ӈ������|*ԕl܌`��������*p4;�B�a�ʎ+�|;}p}!z�4�J�N��T�V�i����Ξ�7wjKw����%h8i>���K��6�g�"��')�Ll�@!���)f��:,s�68�gx���!p�y+����e����]��"U:��E+��K(�u���R׌�AXA����e-_�p�7m����n@��<.]c$�X����PP����n� �afI}��y��ll�����u���_Ɇ������
L��MP�/����efF�y?������ �"�He�"���}��T�]K=0n��z6��HXG���*A'�L��nn�qX|�tMa@��ʅ���_=���b�M~~�4���3�x��<�����}�q�pS��w�~@N�ygjA���+ooOŗ�+���+E�>�VS`<ܦ�&��7ia�k�nd+�$l2w����q�Q���eø����_Ơb�}�V�u:�O�	�� ��y��Zj}ny���HB��T�� _�;�G�9c�oZ���/o���LK�{!7�fDk0�t��Mҿ"/���գz6)n�!�za��E�Q�K�͟�h�2��c�	�&RA2��g�J��dR)��O��7��c /_%��LZDY���zX�	�����t�O#,Љ�oA�|b:�Ỷ����='�[J�
 R%AG34J�@\�Z*P��+������}�{����#ǦЃ,$��nw��!r"ͅ�����Ռ�LsM�?��v�v�e ��V��������ڈ��%�b�ʫ�u�1>���ܼ�Z =t�Kj�/���Tc���JN;D�I��*J�оV��
v#.���Д� w8�`y�O�U�ɰ���v&C>����x���U�{PY���������s-���>ʶ��Z^٠���!Amƀ��?�����<�ˣ��S����܋|�������̒�vCF�� i�y_dt˞�e�g��p�m�����x^�O�Av�f�$��.��	���rqM�!��Z�u��v�K��,�)����'[�|ڈ���4�*�B�UP%��=|bh	10*��#q�Z�W���A
ؠE�m`8��e��*�DS��1f��U(ٺ)\�K�1�Y��:�����a�և+|Vb	��F�~}/RFu9�1���?�J�l�Z���壘��H8��G�.
�Qo�~=ŗ�0�7�!��c�i�������m��P`[�L$�9���ԣ�EGlp�*�A���|��r�NK�]-�a4Dˀ���\���vUtXc��R	�d`�^��<���&���K�9�����ɯ��C���ǲ:0]���b��{�7h^oU��"gg�R�AU%�T/�N?�=y	*y��GrD"P|�g�9�c�HF�]�����k�x��jeD��N"���t[���z¦A�����/�A��m&co6q[��m�O����r�R�,����v��ԇQf�#�!yi�# �
�ʳ%p�Y=��ԝ\I��A�摽�<0r��US��[r����5�ez�+����6�,54�Y�ح���L��ڈ�`a�S����e�s���!%���t)4�c�9��;����\�b��(�q���lL R�M�.<	-F����i�ۚo����Ya9и�r\L��͘n�n_���Z��ft�~�6�.us���_i�q���A��O� W.�@��x7�o������t�	�l%�,��M;�!)�#)����KhF�	Sb`�p��2���3֯�"�~�ћTڨS��PJW>[�Ay�h�E$�S�kE��'Qog<�*�JS��������iO��kk��S���!jY絍�8=uO]#[{Z�b���)ºpzN75ٖ�����#ִ�����KoTHY�k��E"����w������l�a��c�P�k�|{0��j� t	��q�7��w�,7�0�5�!����beS�u���cvY�d��y���I��u��A��G�ak{y
��'�>�����P��4BK#�q��:C�P~��t��E�̥+�Xr�}��uȾ<���5\���'JT��M�%�Z���g���#V���f����D�wh��L���p�B���
�񆧚�2�(b.���>kb2"(�ԧ��=����J��Ւ���rF����/��8ȫ�Z����L@�]/�Q�v��w�8�����8�?O`� &2��RO��N�1�zZWR��%e�PX�{�p�C�	��/66�-LO�ԇ�d�&�1д@�m�X��е����4�$�̤��*�-�	JBeɲH��s��u��}��+�Ʌ%�-k�6���!�COR}&��ǐ��f��9 wB����"�	��O�Z�떿�p�w%5���4��B��X[�B���93&*�7��a_��410�I���צ�çq�(d��:�fCU�3i�)W�(�d�ӏ(��sZ5��A����!�Rz�w��?#��G��5z���%,��HP��D)���bC`��^n�?4L�� v��1���Ļ�AƔ�F,�XBV�D#�Y����]����܍��m�L�^!�w>�ԇUY�n��P�(]�T�Q�H��5$��+f��D�
S�����>+��������$/�Š��N����9��{ш8 � ]p�F�<�I-���^9�y�kWL�?;vJ��\fF�;Xf���9���B�|�9��o�=!�[{�#4���0P��b��EH��O�������k����ܮ3B�Qgo��Ȇ�WN��?�qS^�Ӆ���R	+Z��]Ϸ`'Њ�T҉&�ǈ5�9/���i�k��Z�v��a�9Y�TFQ"D:ѥ^���� :��<��{�Kh�b���L��$����Uw<��T����e�}�����Z�Ev�dCi����u�l�7ç&���/Uc��F�fM�go�Q��nA���e�K�!c���=b�	�w�%�{���T�z\�ban'��7�؂�C��{{�	 �f�Az�?��<n��S�uD��pF.D-TQ.F�R�ϰt]��꼑b�	�D�
��}k���ׄ饂���*fo�s�gG��b1ӱ���dW��	V�7D+��`fXUQ��ZO!��S:���Dde4}�p����(���:y�08����S����a��l�Ǿ'��PV�8��'���3Jįh��Z�}`s�:�}�L�]�
U�Yk;��%%����3�jF�х�I�#�qd�58�&���Ԗ��& ��獞M�t�li茝�cx�0����v��f��q�3j��4$�s;\ـw���������S4H\]�i�Oos��7�㠫��]�~s�-�Vz�:n&�����#�TwF�@�;���J���d,�cb&ݘ���E���P�p{�$�Ȧ@�~����D�8kԔ $`e�S��I�"f#�CMx����m-W��'tiQ$�}C��w"������g�d�A���C�UF�;@�t++=;E`��cV��sc�Fs�;=Q�5vRH�,�w��e���?�{�=�;=\>hHGs(�
@�L��^�l.]Cy�S\ Qi:�];�9 �c�-7��%��i����I�;�w�����_D�8GѴ*��=>��{3G=h�I��5yB
ޘ���϶X�	�w{Gk�͢�(V��E8�z6c%�ו��B�=̹�e3@�>���z��7%"I������A�w0�ڮ��eT��%�L�׺��޵Q
����7zQ�@P���ך���"-]���e�u�OҴA^���]��U3mJf~s�N��s�:�g�}9�(��НR��$4ۓ��@���wy�3mO�N<𨤹p��<_LWa�����#�q_� �A�iθ��z�:c1{Њ*�o�y��49�'��b�?�O�P��iZ����l�;��B�^���Ҫ�"�w��T�\LB��q�0�A\��]�Ҍ�����D{��$��Fe�RK�$�!6�F�+�Q�#wiݗ�ȷ�6r�SO>�	�ǐ��(,j��q��Ss ��Hq�=O���A1��m3�XW}�H������)rĸ5�I}�՟�,�Ĥ�	[8KD5�Q�Yg�����B>��;�ׇ@�̲;q�W�m�3�)��7 K���F/iz�CvdT4�&q�.
)�H2,(Śv�@f���p3`��������l˩nFe`2�3�T΋?!)�\Ѻ4"$�2��Ia@��/R,�QQU�t��Pޑ�O>� ��Lo�,����q �����ä,Rt�+�T�@��;�4�m�	�f�[m�\��d:uY�
��t�f�^�8Rz�a��P$d���O���B���-f������H1�x)~�^���n�s�w�<\����ɪ�|��9�j�z0�Qs�DK���f��Bf(%�"+�҇��v5���]TL]�P)�1(�=�P9��y'v�l�(�,ڊt)��˕�;�onCz�o��&Ӊ5
��/e���1էc����b�On�)�,�1���#ȉ� {\�5��̀,5G���g�m(<F�	����& Xy  	$	�w_�.fe 2_3���T�5����mp��(�W0���Еf?4V���z�r��BMN�Jq�1�r�j,�"�w.��L_�e�g�y�ey���Q`���=���G�$�JI<-T�׫�3UXv�4��	����?��K����+�9@�|Iߙ�u�����V�h����j�Ό�j��?e6�]��B��PH�6P�<c潿LC��Pj��8C[�,�Т3q#�x65��1��'�:�F��z��B���ө�����c�b�Hء\X����ʦ��dG����Iz�����!�hUh:	�6s>�z�EB4䕮Y��[&�?1Ġ1�y�`x@�Mz�(Ya�L�7րsN�h���ͩ���2��J��bk.�������p"���?Q;��DJ9�i1{$�Y�"`�>~ch仛߬���.HC��ଗvy���|�9#���8���$��M�L��>fO��{���*t���|�'��B:=6">�_�>��)�wj{ϵ|T���Rn��^���a�&++>[q��� =8�m�2J�/�@�H�W�3ӡ*���������2C.2�ר[����7����`��ʒ
����G�Ш"fj�P�a�=h�Ln���@.�|�vn� <����}ț"������g�'Ԕ�b�I��T`H��W<���M�r{�a�����>;�����+nle�޶]���c��ls΅��E-�1E����v�5M���9��L�,��;��NY���L����B��@�P�Ѳ�S�.���ĞSC�t��L�:.�`�Z@�5yL&kԀ鈥os[��V7���芑x �c��W�BMI�!R˄Ւ���`��oوi�ۣ�PѡJ�O���!������0�]d`�K�|m�7u)�4���j�T����u	;�1��)�w��,!��g��_�"�[�G��c E��i��ez9H�M�/��,����.�8
���G�m��錷c7�/-哳��uz.jx�(��YG'�.�U�)\�@��5ЂZ�\���Ni�Ԋ2W%c�%Τ�_ʞ�B�m��k1����\%SY�{tG	���Ɠ&�y�x�TM;aO}�\);��LwIQ?TcRBkU�(��0W`�c?����R�2�W3�U�o[�(� <�X�A ��gy;�������͛t�铛?�
��~-��r��[�ɬ����}o�	w��������*�-�q�~'y���s�	G�D��t�}��a5E I��vK�P�}f� ��X ��O�s�����[��S�u��x��1nl�a�
�X��1�n~��w�	b8���Ǝ>��B��E\���e��xP�KR�iS++��N8����k<%\�DC;�*�9Q�Ӎ�2>�+TDO�K��#i���L�߹j�^w���:?�=���N?�a�)�;�����gk�W9��g7��%6�ś)u�k��&���=Z�аM����rI!l�(�c�:b�����Q�'�=cW�Y 	M�t�ʹb%p�%SF��F��O����YD\�y�*����5_�7t����ߵ�����9��1{C��j�x�����OLhw���x�(�9�tˇ�-0����sc)�d��Z{4ۡ��贠J����dL7�y_�6Rت�'���)DS���R�ت��
�1�iq�u�)c�D�/:\A�?wH���}��&�������'�	�U��w�X�g�i�_�=[��q�~�5[���ۨW�X��5F�3O�����*��M�T����!<]y�7{�)�L�bZ�KID�Y,�#��6ͨ�һ�������;�T_���#�4�}��3��J���6	R9����c�&��-�D�3I�$�p�թ�!=�@o�,uO��`�sd-@"�����~�]�0�x����`���"M��ɳ;�G��$�E\��.v�ً������ �\*6�,@�V���`�LF@�c�������Dt��[�-=u �h܏�(P�=���+Hތ&�:wya�ɳ��F�m�F��b&�����
�Hm�d`��Ƨ��$x1� Up�ذO�#l�Fwܠ���j��S�=v��*��
Ml��>�mg�^�W�0��S�k?GK+o����^�Hk=T� 뇄��%uX:�l�2�^�؄G�a\��E��A����O�)T䪍2D��	�N%
C<*[2-O#�=��m7
��EZ�Le\1�
�ilc�<���^ce��;ޓ��:ӳ!YH{�����wiD��UnNё��"�iǤ��	n�����%: �ـz�s�f�=�?��;�F�F8����X��9�J�qk����ߣQ��NA]�S�U@@u�9�}m�Y �"�1O��= ��y��D����%�)�L(�K���rI°��쟄J�'�?rϵB����5�>.p�or"���Tn�"Xw�@���Ф�=W�=�"#}#�H�:�5,������3��!�?G��X�}�.�rqi�eA��+�&���O��bV}\�V�f�^�@��_zi��r�EB�P��e2 �ع���d9/�,���u��' ����R�(����/��dU"��Qp�3Ž@�/qg�Q(�ndQ�+*gy���0]��
��0:�l@f�9⾯̙��˓�Y��^@{#��ܺ�k�b����C4��	t�|�m�e}oC���j(^��Av���S� =[7ks������?����u��Bퟁ��
�GR;��l�3Q`�:0�9����)d���xRt�xE�2�����)�!�	�q���?8�8��l�֮���K+V :��?L�A�f+ҝSR���s9<k�Z�_�H���{�fk����8�;<]4i�w�▓�_�ĞN@�R�,Fj���q7�����{�K'��<��� 8���\Z�w*��[�z6o��O��
�qQ�]�6"SI@2t��:�}.�����i��V���xs�|�=�`��7S�="L�M�V���H�u{I�Òz����=�Y�Q���_�Hs���}�}7���߈�#�x�y�|��>
�j�Х��G�7�x�+sa�|�5���Fh8� �ը����8�Q����y�P�P�P{�v؂�)n+�j�B��'�<��k0d+�qτ�b��i	��3I�BJ3��p;�M�j��b����f���M�����-��{T{D8��s��P0��l:J 2
����ĞA�B�����e1W�ůϖ�M�4�Eu�Hp�,S�/��d�%&��,�^�踂O��u�$�'�#Z{c��=~癩Kc'�� �`��73F6{�q�z�L策�%��tO�$㇎&���#?-1�z��N��/��2YZE�0����\�ޭ�O�o����	���u�}6�y��
v�a(2L{(��g�/U]��AXs�_5c*��v�y�����u�\XZPl����Fj,+Ix}�>K�����bP��"�*�д����P]��C@F�'-Bmt����[  �/�g2�� |�ea��1��y�&�ܪ�*f�#:�ׯK4����2Ɵ)�ޢ�@Y-��ڕt�+��N�zԇhK� �~�L��<C���V �N�)�N�F�7Г`��=������7���Z���G#�KK���5����R�� O��M�E#���v�O�r�u`1>�����&���n�mϐ��T�Q��|��l5/+$
|5H�))�n��h���R�'R�w�{�>�V������:F7�4�z���.��ވG'��M��M	},b�T�_i�f����n�t���p��ղ�r��!)B��vm|�<��ܧ��a9z��<����!Q��{�rz�!�E��� :%�0��fʢ��P��v9 3�"N+�ݚ,�q�Oh��x ��Dci��~k>�j�Q���*4=ݛ���*I�ϪK^��#����6�,����?�X��-�@4�z��+�2���0ظ���]�c��]'�t��/3���P�JE�	�l��[\�:�y�xN҅��W�����op�C�]��O���$�)�f3h��.V`h�l�n�47����}��h��8�DG�3�pH���?�6�N� �y�ϧ
��������O@Cy�JO~�u���V��(��ZD
�*���eØh����Vآ
�+���(��]�#-�։w��ԅ6*��:�`ö��ΐ7�n5���/��gM�)�R��2�I1�O�����p�O,��0��+.�7�)EW�� 0_��Sj3yޚ^����   6�؀���W�'�6-R�'�3p��	�q��Q�I �����J3e�����oɈ>UIǏA��R�"}�g�t��HJ�E@�m;!+ %�����_H��(]v@��7�<6��y��]�)�h��ӈ��ȕ=>����~���_W/W2-fk},�_4�h��@��I �g3�}gA�NA�1���C<��i޹��h�u)�/jK���~(	o$� �M ��Nq�$
��1�3SU���i����4�	:�8�������k�'��y^��@"B�Uj���Y��Ƿ5�)K$߄83}�T���^n�M����#O,By���a);������ÀT�:7�+"���|�o��	�@qO%f"�v��SY�:U�3�����G�T)6Ou�C�5!���Tژ\$���ޣ���$�<����SBiE��V��,���ar�/����H�^C�|��҂�]����!M���D��T��Du����o����6;NU����Ԇ |@�P�<��nc�7�p��j��n���I�sʔ`�}]Z�Sn��]:|H�׮n'��j��S7L�MK����<��@����WlR<x����c7��?�?��w�*L{|�������s�`c�����B�����ń���UE��W�M>(���< ��Zk���D����z�\�gȤV���2t7��
�Qf���9��N�Nz=��)���C��Z��VJ�����5��K1д x� UƵ�7=�%;%�������d��� S�̈g��-��p�Ѧ�|���k=+
&e\j���b��o���U=+�M����D���hRCx�ԡ;,�����̂�a`?�jU`6���L�{���p�ݡ�&8��#�xhæ2��	��`��k�Z#<�ۅO��ؠ���]~�8���C)����7xk�+�>%�(c�(���� ��k�xfW��'��$n&�J�g/����]w���ޢb]\���X��㥜}���R�Rٶ��) j]��ӵH9����,�3��Y@��SX�7S���+þ�PIV������͡� !�}�����`��1T�3>�Q3V=k@Z�(q�E�<*�Ħ;�E�)�#n�k�v%�*9`U�fb,,g�B�E�H�>� �*i�~�B?-�l9�$��&��x�����:5�a3	����^L][FDh�#�-3��?��5���=�З����;��i+�J�0.���17�yϷuK�����5_����CFH=����/���cn�2���/ͅ�D�@�G."FY�W�RT���!��=oB���[1���9e.bA�-?�5������������V~%�-}����R5���D#MM"d��f������K�x�UN+�(�}Ld�@:9%�� q]�r��B8JÃ�7�С�ي�ݒ�&;���.�Ѹ3c�Ƨ��La+���i���7�(���v�>��B5��Ae��c�C84:+;e�곭kd���̢T�#@ud��4���F�I4v��J��(PےFFϦ����D`�<z�BX׈����~�0sp{�H^n�6��7�c�P�g�:h�Պ���3����n��2�}Ȃ��
S�y�[[	21��W�X,�Z�����������Ii���f׳���ս�7��q	������F���W#t��s��i�Zf � ��T�3n� �e�t�=��jo�q�sv�x�u���
��/�K���(]����6e:ӥ><�V�)�O�݅{��a�����L绷%����;~�gQ&��T!��G�e�ǁ�ם�b"*8T���5�4}��x����'�<KϦF�ZT��[=���X|bT�߅�#��Z��t) ��+�5���\�~�X309����;��+.���91�fS�[�:7�ZC3`�n�t�y����=N���p�پ]>pd�@|���.ܶ�t3 ������� ����Z�̸>���:~�q�iՂ�_,�s),#��%���������(���3~�
>,�����828�(���#�Wåe���~�l����D��/`*9�p�2o>��X��gV�:��tQ���l�"R����,(=�F�����g�d�W�z7��U���HH�ܗ�������l�WT�ۯ2��s�碑 �K�wT�]�T����VȈ�jJ��9dר�c���O:O�
"&TM���X����e��?����VA��
��9Ǡۂ�h�(���RX\����o�Ϟ{
�a�C ܨ=������TF�����&�����^aV���^��P��gt\����G���~��͹��47,9�h���&�V]�����^F�:#ss&:�p��"/��|�Q��-���ֲ�c��O��?5V��T���GG��a7c�<�ď�㾗����&���r�<�!�g��"�W
ة,;wR�|���ޣ�υɉ宺���4�'$��;�_Î�0iK�L�Լ�f͢�l�M?H��xC �$Hn7($ò�~��AOvK��T[�Eq�T��Ļ�A��Ä�������N0؊�s��d/�-6?U���>A%��@���7h~Jxt� ��ۨ�,����_/T��`K={$v�g��*��|�Ձ�bWb������&'^�R��泇o��\.���o��<�qm=��w�e4U��1C��6��ds�a�qĝ���}
�B��ҀF�ppx�͎"Բ�I��/�}̣��f�
n�����v!�U\/j��������R��,t����cːR�r͖��U�"�/1OɈR���V�Ԗ7�C��2�2��Ue%�p<%��k鸙��ߨ���9"h�*I����4�&xg��rJ^o�2q=R����+Ը�{j;#e�o7'���ȑ�6�'��o��S�v��0�]J��JZI�pΤ?l�i׭-�1,�Fg��UR�}/�<#���EЌW��ǿ�vEΜ'�D�,+ѩ�Cݔ���t�o�@�RR��J�Ǜ�����Y#,d+����̷;�v��O{��>D�^5��f6<������)��c�	!�a4��Q���g�i�Ι=����ATB�4},>?W=c��;��3զ��VV���.39UY��M�%*Χ��Tp���V�y���xfh2c��).����#F�xf q�Zb�W��/w>	[�)��,����G_��"��� �[u�*;��#�I����_��Qx�}�c��5��Y�ʜ�����F�j�߾kՅ�$�f����<�`���вa�j�x[@���*�oZ��.3z��~ڀ���������è4U�}�S�ٶ4�^!n��?K0�A9kn)q&�1���E{�pG&��h��8���)H�6�Q�.��Q?2R~��v�/�&͏��c񮔓5��T3d7����:���`�̋g[a�t�q?&'��8�B�P��;�B�Bԝu28����\�1���qcb��md/2&Pv��7�fB��E�<�c�#�a])��b
��5��L�h\T����J��ݜ��JKjBG�����9H�'���C[�L�IM�X��,��n�X��?�3�������3�A���P�W�]8[cu�8��[��ۚ�iq;@k)�5��������z�n?b�jA͠oy�d��7�K�78���kh��v�(\���	9 �F���"'���[w��+>䔗G2�[x0��q�XЄūJ>r.� @�^�&h/:�l���/�t�e�	����y�c�|��=G�%�X/�<��M� .4K�<
	E"���N��b��U���@)�b����Y��K1��R 	 $i���A ,���lYV��(�J��U���D��s$���)o���ËK����Z{����"���uL �������i3N5`ɴiD��h��@��`����8���{U*�1Y���0a�=���a0q�~qJGkO���V���v�?Y�e&��u�rW�s��e�-C�no}��7bvF�k��g�T��EG54���Gv �H��@�臍�����_�;�~g-PJ�
Ea��[�[Rٺr�:�mI}T�	Nx�?� �X5쎈�*�Ψh�{[�mwTRH��z�捬bxGKc_�:}NI+�Ǆ�g�D�����]
znZ�@�Ű��<ً���t�АY�-,�?z�J��C,�{���=�s/T�
V*� �a�����p�ß�����O����Q=�������� !�7���sf�n��Ë4�?�9u~�W#�~�4����82��`�������N{�����Op��g]6B����3�л�0�|�Е�0��;Ȏ�4�a`�B�b����E\��/�C�]�z��o��H���Z�3|"7�L��"�,ݠ��}�B��r���~��H���6f��Α��.��������.���#����x��p����:y�4Cuh�Ln�@�K������ͼt|['�a���6��
j��hZ$�2���dD�q�]
�jϞ!+�\ш
�F,�3t~�|�~��<�-[Y8t#I�R1i��oXK#E�xxp)��B�x�վ�'�����<)����BE�� ���"���{�5Z>����Vj�s�M��w!x��:P'U\�Z���6H��k<�v��'����v�ϸ+@B����)��j.��)Ub��ԟQ�����d
{E���9�V�
��p��Op<x��k��	L�^��o`aw�h'�k�oz�����Djq����-c��e6�JމǴYKg�Դ�p�d�mG֤֍n���ʂ��8_��zW�	ł;c��x!
s�~�h��1���
؍d@@�%}Z�E�)�v�, ��-�+V�y}#h��,�͢|�ׯ���T�a��>��LWҢ��0#��T^��FI9��7]����POL=�ڿ�r����y�;�}��ֺ
�V鑋t�@Pa�ŷxyi�Z�?�y����Q),�t���bP��T�7ZIӃq� �\.Ib㋘�3�s��*�5,����A�1t>$߂�*�g��A�L���n��ד��l֙�I!!��A���a��[lh>ǤU�F20�E-GN�dH��ѧ�ĥ#�$JqZRT�3DFO�kp��(����d<d 9���"�N3m��Z%�_�|6�h��t|�P�,`=۴��M��|���uvč�7h5I�N���$�ۅ{������N����ʋ�vBū�94sky�W�=�`�%�=�K]tm�Z`x���ڇ�6�r#5��u��xPД)������" ޿�<N�՝I3��~ ;42% &Q�=G\�;i��N��hϔ`�z�:<M��g/��1��1��	��9󾪨y��@�����tۇ�c�V��ns�� $0/�\���)�ŏ�[�y��$��e�h���%�#��� #̉�؅3V��	[���� :&L%\�7����G�h,�&��6�z�=�6��u7�[���y�n�?i���"��P@��c-�'��ͻ���9�EI5u�����?tKHܣ�Z�?�HՃC4V�F��a�*`��: ��Z̍��%Wn,_���s/Oql����wS,N�i������d>;�`X�?$�+���0G}&]r�Y�~ޮ S����8$b!B5��ܩ9�\�)��"�ӎaeiw�C�։�	�Z���o��%���}��2�i�G�q4C7r?���5�MS�E��̫;~�}�s�2��lLn�@���7� �H���46l;��[��7��u.h�er �(�ipq1��*��˭=�C��[$0Tb5vO��5?��S�܍�G�������}y�R#��T,<jq����fW���Xٓ�Υ�<��i���)2��"e+:�FIu��R<Z٢Ǌhc�&�q�%�O�3raGQ4ѩL�S9��<5��y�,#�D�u��.�[D3/U�i�&u��!7o�I�ԫM8=��_4R)�A������>�hCwtL�p�p 6��n_h7`,�����j	&��'���? ����j]�;���f���%�GN?�遯�<ӂ>0�1'�zp�<���F<�#�k�<N�S�# $���'ū��x�i
b9 ��L�R8c=��{�a��4���
9/��Ƭd+�3��a���GH�݀g�zc��ap���P1�r%��ň�49��貺��+��l��uHs�W�?�VTɣnK�Н{�K���%� G��>Q� �7t*=��i�t��#�7�(	!'���S���i#:j��#�,�q.e4��2u�4���5c��	_�vSoC]|v��.Z�l ���XQK1=%�����ه�{복���Ҵ1=���ȔJ[�<RM�0bt&/l˛����ԛP�@���@�U�D�u��\��t��4�ɞ��$��9�C�зV�=B�gȃa�|� ��:kKR�y�,�K�˱�z�Sfm�5��h�;Qlԁ�%�/���Ŭ #��o�Md5ej�M.;��mTص�B@&��_RN��D$�5X�`���	�Ǚ�?�$�`�������j�#e�D���>�\`k+>�/��`��r�d�� F��!5~������]Z{����+(>��P,~�B225b�h����vW� ���៷+I��N��,�;�%��1����C8��)�lC6�.�����Dn>>�
oX�l���C, �y>�)��[w��o�=!��Rc�U�Wk�R�*�@A�����y}���N�j8}� 5�k3�x?:�$8��K���˂�'�0Fl��;k���UJ96	̎��/��Q)֨�.�?���q�V�G%�/k�H�x��䒘��Z�-��򤴁`l]��#
��T'��ew�h�UK92�*�"w�Ig�*_��(�ޝ8� <�JchFl8 I'��熯�i�4Q_Z i��ڴ_[��������J$�Ztq�(O�	��\�tˁf�aJ�Ջ�4
)h @����C��x���T5��TVf� �c��Y��S��f�X�<%���M�*����N��-iʤPg�ڕM����{��%)����i������H��{ڮ�z�$�� �g�v�ˮR�(�O���]�}��~�ye�gɡ������70���[�Z�nA��eJ���r8�����[��{�O�*�W+x'�mk�!sd$�V���"�*-s�q	D�O9��\NU�����M�k�	 t)�[(�.k� G�a�}��䯊$.�#e<b!����A�j ��	^�̺l�?��b���Q
��� ��Ѧ��5�� J�nO9
C��īf8�m�����{xI���|���u���h�;�w;�Md4� eVM��C�Gʦ�!�?!c�c��OkGĉ{�W�q�d�����T1I�K[-i���=Յ+�����p�G�I�A��B�������c~�D�@:[d��<Go��H�Cp�ȕ���R�&e���I3C��Fy��������������B�JD'��pX{iQ�}/�P��D3g�h:�ׯ)⮹r;���T^
����{Q}�D9o�8\
��2筩�p`f�Ṕ:�M�/ھ��Q��)��?&z-�@���j`q�A�i�a�}2� �����~�j2re�qi�#���0@Z��ݙ�>��� ����eT� K�o+1��|>��th���BN����߉p!�p;q����]�q<���y�.�(_3Mq�i�-�Dfk	s<F.~"���2!kvVӵ�,S����sL��s�"fz[ ��L)Ԩh������8�EX�PĀ�p��g��s�d�Y�d%0ȇ{�(���۵�t�����<�`��ѿ��!gyo�(�.c���&�[R��[������!���G���lS]����OFj��7���>0�{)�+~{Ў�# sݪ��M��٧���L�M��||YɡC�Z3X�4y;�������k�
j
��o�*�� ��_��m������'qA��h�7d�3�\��N=��@k�B����8һ�
�t��!���e�py�.qΙқ��*#�z�k�=ݵA����[!5�
2�#P�N��o�A yk8�5�mV���LiW����ie	+B��L��"��@�$�g�K�k�[pF���5��]���bϵ$�d�5$$�p��b�<�L?��3��G������cx�lA�w�>47��R���V��ZDԀ+�K���::y�������� ���W�g�X^�|c�Hq�kI�y���0ƽ�X��-&��J^���bWE���K�~�r���<��܇ex(��g�)��"#D������#��$�c��/�*^���J�N��\��oV�ú�q��..���}$�/����[m, k�RXKfG��@���S�O=(y���kU�_�)HH�ҲT�g :]�D��.����H�= �݈bpZ��lR��C��^�I��p[}8��zz�5M�%=I8�z��e����q4��:�_^�x֛�*Τ�r�	%	;��D�D�v��0F
���$�Z3��|g��VK�ņE�3��+��[ڝr��ȶ�s=p�\sLu5�ߔG�$�J:�'j���;� �j)Π�Ӫ�0���N�
h"�᫟�#�����g_�:���2
��H�_�\a���1g�����9)X�߾0�9�Ŧ��@u����f�7z��U�+����}(E����9ds�
�Ύ7�]�@?�ˈ��R F�ˏ��!�]����;�]��؝���s�[����}�BA�:�!o/őgǚͶy��UI�F�l��|�u��&�v���7�>���q�����b�:����&#��F���].=��T�{��{5%>��@l�3yy�T���/e��`r����� t���eR�H��� �5ih�|�+��9"B�T��©Z˿����S���W0��؉B$�-]�ּ��Ę㠟��Q7s�T͖Z2ΌA��|�M����8�)]�L���b%�-D��~ꉐ��V��@���M��V��m E�f�����'������L���K(�6�} {���'v���k��I5�)��|պ���~힫�&j��U�_e��Vg����<��Q�{�#�����A8��Q9;����جy��D���%�d��̿O�z�e� 4��rT���nܧ�����(
m�Y�H�-���8�� ���K[���ɥ�3�tnuyl����70H\^۹Q�	�ġ����Z�ev7���%��C�����N-�d�Q�`ʞ��p!G�t%��%�1Kl�j�Up�4�!�u��I��H8����v�����E�^��T��Q��]�g$��)�`�`Ã��{�#��w�iS=, �Td� L�:F�iϦ�*C��9
{̧"'������eMP�q�ڰ����̀̸| ���m�ٿ5��?�61k�:A�9���j`k�����V��9<=K�p+p��W�΀	�3����G�pVH��0��V�i�(�x���d������̦(��ò������W�+,D i����7'�|u�(�`|��FÍ����v��6��K���RT��++]��;�?=y5g��,y�!R p�X*��9�"�W�Ƣ��+�\�I��(n�-�1t��Ȅ�Ԗw=P ��#��hE�ʩD~ۧ������$Y��K�&$���#ʊ��bٟA���ʈ�j�[ �����ƹu&���!>�ϛxY�
�<�[��8 ���~(N��)�_u@��Ӌ�f?����b����2��e������ mx,�^���e�	#�/�Y�����j�]��ܹB��nG6G|��Y��T*�z�c����@֪�;�l���1����ߛn�r�y�&:�Qs�Y�\��'��wOnrS�8���i��[8��d�=H��k�}Ij��j~9���B�.�J _�Ƿx��w����C����H�ܝ����TK����`������;*�P%�g�l�����I�1I� ��s����� \(��O`q�t����ۜ�k6A�4�*5(�d�Cs�o��I�Aoy�ƛu��[w+��cq:jGU��q���P�A�X�(Lݥ}ր�����A��W��E�u��f�4+�&qv��q�K0An��ݎ��{���L#~���`�WXQ5�eW$�3���( "t+�w��B�W���/g.�F�S�dvj�F�ru��{B��xe���`�D<���j������jM�����>�$�2Y# 1�N��9�I'-��K娡��H8�x6C7�/�'�kVɘ��ɓF�ةۡ��+��'���f�5����R��S��Z��J���ޡ�i�`;q��go敡��_H�Y\��@��$E����Ƒ��y���b��npp6E&.t�_�g�$�#��&�\��޶�-c�+�C4���<P�ujɤ�S������89�6e��!�x�y��(��$���i�[1>�~7��Io��䟄Eٞrr�rW�8������2r�<ҡ=P����NG^���I��8���έv����|��9���B�\s� H���'��YD������٢yI,�ُ��f��BW�u�̬�� ��,��� �p�&9#��H�o��&66���0\�c�������4��s$.ſу���ɷ���C=�Q|A���i��\��q�K|(�3��c�1͒|�kkz�5�?i�u�p��a@��\�"�=p�K5���V^������ Uc;�2��YK1S���G��Wg�r�{�,|�\��0;D���#N�H�y2d^(;�G�7l����&�Ý������Z6:�yrU��`�[�L�$Z̄��ט���x���7{�]�ϔ¾]`��b�h�� _T�#;$��B@$!(�t�Maq�G��b��H }*��X�-藈'��x1�o�pV<�c<�\����A��N=T	Ed��b��~����#�S��^s���/���#���rD������S�h�N�۲�_��6�9P�ow�l�G�Q������������#�������/"6O&�*	�'�^���=Tԝ5؇| ��`��j�&��h�"
��'�ǹhfL�ܻ�3�b���G+���$��[k%�����0�f�I�t���?�d{��Fc�y���2v� �����$q&�������+� �
.���05���U	;�wL��%k��v�ݺ�.�Bc�#zDXu�Ǫ䷳��Ħ��{!P��d��\�)�?�w�@�&+N�A"|���S�Ex"I2.��ˤ@����\NO�'茰݆�"pz�=��6��Hֿl3��ץ�n�|�.�-vz�~��J�_X)���^�Lޫ�y̾�##L:�uź}2�Fnz���Y�"^>+�n��{Pـ����h�e6�p��%�18��,*Iִo���IE!6���o�5_݌���7�c�!�fMO�|.Y��E�n�3{�����>��ؠ��V�h��<���b�ɋ7T�#)3��?�=[�(��D��~�W���h�V	(F��X:0����w���5<�B���>���4լd_��D;�8�t�;0���U�.@ӕ�~3�$�'����TM��ЏZ}�{�7(a}��I��kD�����y�]L���h2����7<��� ��h�V�Z"Y?//`�0)�-����QڟE��`��(�G[����S�ᰈc}C�^(FF�����0d	��&. ��ֿ11�'���`gL'�N��V�1�?"x�$u8{�p++xۨ�����#p3�Z�72���V�����A�@��r�e��崍u9��zح��C�r@zq��d�
��p
I��$d��傒�B��D��&O�/4��o���'+�j�JU5�tH��(��v7d`}w�W�É���>0>�5��x��w�Ϳ�`�&��!�5)�-=x����4Cx%艕�CɰV	�$H�A�#A��P��/>L��04D�v���z�q�y=Y�9Q.|G]V�)D1�([��:�P��3C262y|�e��i�B9!�^�LSl�e��]t�0���|�_��5��b����"���x�V5�n��T&}��4z�:AQ�m��q�l��ȹ��V%�1������#�{D��ף��T[��m:�[k1N�9�k�RɟC��T8/G����d� ��Dƴ4< �IC�1��=�q������?�L�W��I΢ެ��@;�;��v!����NKn���(���\�������<܈ RH6kw�Հe9���6���@}")�י���?�G��ő�{r}�Y����5�l2��;,G�9μߥl�����P�C��Ϟ�{fC󉷭��RXsB����t�@�C{S��A�ok���F�����$��}�M��MoA}芙�c�\vo�T3.���;�YI�x���&��hl77"�;Ke�/�V���D,��',�9a|$٬�
�]}*2�v9�Ԋ�ſ{�Gr���l�F����޿c�d~��2,��]���
h�����v�_��-B�Ͷxz�f�q~�i']T�0J�zǻ��ω����5]�Y��s8���q��'\��c��C�C`��s����#	�=��8k-Z\w�
�n�c�����0���O
{1)�=�D�iO���%M����G�m�K���{� �����1S@�p%�Y��"�Y�ߢ'g�!������/�^�>87�D���~�3�N'��}�̍�� �L��2�����si�� O�9v�ww���k4�ꎊ�Ki,ӨI\����b7�9��>������z|[�#��4L�b;��PӀ#U��H;��7a��AF$��x�ǆ@��
$)�'�3�'���2��ZԷѳQ�|��h�k�7�5qI�L�xPź�
HRvz5}0���4){����~q���'T��{�	�H N��a-(�Y��'�o����V�0��$���_�cr��zũ&�u�bQ�}�ĖH|�-$���,��k��5�&��3��i��W"��z�j�ԣ��t ��5o5�������b��`L�"v��V~��!����`iwm�-|��y�\H1k?z��Q� #�;�5�BT�HY՗��aW4,� �r����[�*�f�L1���i	~��+�qh|uM�ޠ��Z�1��t�"��x�c�(�ן>��1�6mdYx�uq�9�^:ˠ�JC�Yۂg�� �+{
*�R��8�[�N[��	l��2�L�h�-؜�kSxO\�r۴�z��j�V��s��j�|�ٰ0���f/�L�ۜT�%�q��1�G-�a�nd6PB�,m�y������ӻ��}>��m�Wh@)^}_��'��(�;�֕X�\�no
>EFc�9=��!�.�3���LG���ULⱒ���T� $�̖zn�����&�D�U>\\�_n����b:¿���4���`"�������j]K5�,���c��N���t����32# s�Z]Yy��T^1Ngz��bS�]|$%����HR��;Z�D�p����W5%��+�;x�`��4hD������6�7�·d���m��Q�8`k,�ʭK���}��lk�(�Lqn�ꁦY�u$p¢�_�g#M=JRkF "� �葹��e�lv�11i���6f�G�RP���5�)ۖ�čwG�8�%����⋯�������7�'�raIy�蒚�*V��s�c�ś�(4�����՝����V�&%~�q�)�W��e�j�m���&v	ώ凡�1Sl��8a�q�T�˶�9d�s˟����:J�"SŸ��On�>l�a8����a���I#�rI���Ȥm�gOߒ���v����*�����y�RNCfo,"��}IE�bY��|�tjf�΄N֩�Q�KK{�[f�su���#A�1�O��s�}���ǻg��
�O�Z���C�E���4 *�d�_�|&����L^N�๟��K���^I��U(u5�G"�,��'�\儧�KB�{/���@ݎD�v\�;F���'�BI������p �*��+��D��zg=Q�i8pQ�{˔�M��O��{��s'��%�Z����~��� �H��J�AH5�7�%�2��5��GK�(k���Gdf���3�
�9w:��;~��"X�;Űs�HQ���狹X���,��VCԚ/�>kDHRB�|������i[1�����76_�C}��|�#��j��l����h������|��f�'��hT�$���̟OS���g[`//"�ߨ^�7�_�1&��M�κ�y����yP�^�O/�h�@��Ȯe�4><��=���'V���cZ��,��/8�H)efu"j���[,��i��DAqq.�J��� D�şP��	�>ط��t ��`D�&����֓��PHk��O7F�_[h�X�!.��B 3�@�(7ZB~�B(�8 s�f>F�����}�)�T+E�I�'�fi���S�H�.	p`���~qrY% �k�D뺿}���a;IT/f|���;�Y�z����((C�'m~��M@%�e���`������&�O^�k�Ү�����7���(�A�*$�s�?��^wI	�8��M�?V�*�Q��r���+�(�D�!��[<�+v���.�^���?j�7��I�}#�}T���%3���tjD�ض��B-��q��w���2Ɍ��t�3�_c� &;i��!$�>߼������R"��>�V�_���m��Ʃa�W��_
KP��f¾gd�;�9��l�Ԥ#�0�s��O,�P�5�yԚck�i�"�@���/�[��E���}����0$��)�tBǓ��$\;��!�W���Ϧ٭R����
��i��@������=E7�]>Вx�Y�D2����nt���r�V0�R�2�8�7� ��oeS�Ć~t�#���_�Wj7X�\	�r2�m�n+._�ls���R��+�%����W�>T�ѿ���I,p��b�sa7|�f����dS���Rr��o�64�当~�U-�D�5�md�$�c_�4Q��-t!+����YV�Z"_�[ktr?�*�*Wy��ǉVSYǎ\M��9�C�+�`�9������N/.��*�=<��$�#"鹾s�:�_�n�q0!=Y���J���"�9/}��Ż�{�@J�aw�}��С[]/��B��D]��=)l�!G��7�G�]�����P)K����;f� 5������r���5��l
����\�3���p�y�"�B��~�vt&���]R�L�y���g�=&ώ���עF��h� k/��YP �y� %�����.�~�K��e��z�ْmE�T�%��<m?LJ�[3�T��l�G������j��H_ۃbx�{?	�6Ne��^�6T§*��$�d��N率�r^7X�I}=��8:�g�7������c�j/�(�]�;�gzw7�~�5V����-�6&�ǘ���\�͒��ĹF��0�^Ö;�!��=�8l:x�N�;'0sM�JzǗd* b�%"P��A=T8�C�zS��_�s�lՍ.��A���pa��Pd1Њ�Y+�f�|�P^�t#\a���/�j�k�<"��b1r���ȗ�I�t�w�&�-���w5X8BѬ�o���d�����А�F�]�"��S�p(�f!�Ѯc��#>��c�JS�ɧ��0�0M�x8���7էJb���ޯ妆d��}]��W�G�)T������K|��B�o��z�#�p7yA��0���^�?������˓��3�#���Ѻ����W�y�푅NOp�๟���>͕�c����g߃7f�c�iP������� o_�^���C(�7#�/�cm�%��zŕ�&{3)�OcJ�?&�s��P��њ�Qc���>�Oj���n��eP��(/>ΦΗe�L��v1�lOȿ�Q�6<M)Ļ�$}&��Q^�C��6[����t�q@kY�I(�\V�<F�6���+� �������̤��[��L!+�R����m����ت�����F�aFG��Fp]�����N�ZRr;]p���д(�9Di�����TLbg�E@~���r���yڮ���I�=y\Rs�<U]VW:(�$�����R�&���a�M$Z��N�\!L�U"��]g,�x%�������/�k���n���X����ãK֣�1�h��M�׌�7+��9q�d�xr?Ԝ	t����*Z�q���b��'Lڡ�!oJ{�i1Ҋv�)�VP'(���m
���v����Y�7	��FWZ�x���C5��
	��k,�����ra��6�����^}4����Pű�ۺ	�(b8�
s����]Z�v��E��O&TN����So&c��0R�qơ`Yw1k�EEW���o�M�~G��@#��ۋ,�d��>�NL�*��]%b�*|�rbd2Po5W�����s�MdlG9�;��Bh�a_�i�S�,�w����8wt�P��:���c��*i�l��Oi�;H���i-H�{�od�W̓�;�1��j�@�j�K�Y���B{��:=M[��1ޥ>�,�*1P��1�v\\�/@h-������s��ikL,g<#�q��4��D�$}����`�s�1���{��*�g��Vr�FE,�:è �N}'��1��a|&c:
�w��GU$h�r�E��3��� �)KzW^�̧� ȭ�����B%��3fREw�,OC�{X�\S,����r����疁�E�^��70��&A��k+�IHMQW�iʐ�: 
�s8��S�4��e`����mm�)�1Q�n�i]���*Ҍ�ٙ�58�������`з��ܸ+)�^���f�_K�[�6���FT���IMFX!wٳ�H���sv@�I��Ԫm}�0��qcj&9ݟ]��c��G�ؠ�MoŤG[���֫�]���N�c����^@Z*�'ڻ#$�lY��t~)���\����x�P�{�6����w�R��3�z��_��4�UT�U�9qf0cW�?&�۝��� 5���#���]�-'j��o݈����m�9�]��K��4G=ѭ���IJ-c*�C�%�"�\�|Ь�	�D/.4f�|��M�����܀X8�KwF|��]	B�P L2����koz�=����_����]�ş����G�~��q]��/2-��6�{�ED�wtݍc�J�R �'�zL�d���L\�B��5��mWY������˭]���S�j�N���ƫij�*mG�ǻ�q`tՁ�A��l.~�H�p�5�W+�c���F��3��R�\:l�%R^#@h�X7���OH��W�QC:��<������*";}��%[�/�F��q��wQj�K<^�XrrV�P1�#��@��%���	��=����hS��t��������LO�`��9px�&� ,6�v��_-�ASH��p]��`_o�xX�lfaX��&��� ���<��P&ƃh� ���*�AQ-��]S��_:�l����D���e�u8S�:ȫl��h���+ђ[|�2�S�sإ��I+�J��M��8��J�ùF�WTע۪��7�2�׌;+�����y�֝B��M@T�X:�*ڃJ�j�����`bM31U�P a��=�u��-to��o�Or�]���ʬ��o����$9䊰E+��|���ɭ`�C�	�����a��&�����㒯j�s�xS��]�������	C�����<�S
�i���I�R�%,�3#��;-x��q�e�rě)�*�3m�w_�ʏ<3�������;9Zqwq�$��^ʺ�a�b�4W�Me��0P�1�dǭ��TX�1R?E"��Xo٢��#�jzY >��"���~����3�;��]Lue1q�\�zJ�������迵kg/�Zn��à��׆P��u��K%�<�S[.�#���
�7 w���
����FЬz�`Bςw%l��DP�Ϡ҅����w'��x��X�<d�4G�i��j�P�� �(zs����*q`@�_˯NLc�-~��t���P����Y{�	ǒIGr�ݖ�,qv�Ι��'��T���������e3��@�*�`�1���k0���="���6J� u�w�DZH#ȱ�o��X˳��\�
F!�z���`�`o�2P����ю�h��p��tK�iH�H>��D�To���Bl��)ZS<�D��r��|��6i��Q��
�g��d>b����C�0�g�A�sƌ�_�u,�a{�y.��g��ڟC+h"���Bצx�����N�4��� �8^���m�i��`�<��)I�(����H/ћ"�F�9}gh�B�J�
.G��9�X�y%�'���(��i���P�y����!�d�� &�Sp�Ĥ����	&+>�$	�;����}�:?�<���E�`B7���M�@���*����:g�!nO�T�C�h�^K+"��J��m=u���P�R<F,@ٕ�D��%�ȈG�`r��T�� ���Ih�S��m�)�@	��b��M���3�fy�@	�!6Y22*Պ"l;�l��z�|k�u'�D~�}rN��N]�;)���:+�Im����j���\��$��g��X�P�����`J�7,3ώ��������N-��|y��4�>�!�͂��^]�̩�̙X�~��/�Ғ�j�S��M��3Yy�,����֏w�ՔG�Vs[G&���Fk���n�;ES�dZ�R��M��#v-�,��F���%d��?�ڴ��C���:��j�'�*�ݥ8��U�� ���'�h���(O��۸�^0δ�+;C���l����?�L%ɤ��l�-ó����4���5@�R�B�}
�X�CjEv��iO��/H tY'���ܖ�kf�no���0����y�2�:�u��[�%$2���V�t?,��3k�Yy.7����XI��z)q�N]�9�}�3ym�ì����;�6Aeo� 	y�G�"�������˗��\rF�'
����G蠘w�RVoK�`�e�u�K�|/oy�H�[��J_#��X�����CbG��D.�+�5�X���kK���ڐ]n���sx:	h�T����m���v0mB�|�\���:��Sy^KKY���E���7����f�?�};�*���3�t�W#��?"ר0�	d��z��<4�u����J�ֆM0"�EΙ��q�K��f�&������k���_D�S|a/b�A*� 5S�9����=F�
�yZͥCL�"z��{�%�f���5�@��ȴ�."�}�j>������Z%PnX	�����<mE[��'m��&J�����	��1A��^Eѥ��.�͹��N��6h�����iO���3�=���$�B�����x�v�)oME���f������WR�$K�&݀���]��&��I���3�Y�i����C���+5�r@l�cs�ѹ��H0.�SJ��|B�>�Ygxʚ�bA�f
3[�IR�- �k���ϑ����t��0/2b�G���N�I[�\������,�M���	E$z/�5��U�V3f��
l�p��)&�`�����Y�����F�Q~�c4�&�ѓ�R�A�da�Uaxa�q�&2����(��st�M��k!�S�V��!̄3%%)M/��u�9�$��
����{�أH:<�N>J�
�$��$���}9w, �es{b�aᢠ��xɐ�eA�6d�)�ʝ�.A�������QB9lL�o�����^�;�c+jn�k���R����-�Ha���<4zm�~��M\7D�Nx��;�IЊ$
����{�w:&͙1�k���/�c۹Xw�ff�ʟ��^�������h��=Ћa4N��f�l��̔1;ۖ6<8I\�"�(�x�~��SC4���O�8E�ӏ��d�jе�d�������[m���J��rT^"Hq�1���aN�6pʘ�ݼKw�����PعvJ5��;ȏv7���7����4�,��M%^�Y~�����RTB}�5փ�����������O� �����ű������`�@*��QZ|vy��`��]�|�྄A{�J�q��ޅ�%G�D���E��ݕ�(ׇ#�y�K�<�r�O� ��٘ ��=a�jo�j����Qg��Z�%�6�U�yiZ�v�MM�:j[&���^�X`�<Wu�_��NW3�L�j=���!P�N�u�A����EQo���C���;��s��D��)~2�����&������ORͦ�Vg27����d�"���R�~�_��6ӱ���$�
�4�C�][?�ɟ'��#���F��C�/����`�9�^6���K8�c@R���+�Ւk�bi�.IZ�*8cV%��OE��b���a��c'�WxfC�E��~� ������c�c�lpN�ٍ_9	���7������)/�JQ��&9�����.�@�1�0F
���\d�6(>���&��[�w,��`1�XܩE"��''q �G����=��?Pfv�UM>I(���{�pr�������{�J�3T�3'��yG>�T�TV6��Ƴ��&�e����U����6$N�u\�j,8�jU��+��)���Om����2iS�p࣊��n{�%R��7�q��f/�pO��Ы蓦��h�o�l������;G#,A���_3E�ۚܡ�1c6K�$ 
4�8o.�����:8�y9r
��С1`H6 ���%א��=�b!y��Lݔ��?���c ���0!�0^G�F&��건1���)7 y��:r�dv�N�l�Wu�J{���[ ���B� �s���Y��ꔔz�OK&66X���c��%���W��/�ֶ�U��abh�Ip��WK�s�T����%A�q���N�6�@�'S��׻�1j�v���;V@�� Zy�5	��y\�<�ASI�=��3��E�,����ˬ�h��2;�����2�0���]�XT��~�F<quC:�N ��X�w�w�R�j�$;�I#h����
гpQh^n?��Ө�������O���HW����8�����<G%B�Ԟ�E{�i��~��dP�OkΛ݌��[�S�$B��X`�Mқ! k3�/	~\�E�1b`ɉg\���W�n�a���QYԞNO}T�7����?�zk&����Q�$p�#���(avYx����c��
%ԯ5L��o���c(b�m`@���~�Z�2�Fi�,�J��T����r��4�!c�2�7E��*P�ܙ���h��Fq����3��aE:�Z�I�?
���]��+�����q�qA�� [t̇ߓ '��L�����rcyƞ;H@�Vﴷ�n�~bw
d�a���f��(�꫒�[����O�s���Ih��	_�<�*˄���X��v�N�=�8y�s���Q |��"��8�Z�~��ޡ��g�0����r���]#y�Rb|�_�Zc7��� A*����LlTg��	[�9��N�L�~��c�~#օ�!U�"�u]^���"Pi.��H�����v� ��@b+m�E��N0(�xϮ;�,���t�h@��ËM�H�Z;Pb��Q]A�n��sL�W� ��`4BQG�?z�ʂ�B�G�=Pa�Y�4�g�"�B"> �T��s�H� ���_SݰF:�d��"���Uu��X �$W)3��*I���P 2+�ioÃ�jDD��r��2���!�DԺ9뉈��wݔ����:ך����Pu��k��E��L� 녷��6��5�(p��,XF���I�Q��n�&��9�.��T.�J�mƼ����|���iXvc-���X�j�������QA�
�Xť{`�Ev��E@渦�~���u�3c����+%wþ������WڅfY����CEq�9�uɫx�!���ɯ�a����|�ӪSz
��9j1���A�}S�<�'-�&����{�ӕ�䥁o42g/� ��I�����_�e�ۭ�	b���ɟ��A�?��V����z���0z��w_@�F�V	4 ��3ǖӠ�4��������U~������Y��5E�8��D!�Rf�;�R�2F��7oOK,�y�W�
��2���s�8�\�/��cO�D���x���[�<�Nn��H��^��M������ߔ��5(ż>��:b�����͒B���䂵�SX�N���=4?���艍��n)[$f��އ��,W���E	��*O&���	:hH�χ�P�3ͨ2x��5Rޯ�vT-e9�	�ZT&��A���a�h��ru�>3�dn��>�&[$�E�+ɓ{ip:�8%i0Kd����1XN��o��[肋����-O�Y�����;z���(ҭ�_��^��T��Ű-fP72�%��vK��a:4�qq���?t���\���IiM>2	M/璑w�xx �>@w���r����!k�T6���<�G����=��X -��Sk�2n`ܣͲԎ�t�+?�SǼe���w�t�x�mѼ�7�����7�D� "���B?bO[��Fa�ٌ�T^�IÔ�i��n�8�kM��sO~:6_����*�xT��`�����	{I�O�c�s
�����b���QR\�l�ͩ>C|.�#Dh�9�h�Gs�0	�m���S~��[X\�ka��1�?(3ͫ�Ȳ�(���@J��ƋO���ǎ"�O#)�� {&�emX�{��Sv󛵋/|���H>��1��y�C�������L�,譬ФI�5´��^G�F� _�~
Q�}&h��̡f18�f���X�����_���eN�k��8h�L�'�H	��j�]�Ju����ܑ��o�=~���L���t'q��ߧA��}�m^2��:����0�rd�^�r��ߢ]��?��hh��6�5��RM�`X�|�DHR ����ә�b��Q���ƣ��'gxt��w����gs/iD�۸�U#��q0����<� v1ۨ�h.��友�\[�4��H�����KկW�-�$1�ˤ�q������d��|1��+3i���6��'l�@`�jF>=��+�xf3]����h�N����%�XVa�U���I����m��������ߧ	.�p�0�hȘ?7�sx�wU�'�r
�Q2��&�gOA����w�������^�X�@k,1�]�1n��"�C{2*h�P�v�5�.f���@�-ۄ�)�(�xU�x�'���c�m���ܺ\��o�#�'�\�9{�����1�>����[(��1�-��_^��:86k,~9��5�?P����zu:\�� �x����_�Ǵ1T
�KJ/�yՕl���&��'��s�Q6ǟ��3ǣD���ej�^��1gz�v+��{�?�&�U�-�/@�pL��ė��	��"��{�?�u&�:1O�N�^֥]rn��� #���z�c1I���w|�\�E�
�Q�$)����`�;,�����iR��Yo�F'V��9E�Jxq`EIH��p؅�,)Ӎ�Pj�ǽO�V�S�R�!$�v�a��L1^�^#�w�G�[�Q3�y/��Wx��3����Y��h̏��Go��N��O����#v�9l�0;�d���� O�DּD�655^�8[�ފa5d���b׉���]i	5����4ks{ʦљ\@��7]'=l�c!�P��
ك��a&�Y�j��}����8.��V�[{��-S��q�7����|�-R�y��ᾀ/�ҿ��#�{āT��<ݧB���@���jro.�u�-s0��Ꝙ̾(QO*{���Iߣ>�%"�A��,m)��ĲW�ݺEV�x-=Mvx�&"�h
ʘ3U�����q_�Yu�&)�Q���.XU$��@	C�#HE�&��!c	�R[qlJB	�ؽ *N2�h	�Ux��F\05=��A�(�tCj}y���_�?���M���/¬��U�
#ƂW��Kv�4�b��o6�>���!N�2|@;���Շ�g��E�p�L����G �h�Mզ�Mǚ�75�Z�N=HF���$}�osu)P��ؠE8{%�.��af����?�3xkl�1���eB�e�)?���ǧb��V��:\M���0���|�'=�����:]Up���G|�@O-oy�����·�b�b
�f�$- ���g��rO`�Ņc��B(�,֜}F�x����i�,���p���'^S�pպ����}գ���������1Ș���O�fSa��*�z-�d�$ d��8͵-���!, ��Ơ��Sn��hꪝ�Љ��Ԝ�_ �Mm�O��n5]T�	��*ݣ�+VF}at�m�q$������v�5��Ԇ���<Ί%�)�Z��~I��tu��ʐ�;��0Yf������X7'�
q{��|�w9i��^��+�E�i����]��P�y�VF�ʁ!�6�{�K���i�Y��t���1�`��Lϵ@��NV�������#��/����2}P.�[| ����MG~:ݭu�q^��yI��ŭ�@uqZՁLJ�y0�q�|��b3��������@,wz;
�Ql���.sݔ�ʉ�R�ͱ����
h�ӝ���4�B$���Mm*���R�A�S4��li�8b��UN�a\g1/�A�FE���yy2ϖ���t��ˑɋ���*�Qb32Q�ʕvD�W�n���9[��9(��;��Iz�YH?Z��!Bt=��Pv�`{�Ո�qB璖�ǭL��#6t�=�YO4��.%�u�M�0��;�C}ə��2�3W�`���_���9�,S�_����8��a����gI�]�Y	4����'M�s�����E
8k�.���X__�}��
-9$T"�����=ꯂ�ܨ�|"Ż�G�rYp#>xUu��
H�����Żg�rރ�k�o�%��u�̞�`Jg�L��=�%�g�l��ɂ�ew��y���~#>�kN�3�>��f���#�bt� ��I�l���� ���:�z�[ӌ��و }�����$��!>�YI���N h��"��P?W]����8��x����&5Z��u+���� I~4r���S%�����"�XCGc61u3
T�c���u�d�@�J��\)(L�?�0D]�ܶM�d�5�B�0KO��n�(v��S����gt�~n����#ʧ��F�,�pe��~�-�xm�_��
�R�i��vP>����XN���r�÷\!�U���h����FH�(��f3��@Z�i����d�^��[�4��8�'w���] �=����쮶
�� �]v;������4��\�sJ�nY�1�~��,�qJ
It�S쁝��e8��m*�L�$x���X�,�Y�.T#�μ�Ki�Q95��t;��m�:�j�R��,r"K�T$O�t�B�.��� �ƴ��|��� S-]�D�̟�潻�N��P�����L�pM�1�4����p�sg��_�"JĊ�~�!���������26A�V7���B����H͌��"���
B.<�W�,x��yn�i�'@��X��Ϫ�������{���f!�r���K�@�v@@&��m�~���m!���<��ɢ�o�t�_L�~}���(\�u�o�Ҫ8/�$
�Ꝡh
��z>3RSM
7����8$�鄟~04�A~�7�$��m�o[f��&�K�a�1�&a��3(��V���f�`[���� k�Ȭ�3}������0��� dؤk��Ld3~���S�j�
�T��5�Z](�M��)A�|��g��|F��W��jCx�2���[tP�~�P2��a�U@4�CHQ����1*�Y�D��((�E���y�^�T���q�7C�Ѳ���^ld�t��@��>����$Ȗ�c��OlQ�6�YN_,��i����9�� �K�����N� �ԟ)eM2���&�#��.ļܱ,�7ip�m�$97ó!��=�}GB�E�x�{�U�e���W|\�$a��_��[�n�~�(>Ů!P@��Zl7��$�
�
=����g׳`�e͵�[geL�4���ڊ��5��g���C'��,��=�i��I�(�^ZE�+�˝�>�ݹ�?��Y��r��6��R���]��F��5�h�@A�����p���`�T��Z�4��FşQ�ɀYzF�KB����t���n8��\�ʙ��f~C��j��V�u��Krw��8�[(XD:ܫ�<- ��#�dM��AK�ǳ���Al-{1z�}�i@�� ?�p38U���W���b�`�7}�[�Mg��k���#�/Ml�>V�l]Nx�^rF�g�}�`Z�LY���ͬ�)y�[�����*�U�7�OC������8ui8s�n���w���}�5�[1 
w��ěo�n��i�b�#���3��ÊKQ��[>����䈸��	M�1�tD�{\�i�Ѻ�
�y�!]�;0����"c�qZ�a�ۉ���h����ʐ!\�v��<�V�T�J9��oi�=|���j �3b�~E����Q�A��z���/+蔶�̈́�/��tZ�wͫ���f�=O7\:EU��X�<sX�O=I�o�1uvH!��Q��+r����'�ճ�v�t��%� 8���B �\��}�N����\�c�����
SV���f��t̳�+��O�wLq���ck�'w�9d��!,��jd�h��S�Q"�������O�#0�5��� �	�qB�
4�������8�}0���)��^;��	���I%�Μ+]�1~#6��%	.�Y1���S���+���Ȥ�M#�J?/������_~���E�O�2m�F�/)+e"�����iP3 ҬD"�tii7�t������E�q�O��߱*�GNż��i�]���ɶ��������t(W���j�.�XK����پ����X|l7�p�� }ɾ`�I�H��~��E�B9�/�7{���TG"��{���L�8̦�J!㳪Vz�7����f3��Ƥ��,�d��Q>HV� ��*c�& ��$<��b1!M���%
p,}	��~��qۑ-��&ŪX%cSK]��h���+ImӰ��w)O��V�#��_�Ϙ��W`,�t�Ůɉ!��V�3�.����o�A����ѯRg�!�ˉp���D�w���)�F d��G1G�1Qgwa/(�e�u�%_���\�{W�QkEs�,��fW��짊u��ha�i�.���^�KCأ:���Q��cof/0~~�����}u�e�L�(��AQ�e��?����N'���a���n���]x���n�SC]ԁ���Ql�bJ�ր
�#*�w��e��`P��Ņ�����{���6kByi�tD��]	Ym%����x�Ԭ�
�vl��Q0�4�"7y��ӻ��̡��fT%g��М�*��"�+��+��FP �C���M����x����	8f=8K��\�X����|��lϹ�9�4��k�u?��;�?(ү;��p���%Z�+�t�],�`��*�]o�ou�L����&��g.��igd�@�sW�shc3�x()v(=8H1+�m�����|M�}ywҭn�؍�grnc�]�]i�wc�����"�Y-n�7�T��id��(��&��gt���_v�{/��}�RF���87�L���4�gJ�o=�N�A���J�R�aQ�����:m�և�m̯��T�ZC�ZKH�wn.��=Q��0{J�F�|���Q(���=���&#��\��B㕄�T2O+�J^^�vŹ�Z]���G~&�K"����y<��-����G����M�<	�|���-�:u ��d�~��&K+y�F��2|k�F@�=Fp�N�B�<��b<Pm�>dLӯ�q��!��{��/V�4��mHM$@��I;�<��q�[ϱ<��@CK��d�(�Y�a��T��w�Y��O� {Ą04���I1S"|�4�4귱Um ��zTƋP��y=�pu���*ш���r��������̈���>D(	'��e�2!�~Y4��չ\�o�	�j��{_����K�*[x���P��RUE� k��a�:��
�>Q�^��CBf�c�wG��}H7��+�`�&D��@��:ٓ���H tSi����Ei�穢�i�,�Y����-���+�=ŵܻ{ �'ME�K�p#~��)�6�����^wc;�5��r�C��� ��>�o��R�/��rx��	%h�N��]Ս�6W�1R���A��!%�����c(ڀ��� �M��o��S�����,�g�ܶځ��|lS�,
e.�<t�Y���K=\LB�%A�z����V�i`�q&�y�B4,|p��,"���^�h\�s6��պ�i��ڌ�?�v�ss<��X�?c8G�E*ރ�pJ ������O\n�T6{Y�A��Z}:�Hъ���s��e	͍�����}�K��w3�@�q�Dc㲳^�2�Jc#3g"����U&w�W����I��e�O�y�D�{��V��H�t�H��|I�Z9"���X�3+�t%�p�X�8�$�cee��.+��7�W`ɒ0=��
�7m=�������D��F;F^����#���Y'u5�����՜�Yr`s}���]:ʛ�{����r�E�m�oz�����nz�^�Ul�R\I{��0��)s���[� ���'��4�Ȗ4��d�6����p&�_#��G���B���=y�&�-��eH���2[ �?z�ô�5��M��Py־�Hn��N���k����G1�)��ồ��u�nU����ܨ%C��4O7�
a��w�t��7#�fn0���6^�{L��|=~�5�?Q^����υ� ���:\��D��#��\�v���S�!"����Cbnsz
R^��fʇ	�',,{��������(h��,]�֯���]´��B��0��DU7 ��D�v\l�R4M�ۀH[���0#=��Ҁc�6	pG-v~�e�ן:�Sj����o01��?f�w�����!�E5������Ug��od�),4��ɝ�>Đ��|�w��r�jik�
h�z�F�g�*�tGSR����/��,'?�Y-w�����ޱ1��(���Y��t�ޭ��stw J�b����v�-�(�}��t&{ss�z�oZ&���\j�m	2��F#N��xt��W�5�)�|l�Ki'��ԕQl�ÖdR�P>�����O(sz�ITw�u�T���&	U��P�S��K��U|{��D��(��9Õ4�k8>��Ǐ@iPB`�/!HW7:�)L�k!E���n�o$�5ʵ� �s1-��_C��#�؆>��/�?���6Zt)�e����9:fg�yR��BjdO�m��}�Ɣ
Ѝ��g���i�de��;8�	�uPrƀ<CS��#o�h��5K�>���PqԚ���H�Y)c�Kf0�L�,��� �jD�������T�?Lc���]> /MBG�جXԉ���,� y��t^g�xLc)��)����`T���-ض�����rK��WK��ŧs74����KErf��?ɷ�?�ԙA -�{��/�X�O��F
�k	��G�O�����D/ץ$��x��H&	�����(�E�(Z��� ��E��m'a}���:��x�.�4%�
Vx�.�2Y�B�	��fI��ZJ�Bi��ǀ��I �TNg�A��jշ��E)�p�\�H��D䏯xͼ�o��a�k��k
9 �Gny�r@�_�k�ӵ�Fʸ,i���l��E��'��R��A^SY�"n�Du���)(�g�k-R�Ah��/���^�i@�D2g�Ժ����w�{�����U�������!\$�������A~W�5�kO1;Y)�E���d�H�3�0�
���?w9ͭ�\��5\����s�ƛ�[k��McX�&�mt9�5 �4�ƳG�"�a�.�p�e��KG�y�;V��v�v��tE7$�&��-���Ò="��n)\�Ҩ[T-)����J�:q% �)JaKÅ��>"*J�z�=;�뗲�mG�9���@�t�XX�s��j��0܇����"ȭ/J��r�f�����n8��`%7�k|C���}�V�<��b=���dLW����O��f����z��IxG�̙Ψ�S�H)�fҩ�<`{����k��	���&	z�=��U��&��f'��p��A5#}u������&�ޖD�"�K��&@?���g�Fc:V�P�Pg3���?��dH};�\���4#�����_&8˱
R]���~ԩħ��	ӜJ��)�\ƺ. ���R�u��,,D� 0���C����L�ѩ�>[�`�o�>��ǹl�0�rdjp�MG�dw��(�*�s\��n�� �"oSL����ˤ���q7��k�P�����?8�9g�Z/8�iBG�����w��q	��r~����x�ۢ�N�]z�ݐ��h�^@v7�Mb��U�ּ�f��	��SyCK�R�X�ӗIM:\޺m|	Ї��aA&zbt��彀:f�u6�K*��w����Yz�KP���u�X���W�z�P���;C�4�Ly�f5�+�/���B�a_� ��#��|S�D#:�)�_��5���-�dN�u�$�c!�9x�4Ƥ oXh�l������ k/6m;��HR�ɫ�0��s���"s�;���:E=���M����|9c6�Jl�W��eL����:Ż���ބ���<g`PG�exDn���i�᝗
@��מL5���cdK>CrG��Ϟ �?�~��Cy�=�I�1�}�hR%������к/�ʖ�3���l����N)P�X��VP�S�PRa=�0K|0��#�&fa__�t8��}*/�4��o2���C�����P`4�;��k�m�u���m_�ec�N'��X�i���%�K���RBv)&Z��)�,A�}�wԽt�����l��;�u�c,��*�U=r�;�o�9��>��(���(>V�)r���<a(5LB� �{���~H�� �7ry��(/[��@���c�M�lAQ���|r|jA�%C;��JBW���Sb��3z�P�V��I9E����C=~ �qpM��r7�F:��ʯ�Y#e��'��o�*��r�o�X���?P����%u���h�GV�1tB0hB�f��l�Ln�T"�=p�Ws�.��_������
��g@]�Y5�:x,-�� o|��[��F|b�
�q�[�1?���������s��psS�d�	[_���Ep�O9P�F����oț�������rz�wW]Ќ�Y�r4��/��jm(e��uf[8iSt�'�.�uF��^���K,�Px��@e@����{�%�P2�ZA�`o��D��6��1���bZZ�I��$���&��Hŷ�P(�,k��wF��]1s�dj�,�L�%[_)�Mh�(���\��閵��������l������)�C-����Z��c���h���H'ɶ��s4���w�V���i�7/1\_�_gu^[��V&�;ｬg�]��9F~$,U_�{0�v��v�:L|pt��Q@��"�U�c�?ħ(!6�Ϥ��z'�{j�8����4��+K�q�͛�d/=�%��D�G^�0��8��v��7��/l9�!_�%���Jk��5I�}Bgc��f	A�EK /W0m�?�l����-ĵu�#�	�$��<S',����	[J�vv�����!{����"����) �K��Z��Ś�#{ �l��;��)G-lǁ��������p����d���5�e�'Vŉ?5!_=��a2�Z�bn�7,�ל�J��\bH��Hb'�x�|њ�>U"�R�"јp���<���S��t����$�vS;uxVSfHSJd����J��..���,�|�v@E_����S��e%~79Y�zb�D���ٺ�%=����&�=�W�j��d%K���$R����\��E3�?�=�cz��:o��JA6V�T9g�V��CZ�<x;2���9��j"�M�0Hǐ�af�h�,i�=�P\g�܍�A�����f	sWu��֪��r����|����e�β+j���{��厡O�]tǆ+0�آ� ��=g����c}ތ�has���Wߒ����0J��{�X���̌��L6�nN�Եk*�&՛�yf�D%�~}��8�%⽏4�YΗ쩗<��V����)������o� D��s�AF�@�=,��*��Ev�2��dݻ7�+4?��83CČ7��ZB��8<���`�k��(��e]�>&FN(@�,W�Ji�� ��KZZ_��%6Ǹ�����,ˤ�B����������-�S�g�l�'�9�0�s��Ңf����8�妝�� е��L{Q�O�c���%;�Mt�%��A��պ2�Ȗn�}�'W@P>�e���(�Ꮻ�Nq! o�
xFr�:#<ZڑsϾy­Ce��:�ׇhJ+�u���Y��Gx��4�QR��V�U�B��>h�f��TIP��\�ݓ���>��1���a֤�48]�������Ht���|c,&t�zk����x�Y��>$����p�e�*�R;���D�6�]��Q:�کԽ��	b���f( ����aF��lzze;X�&$Mj�(��Oػ��y��ő�ɾ�v阪Qs�,�a�r��Nj6�̨�&:�m!��{%�r�n���F5�����H ��]�	fL�w�r19w�����^ZiI�G�,ū��J��R1���Q���=>�4Y�,��G�ڸ��3q���������5��_]M-[�+�� �YD��~$��
���Y?ذ���@/g�|!�7��Uc�{���R�1�hd����3l�ɟ���I�W�頫�~������|ȫ l~���F��ߖ'U�4J>���MPB�y�|X�̨>�d$�B��ڱ(-������g����:i�D�,�0H���VĨ�}M�!d2�6��p�w�7[(��uy!�ܳ���t�[9xM�d�|ҋ��˚� e@g�ܜ�fz9�"�MPԋ��
�uyi�=tR�|/o����P�Ԗ��� ����K|�=��.b�\?�M
�"$q�;�驑���:����!� �@��F'�@���>�)մ�W�2wa.��2�l_�ԝ4n��H�~�ֿ�p�`k1�M��?�5Y1��Ƈ��Ȧ�=�ä�X#3��8\�u��x؈;�l2�R�fV-�	e����+�nL�[W�8B�,v	х�a��h��	���D��w6�R�n|�,�}fX���m��]wB]:�N��,�,Q�{YUO:����X��C��߾��=�Y�5�߱��Y��e,���{HHO��3�h��V��E1��u��cM٤��#|2M���+�Oe@4��sʬ���Y|���guxg���ѿ��h˷Й��l"J��m�$y�`Hw!W���x��=[j��O���{�j��<~sq�e�h�P~��iI�9�Z<D�W�؍ luzYN�LyjnH�,�RCc$a�?>�C�'�N4#\-�C ?��}V�l�#3�t �.��
NpU=�X���T+����ؕ�]�sx�t� })��u>W��+���\S1*��&x�7Y�r�Cu��p5a�p��G����\��_��'��K�番��$�"�j��Ԝ�`���4�/�д���U��*�h��A�t3�jO~����ol�+��Ը����hK%f�*@-�j�H�A,]�-U`�M$_�L�6��ô��{��h�X�����-������^�m{�'FJm5߸����?����"�D�y�d��(&����V~7�5��!؟�Z9��r��u�����d��G��fu,?!�S��Q{���K�X��1Tw��a���&a�o��%8���rs����$*>�-\�H��
����c��mc�����:�FQxƯ�}�O�n8fcHk/�={��ܘ�Vnd���P���7�\j]�h˸����lܛ5�m��wR����#���F,ݠ�ߙ��	6�~��!��7���<5 �M���m��B�!�R ��FpJ�s̨�iQ~u��*�&i+���o�Ry�y��en�ޅ���������H*2Á%�|�E�ç0�9@�sR� {9ky�T����/�tx��)�vI}�$B!<�vQh�k���4yp?p^_AV.���>��\��l�����A[���$�����M�Ͻ�&�}���	��8x�@�6N1_z�RY3����BڽJ"�L$��'C��ˊ¹�m���֭���f�E�w��sm ��K�%����=����	��y�O)[#|��}G�<��C���R��-����5<���.?�/P�._����"��f<��"D��n��,`�Uέj\�f����l�$n�@�iVP��gm��D�eg��OĒ۞J}�w�S��]�b8��"�����|�x��hg`�����X����z[�=Kʵ`���A��o��gRƨ˖�X��/R�c�P?ӊop!��b�����I�5�+B\��$��?�i�ZYV��Q|S4�9���"��p֖g�P.�6�d����	1ؓN]���¸�>µ�#,]=���7��+ߒ�cKO16e:�WB�� e�i0'@��̥R��"���y5K��S��#�M+�e�έ��<Q��,'v��w)�PK�މu��+�zh�17������Ng�,�2ZH�l�A��������(̱�H�Dp����Y��+���[
�)�^��qY�ɂm�-��OTl�IK�'D��ϵjk�F��2ه���Ŧf��e=��(X��+n�Xy��Yzԇ�����½~�ܼ�w����+0p�<��Rr ,�Q��o�8i���M��& Ph���Ȏ�br��1��p΅�������<^<3ē�ⅆO�GH^䉩mOF$��%�x���{���Z��D&��t~S5�7dIq@x�bH�Kv�0�H.4b}������GS
�XSz��(0�-fEY'ZpfF��M3��8���\N�s��%���g(�^Q�tx1
���y��!��G	�[���?پ��dp=�
a�ef�s����?r�?���Z0�L�y�����t��SA���D�3���X������$��V��gu�搥�l�(�'�$�u|ʓy�ò���{�&����,�I�4h*���A��VdT�.���j+�a��o7�'TWXٚ Q-�5��v�P=G����j;cPT��z�҇R�
z`���Y諒��M���74�Z��(�H�)���=\{�R�z�d���L�މ�3<�<S軀m)�ɜ��Vtl̽��:i-Xc_=EV0��a���	�43zt;5��ݩ"��,囎��4��{����@���V:�OH`Ѹl�J_{Wm����VV��{|c�Z�hR��̡垗��a��vI)��y�7~_�-2��	�0�m���ǒ*�֮ wf~B8!/���F���	^�S�T�j�?a���f)@��m1Gr�0]�x�v�����E&���w)�'���O�hm�e=�iN�i�	wV4��6������
��eC��>߻����'����@��8��ؐ����O�q��+�(߈���x!��ÿ�vN�#%ֿD$��s�p#\	B*������8����(��T_O�*��,�L_�ɝ'��ǃ���0��+z
F�lpp��6[xI���λ��O�Hof��X�`u���}{Mf�Ԕn�0v��f���*���c��3���z�0}Ce\&��<s�F���"Cw��U)�jT��m&��X9�j�-}i�oŗz�Ҥ�Ҥ3=�דmAE�w����ά��+@�����n٠��.챾����4�7��e�۬T�!��+b`F1���ġ�T)�X����ŀ_�KJק뎘M�6,/Z��i$���00D��G�.=� ��P��Wg��;&*������ �V�<�Ѿ��菮�`�iʭ��	��S�a}�>��V�f������Y3�OǺ$��8��鿌��E��H|Cf��T��Nq�6���**XH֟�A���^������(�t4��:�|]q3' �+'9�f�\���]_E�����W�	3�kY�m�� 5�˚hy�f��"�j_s��S��c�u���|���68��gO�&��+��o�
�A����q8�cxw�9��PAGJ���9�F�T�e���ʽ�D-4x���gDC� Q4��%����VA'���YdF*��~AO�rsﵻ��=��L���)��)�(N�3��a����_Ej�\y�$x� �[���Pkl�kϷ�BNc�o$?�Z�� �H�͢>�ml��gvN��3�^�5���5���K���HXZ�d	��O�D��\��( Ĕ�Wi¥).��5`� w�b�$�{�"kj�"/����������,*Hle�0�Q��{�v9���Wj!�q�bִ?o✏��d�������y�TTpLI4�1��=lN�ȥ)���HT �/H{t�a��0�I�>�"�I�Y�q�x
�y94�L��
K�0S�ܱ`��-1�t���1* "��	�q����x� ��� �_ ٸZ)��Г�NE��{���-�z�v�|?+A����<���d��'Z�iy�P'5��j�Q������iǩ1?c�[�U��ꬌ�ו\�ùYh��2��	�>��I�0.\X}��QZ���m;�T2V]��J��G��VH���&��a-�5\�:E�tv>S�Z4<�!O��z2bHk�@�P�.u�����'�<ƒi���Q6�j�ԭ��u.A�%T���|M���t�e�/(���߁�:�tH�i��F'pv+뎌�5�l�'���b��K�|�?bX �r�h�kB[>�d@���&A EN��m}�0&��� #KyJqV��� 1��1�}����ʙ�8s���=�<�ڀ�c�Бʲ��I���2i��er�"�.	mpL���剢��~_�8hꈚi��N-/D�.�g��(n�r�Q1�T�����a&�3���'�C��2,b�Q)4�X�0��!�z߇��,n�8]bEcf�_��Z��yg_[��y�o0)���=�j��'8�`�A�e�� i�5���򽬥X�!7��zop+�1�06G���ay��˪`��ѦF�����܏E}�d}��N2xr�cT}2aN�S6��k6 ���G��#�1U��FxɄ�����u���PO{p7٤V �'��}��}��F6������߾��3bݫ�}1�i��7��o\ͅ��o`���gӇՄ�[Z��5ʫ�Mw7BDR���Q�лk���&`q�M�s��|�;U1�|f�+0���r87nV �Y��5�va���<�I,�T//L�/t:�k[ɽ��9�%KvJ��U��*P�:�T(�S�DF�$y*=FK����G������K��q���#�e�(~V�f<9��#`N�\O�[���nB�E�- ��P��Y�#"�}���fU��s�{X�O�
��^bud� �hb���&���z�Ĵgu!A$��R����lX!>+<��kb_�hͲ$wz�.���LR���C�8��Nh�;�'��F	w��sl� qJ��N�?�tIB� ��y�J_���\L&�;^�������>�DO��bl��,y6�T{����V�Y�G5F��/L��Gi��ˤPX0j�WP�D���(�+���(��B��7�a�T�ii�L˸��@���8�޿�<�R�^��/ס�V��)��Wh�z�����-��9�̖3Q��;��+�m_�"ND}X>�/u����]�H��}c��2�P&�G+��Y� �X18������T��$�I���bf��U����X}$��G�0ԛT�s�A��>F��pgz�qă�N����O%���r���"��,0꧄�X'�ӝ%�8�N-����]rYs��Xa�� #�̄�'��Z�w��ҳ�X�A IL�����[x�YfF��ܱ˼AX�:�i_��i��y�`�Un�K�Pؓ�@M����4ET̐���`����xc5�-_��պ%�1հ:�%^�5���b��C�Vȉy­iz�B�����2���=���I��7Tpx.(���Y� r�쩙����~V��x�aGv5�!�7�.7�рy��
ِ+��BX��MHθ���Š��n~���U�D|�og����nv��L���9��ո*r���	oh?��7�8��U���|i�{=�Wu
�aٰu�({��M6���l��p�.�7�&�������-��$Cb�<�4j�U�B�7N��g�\�����;-�SA��
Z�d��Dr�KD��|�7u��N���8J�����[r�=8T������������b�ڦ��7���:�x��I���&�����U��}/(/)@�B�٬�w�:c���lSYC�S�$�f|`�eͣD�E-�|R� 7�$�;i����.}�˭�oz��#���w�������_�!^�'G�ũ���r�)%6�S�D�[�t�&`5� �E
[�ɾ�HzV��D�Bl��?y�9pz�N|[��{uu�C��	��.��ͭH�}p5�Y\[3�k�v69��`������w�(���Xg4��༅k�p����?I+�B6�b�pEg_��Mt"|�;+�l~�L��B���ԭ_�lWL4_6Ԇn�C��*% ����0Ik7K
��L���(§�k��\*3����d�Ǜ�i"�0��H�����_�|+�!��?!�_t���׋�q��@f����5�_d�ۭ(}A��]� ������qV�Z�o�����&<*��qüå�b�5X$?l��xo�D�[(Ie�i���-Q,�mB�H��[�p+u0d"qV��Q�~���k]�SĒ�����D�F���[�4��&�p40Iɟ2]�fG��ٕ,�����@at��:��0$��P���D?Ӗ�GN]5H\k�J��݊t��z	��6]�����8�7]=��,#�%Ij0>��g����{�:�����/��Ip�x������q�(b���g�GiΖ$ҨS�P�&`�o��(,�ʟ��%c3MI%��>��e�2r�7�����e�ȴ8�(Oo�]D� �ӗ�p�i�R��(H�SA'��Sxi3�@sd��0�W��5qx]Wcъe/�:��f	�Y�y!��������@>�Њ�s  C+p*%��Х˅��ri���ʹ~<d{i�y�z��ۚ�l*�ZN���Ë�eq�8��YǪ�� {�|�bW�
�k����.����;f�@9���F���3r4T��v�����0F�$b��h)j����}M0�eT��;p�h��Ex���l����긇=�^y��C3Zݹ���Eݗ�@��%uY%�N�yV�2[��u�l�s2B��@�b��+$��D���j2�w�h6�餠�y=��pur�:���	�,���^'�ٯ���I�:=T5G��ϲ/ҧ�V�R�W���
dt���!�������+CО��,�5&�"��t5��$M����Y���jX$��P!�ai�Q��>~�߁	��u�H�����gyF�����/p%�/J�*T}~��݂���%<���_���j�u��z1(-w�[�އ���N�78���yA��t��*f��Ll;��3Aүg��}%��օq�, t�V���`�1��b�Ҝ/��(@�����3o.?�(�-�=Ԫ�����������\>,6�D	Z�r/
�hR���;,bΤ�)3�t�vr�M���{7����ʨ�J������U~h_��d�2�����D�����`.�%(����вߩ� �������(ȭ��%��sd�� З�����S#����	��7�r�u�N5 Pd��s,4��K:��,4���_� ����4�����JKϣ�R�WPx���̉o�7[�r���^����;�u1_�"�g�0��i��k3�Q��1�p�,�3�ž|S�̛�V�}t`�96A�ZlC�!�M����>SX�M�,�"S��9q��]��&�����IX�լ�2�f8GK�����DK�Y�a��?���H��=��_[�x
G:����_�?�v(�$�Jް�%p��J- ֨�(=��]ؒ����_)��9�c��D�Ea�٘�.�h&�A���MMye�Gy?��/`�ywH{�H!�v%Id�����[	����sxi�q��z��$$m�(9â�E7�Fh�4��:��,��z���gK�9����G�Ξ���&� WSv+S͛ ��妈�]���GQ*�{Ԡ�y�D�,,IE�c8��~�Tm6��1����V�����z��"w��r��׬��y�n:�ơRVi�$D�f�+B�����-��H�y��!4,�;[�BD�o�ߔ�թsoi��^><����5Z��/��ũ�L�����>��
���!�G] ڟy-{��n�����ؒ�ZVt:�Z�T.�F2�cCwv�����87���?���:��iG�g��*��L�����O�bu94Rѽ����I�1���a5��T��	�b�6�	��n�e�_��a���?`!��$�^���^�������e��gz����(��~AAr�sJ�Xz`�E�;k��p�� ��\*j�=
��н��8gk��2�/L����q��� 2䎰Ɨ�����V�+�����ީ�^����_�'_���r����Es�lUL���鬺��ʽm�Q;��[�3&>[��e������6=����*^��M�V�g�J�N���Td�[C�)I\ ��P���nn&,erB���/���(@��ѥ|E}�0�<vǩ��p�Zjb�ݴ]b(���<]z��h�A���cp��

6��"7�����������<k^�C��Y��+4ųŽ���4p�0�jޫ�K}��mG���b��bC���`�hY嗔Ѭ������h�wh��8�� �;�ps��A�.B �g�g��u�H�:hƈ�K���cl�$�����IcF:\7M��p[������6��{$}���^l����@����,�|�I��
j�F�rrK�F~�<�W0�ѣSk9�d%��/͏@H��2B�Ś(�֫�W������>H��-^�
��-s�1|���}@$kN���ة�}����D��RS�Ep�Շ��No�6��g�� �R��݆��p{�'%�RZ	�?�BvQ�+n��?�<�S�H�-t���J�-Ҵv=Y�i�EC1[�*���X�2&#�#}��*�0�0��ӳO��A�)8S�i���B[n���!R<�eq�
�j �!��:��'s1#ˣ�L����Vd�O�ҸX�CS6�ˑaL�NwT�ʖ!��յ��!�:�h��6�(��K��ذթ�!�����`I'�!2Y��_d���(Q��_��z��E<B���~�۝����]Ru��&F��ˢ2��o�Tk��t���VD�X"���%� ���yN$�d+8Q���.�H��vi��VS5����q, �'�9��]�7O�sNs0��$U���ɏ:�c舊A�B2���E��Ձ������R{yfZ#���xO��������KR���b�j�	���iH���Rɮ����
�����^�)��p�W��gk��}!�h�(Ls��+�T����M�t6��C�=��5zqj���u����5�K��k�3���3EӚl�iU�%X�+�hQx��D��E<��In��9�� �u�b��f�k��ʋ���Si�z{WDQS��H��Rp �o/����U<��'�R~~_]�S���U�+��Xv����m��S�	�c#-���; ��|��4fe��e;�p�̔���5��Y5�'���v�t�:���K� �a�ή��z�iO��~��:>�c��|��8�|S�����u�Z�JG�u>��t�֊kȐ����gu#���pk$��7��/s�e��A4�z��}�VJ@c��{�Y�P��ž��,����ד ݲ���0�"Zkd�ʲ�)��vҢ��5�
�l&�R�E�c�P���J�L!�E$�'�.��@W����e�S�K }M���0W�b��[�q'#
TƷ
c�%�+���Y�d��j�� �&sh@_W���2�����/���O���<�&ּe��C'm_�*S�.�,��5j'�U�D��u.�/3@���v�Nz��+�ۥ:lln��&z��
+2F,I� R^[��T�:����T���Ҏs�����B��:�Ӯ���A}1I�Si�N�V��) r�kj�@��s���{��zɰ����BCY�
�uj�8��'E1������s������~���[�\��s�G3߸w�4�U]ַ�e��2�G�i�����6�o%jVl����_(d����A'���5�뫵@ڑ
�Y�~%�p��H�w�PN�/$v�8��Ì�T�e�`�v|pp�%���P+�긆�C�t���'�} _g�<���5̪o����q˸��Hz]���܎�Y3��}��!|� ��a��/D=�.���6q>5K(�,n%#kf��X@H���mg��ii-�e�����&w���#�$��ʅ3�)J��Y�AnI��%��Tm�\T=z_��6x�&���&ȇ��6ٖ(L7��Ԑ��T����f��]p� :(p��\�a< ���gP97�8�ܾĉZF.�����(,��� �l=���x�v~�X}�7����8|ov�>�tΏ[,��vh�|n�g@V����M깯=V3�&����G��I��ٺ�k��i���w2OQd�D��{����5�":Yft�@ݩ�+����V�<�8��"��t�-p�HJ���$qz5%YI���7�c������>�D���1l @���y�{F:04-������b��!�hT�\���.�4���'Φe��-�/Ca��_���"cÐ��+���Il����8�W���6c�R<�P�1�<c:�c��3�w���(�Þ�Rc��Fr|��b�Ā3:w��5n��Ξ�>B~J�_r,�'��t�ڠHNR��K�pE��&w%]2iUWR��j�KX�"�'ϥ�s����!���^*��0l/iO>g��o.�ۡ�٠�
�g �\��A���AQ�U�+X���v(�*HE�t�o��Ub+
�t���O��G5��4��c��1�6�5v�Cm˸$[u�������:����'~�,��R2K��s{*�V���sV�7���4�iaSfq�(S���#�u�{<�3��Pe:�k��1�%� �CM���q�w�[���#�rT�j���8]�k�K�ˢΞ�z���cS��5W�PIdS�l�j]�+cs%�HD=�ĶL�!��e���KP�f��f�������*�!�JN�0��Tң���rߛb/b�}�!Bj	�An�N�RDͼ�q|��n6!/bֲЈD��2��"�e7���!q
��,�$����.W�ҙ�p�]�d�l�ܾڪ�=.�)L����a3I��ZaH��	d�z�丈��z�׺�6S|s㡛�1���� =e�G4�7��8�5-O�v����x��e��V~s�I����R�_`�>u��0��g���d�ߏ($������7#k�a�$��Q�J堶%!�m��T	 <4����b���M�� ��/�rK�
�ܻ5$x����>ӉT��L'�K�D���%$�zл�χ��xZea��.�U��KYI��Wc*E�B�1��4"��o��9���78�d���L0����*�����7^�h_*	�aRå���@	S�ke������щ����� "��*��gq1��=���	��{��U,��r��R��gL4���X����˂u*j}�[eJ�z�\R'� �+$�|*��)��g0ZuX% )|����-�=����$ϔX�kj��������j޻�Хa���h]k��bsSٿXi�,�u]�R��\p"��"P��J���nlԆ/��	�_� }k���돽����j�QvO�^�Zu���~��|L(ׯn�f&�-F��gd���=���t�m01/�6��<�^�تD�e���ň"q�9(4���l"�����#��F�Ĉ��h�4Km����9|��*�9ޔc�`0F���`@�!ӱ�|��9ș֯����0��nΈ^�叢��
��\�9�1p	��{�-��n�ߌVH��T���l��9@��8kw�O&>G��79���;�X+R��[��� ��-fL�sę�?[4Y���������鬠��ߝ�h��pEA�Zcj�k��9Fr���ow�KDӥ �+i�4w�zq�}|����l ��0:�&��!����4�I9��W���5"�
B�%��#5?i����o֏�Z�%d,Dz^'�P%���!u�6���}�����쿍�l�g��wQ��L����toc�|���	��#����E�ߧＣv�M�%��������#G�+uPqqlE$?# �'$3�u�e�5��c��Bg�\f�J|l[ᗙ� ���1��9��s�c�_e�R�rD��~�r�L_�"�j$yh"�$x��|)Y�qQ�EM�����k��]Xս~F��Q����.	�o#>��a���5g�D��e�-�Fy�����U^O�C����AkYB��i�)��R�ĺ)���tH�`т�����q*�'��<lsɪ;��b����U����ެ�s�i�s�>� ����5a$GhJʔ����]ιEQ}����F1�I��*߰i.Wq?���?j �(�Yb�5\un�[W@v��J��j�z��9^�F�\��7�qɟj&�;�Bh�ڤ�*��ë���K��n1EE���c��� Ӗ ����twG'#����%Zt�%ܜ�������H�d��o��)/R�_Ѫ*g�&M����6.Aw	Z?������Ź�'폓�T��m{�!���R ��S�e7�՝�B��֋��̵`�IP\	�;A2�D������a�;��hN�lH����N2��j=�/� ��\A�y�0�����<K6���L@wӝ���b9;�^-��|4��w̢3��ѻǐw#�=�w��$�#�e 癢�S]���[Y0<L�?* '靑v���s��Ã�)�$�@R�%S}�K>��UZ�՘��b55�uDoEB�q�ܤ��lM#\rr4���:t.C�/Ėp8 �Æ������u����+)�	>��U��'n`/�sm�XC������ș;�.a�#8Rm����}WZ�|t�!-��)b�����[�&�&���;ڟ�m��r�ń��mۻ��t�Q�۬�\U��Q����CE]Shl��x��u��h�[_r����Ժ�b�s�Ȑ8/]��˺�x>y<	s�LH�~�W����+�㷴ջkm��sb��$�'�!RGLDs�tf�G�Hpt��<��T�J���U����|ڤ{gm�_=*o{�֗3�i(�z����˺�t��۰O,�2�5)�z�(���s��$a���\Ke2��}�m�w�2ކV'��Y't��9{U)�T��u�|��FCCA����֐�,�B��LJ��zǅ�[^��^v�C�c��� Å��6���*��.��O /:R����aA�Y�%�:RC����Ȳ�6����-�Ay\z.3Sx&(��k����X�)����^T-7X-��+��-���&s3EŞh��A�
z�Ƃ��6BŜ��$�=*B�L�֣/�t 	�^���L�WI�⥩����E��۰�K���*��s��z~�˼޺�;r4ۗ_5�1B�m��/�'���x���'2~44�l�ub�x���p�\u��:�u�JQ��$�F���}!�(�1����XXR�@+}�<�?{c�Qg�}���^5�-�����h��Z�����yi������ۚ�e�↎�3Y�x��f�pE�Fz��2��T'�s��^"f{X��lR8`z	IU�sʔ�� �ÍE�����F��o��u�t���]��t���q��*]����A���fV'S��C9<�y�5C4s��'�c�M�͗4��.6�"�`(��#vđ7L��[r9�.�eV:BRD�w
���:T3y|��Y�~�lN)�����U�{Mg���@�W)�� ���R�3od��#~����m��<+R���k�#T�)�V�e��f�!�/��Y`�b~��q�Uk��͘��B�z���hԷ�!Dv�P�M�E*�*<.݂oQ����{�6��3��z��x�����)E�g�Z��<�Elu�h!$,��[�G�S�P��6�u�A���7���~��Q�A���.���Bd�R؟��u&CdUx*+�gy����5�ݓ\���?G�0�e�E�i5B��y�읛��N��?����jQ�P��OU"*V��zs���GZAe7���&C��*[H!<�.@	A���Mֳ
�@���y�߇���|��ƹ`���_�p5��fV���f����L�Uo�3���)�-QX}�[܃A/�^Ŕm݄�9���Ҡ�޸����,A�૪F� �{�Κ���>`�J�,�*s�l9�����R������l��r�_G΄ל`�v�Ç)���v UQEgL
L:�(�
�ı���רoT�.�{���Ԙ��� �S@�w&�{��a#[��Hs�I xF��3x�vA��/��	��1��m/3Ū���~�旅�r��[T�د�PV�2m�
?(&�U+�;���u���??:ڎ\A��Z#����\h�J3 I T�n� ��P�t(մ�%,��m�_r�r��<qw/��l���#}Y�@�SS[Ώ�]�~�����;xeX|m?'���;�>�?��dak���k�C�݀�˷�N_�#X#as�BZ�LW������ݓY�.����UGO]HL38���?�3o=���$Ѧc���o㫕/9GER��?NP����h�iқ�L1���z��Ë� E7� �8mk?�}8'�|f"�Yd�qw��0�����y��W5�I�0�tt��?��+���B��p@�����خ,�P	����%�G����{���t�?��l��|�������PW�� ��p�D�2�g�P��zs�~��㿛+5���VwH�����l�Q6Auhr�s�;����;� ۥ��b�"�'�t����廗sJ��y�@1w�����Ą���D���,CuCŬ8p�U�#3P�R��P �}<�ln����g}dP?������������t~ʸi�4��' ��Q�DE�������C�ｭ��Kr�K���O-���,�y��e]�:-�NXė'Gϵ�ŶlJk�����N\0�ǒ�Z��[Z_�C-��`yq3N�-g5�\�� �>� 4�F+P���O�✟���H���&d~1"�t��J]<�{T>"��w	nS�����7�!2�>��>����zَZ�W�Xf-$�(�z=�J�,Ykb�c?�g�C�H���ᜑm�|t; �+l���\�l�����¢�НJ�_?uon
mBsO��l�.��$'{cA�p�MzV�6ҙ���q$~B3|��E��G��}�P���}�igD��ke�dR�<5g7�ϧ���;n�� vc��Ө���.B	��kw�6$��w�sy$��f�(���$�E�gS�Q�����dP|�&M���R5ң_k *�A���}vҤU�+{r�ST�*��z�C�z5f�\&��p�������D[�Mdjv���&�ɍ�������X����pRE�f2LGX��ONP�תU��D"�@n�E8���U�\rK���I9��~'�
/�|w������+���IXu�#�;FD��F�5�"��7���|��Eo�������e�����6g�0�fkǜlO�2l�q���˜�2AL������jn�Y�c6��b�$��+���|�����yvX(�]W�؊�ץy�⯐�}���5lF(M�%"��W����覕bs7U}b�3��%��Ԣ��<��땇���{ C�6��U�C�s({*˫���u�m��$	ϝ% "_$��Y��{.����hޯM^?�!��)�.�]U�N2��S4��ɟ�}*��8-�ST�b� ��%~�^vq#QBo7$|'W;3���ݤ&R�0ʿ�(�ܮ�Z 3Bm�mybk�?M���e{�fɑ�yR�]����V#eP	�Nx�@�΢��
�J�⬩qQ|[]wG��|�5�mːD�9�����ݫ��� �,�p:�]��E��CD�M~��QF&�[�	hG�e� @�Av!����%
����C=�w��15(#?�O"�����'�t� �	�SZ��Q�����>Fo�63����&�;Kp*����m��-k|W�����@�S������@�ǩ�㑷��G7Y
Z9g��V����e�͔.ȄאuOіo��cO���Y9C���i��.��/e�}�[�`����Ǯ��򂿺�!+��z��x]�=�y��1A��ef�a��
.s�9�&:�]�w�:�d�^��]D�����6i��Hs������/�$Z?�D���&���u���Պ�)�I��C�B{_��u����L��I�	�����R_�u��2(4u�!��2)n	�"�`֫q���fϷ��Cf4q�|}�"Ԏ�Ӫ")�uk.4P��U8�
`W(���'�$qm/Nd�q��s�A@�`}%9�'(�3���CCu��.�_�~���M����x��6���a�+|�uA{�شM���%�W�a�|1ap���I��$�Y�|��d�H��4v?� �tu��g��;v[�K-\��`�g�k���3��,���{��ϰ��4~��tc}��i���3���a^�+#A���E߫�.(��ŧ���ġy.��x�𪓱�����:mC�?����Wf��gÙ��ug)���OE��ʹ�~����ҍ�u�����`!`�,	s�>�C�=a����U#��r�Wd/��>���M��OO��d�形N���q�ߺmf� g
���p��w`�s��j�0yBG��]F�:eOא�K$ؑU�YjϘ`�хL =�3&�8�f搖8�윟۬ףu����,L���G/4{;on,�5�<�5YK%����W��k�E��E�+)A��&��k���6�� �Tc�(|�(����Sp�� ��+��K��´��_$	pQ�H��vu��F42���)�L��-��9ٚA�{^�>�|��Z���(�f(��(c�ke���.	�_��� ��q�@�|n�<_Ǹ,�L�#�5'[�#�*u�AH+\\��~�m�Y%.38�����K�FN�H@�e���U*-�-|L3����e����m��p����}d����A@�Q#aAu�?�=dr�6��V��ؤ�����hg�<+4�m�h�$$��8�C����݂���-����{#X,�i�|FM�V�Y�ă멉�LO����нE�骳7=��4���o�ޛae��&�0��A�L(	�U5�<Dl	i��V-~��ڙ�3Ñ��z�J��DѺG'dk�Mm1���җ�X��<�5}��%^5@1l��?��9`h͏�(�%�O�3��s|�(C���=0��M5���Y�Q����HpC(��9���+����5_�� �{�=�*��}��MC�s�vtA�-��r�g�2O�Ds�d{�����Xփ�_,\�#�ut(e�v
&ڃ�ʨ�`r�DMW�0� u�:�@^~�@/���M�W���K�:`1�b��/	XL��N�7 �EC�P1�S$_X�`!C
�7�{<��*q�t��㤏��m�+W�	�B��Edkz�H;���|�����Q��o�;�b%�������w�a��ʈy�/7�s�/ƐL���_ÚiLvК�-@�({�|��,V������L��Ւbj�Rv��1}�t���-��E�C:�ǟO���$-�"XziB�l��L>�]a�7�#�NJ��Ft�K�����ֆ�/Ѧ0A��_ǯ��S^�1y�س$��N�+y@\1cF3��ş�T'}[���J�H�ٌ7T�i�J�7S��������2.Ԡ'&�֕Q4K��>�x���!������q�������ڌ���D�]�p���6�ݔ���u��[`�_G�JX���*�1[���&9�J8;f�in4|��0Ul^��t��� ~�rd���M���,=�N��v�J�3�%d���d-���� 3B����:҅��I�S�}������	��{fH��d�Έ<qۿ�v��0g7�����w�Y$t�Z���<�'�8��~1��Gx1[/-O�������ڪ�ה���+×�C����k�I�t�0iA�JG����<�:!Ϸ��y9�D�My����0@�Xv$�x{p���ʵ�*�U����P�nC�HC� yLPuf=*>T�j%Hct�:�^V���ѣ�|z�2���O�&`cO���������w!�O}�lC-� ���c���*�e;��c�e�5tYrbs���M�VS6,��u�T�4�,?�G�R��.�:Q�_.Yx$&��zNYѾ�=;p	v��=�1�� `?�zì�Я�����*�O�QZ�Vk�yNەQ���X g�����Ԉ�,��"�b�+���Sx䢶.���ƸHR�Ig:��D9sR���Թ�pZk$C�[���SE�\��.��|�r�%�D�4V�vG��xY,����b���:r���"a,G���D5��6�+QoV�khW��#�T�SJ�e�+QG�x/	�W�V81w#�ȗ*ze#�'�^�VVu�_��;
��o��ux��4rǼ�7"�ڴ�,w�1��_	S�5�;�����#��'��p�q�^o"�<��ɯl�"I��IV0��\ xO<4�3?�d�2E�����8�J�e�^�$��a��b%1A9u��iS^�4e��2^�n���\y"�aX�����lI�h5�<p>�ib��g��Ң�gT�jl����[D�k)�2�
���jp��%��u��lԡ����v��gs��]�:v�1��>]���F0�->�/���cl2
⊋V�H�����:�{�"S�>����a��7E��E1��[P;c��c=���Y�sI.km�����d�gO���:
�\D�C�'�f^^2�BɐmH�O�/\��+��Q� ���K��'Ddp-�������$�q9��՚q�݆���
i6�q�B�bX�#��CyS���� �f5O=p��C��B�*����^��t�ˉJ���,�_��H��������f��L����$��ə�`�Hf��Qk�~WuX��/�#���)L�~�s[�sZ�*$�pw�q!i,J�[������&�.���;���V5Dֶ�>)��T�����l�Kz�a����d��Ͻ#'���<m����� 2opq7��C�1"JOp�9Y&��מZ1���=|+��hѩ4��%�J_�L!_jGMeOT�@���{Ǭ��$�%Q�=��h1�x2�-���F]�;�͋*J�����^�#2�}�So�����Ֆ�c��~G���"�6 Η���ckC���s�{���u�*��3�i�+�`>�7�b��f��u���k�t.f,���	�1��s�e��t�|�9�^M�Ȅ�/_���R��U��:ȵ���W�����̴�{��u-y���m��>��H9��@Ks ���/����%��۔����Y��<LX$���Ӟ�� � ���kvdHكS(Df0T�B�-yE�w����"q�N�:|�OQ@��.^7L���H��D��@q��2|<b�Z:�9Ƌι�4�W� i*?4ED<�iO(�W+�O_��6����B/����>7 0.["�����`�N���7W�%Ғ�&d�����{.7��;�Ć�] ���C�EyN�?�K&�Y�?����:��
�΍�q&6�E��p6N|�b����rR�/��Ǝ�\m�2�_a>�tƒ�r�����>�+>$�����??V�U���ku"����JF|-^Qq,�t7��ͤ	yj�ں/��[)���0�W� ���7��[��+]�w�
R�������1^���~W���y_f�	A��_�f���v;�$�d,d�]�{gΒm�lQl������>L�<_fs�pcX��鴝�ʁ�'񥰨<b��g������~�Yc �DY�v;,�V:���2�e���J|e҄��Q@�,��#7W+wHX��MB?C�z�+;	�F僆!�"�'�(�b���;��֧����d�RH�x[3,��̈�|XY��G����=>���*28�����߰]�~������7���nA=w5�l�xՅ89
)Gʓ�K{�� �͠`BxV��b�SR�����������&`�@@�q00�˭㽡�
�/�U��/�KI/��|�)�*��'4��<���^=�Ns�B�;L�e��2��1��[�Q�|T�$�bN�l��.Z��o	���{L)�"�1.+��yBC�s
�Ҝ�uY��2X���BL�s�@ݸA'v;Ƨ	������)�����_	�3�`�o�TVW���>(�J.��E�9�0Û4v�`
�����&G����T-�k�c���[��`4��'���W;�&��P�*�g=�wK�廡h��8��wPh�g���.��S��j4��c��z{	$�}��T���L"s�bz\�Oc*��ii�`��&��ӯ�і�F'cD+O�Q�4�0;�me_v�";Cu�{أ�t�i����e�� .���i�SKb�^ 
�@��������	�8㻢r�(��?:����v�Tv���m�ŃA��7 ��rM�#$�����cQ��ʍ�F�Y���4W��tfƋωË�t�5v-�t��4���c.0�5;ѷ���3@�I�Y�}U����ƈg� 1M;4�8���S(A2�=��Zdk�q����1`��jLOT@�>��%K�n~h|�K,�t�gT]6���]��A]�l�(l�5�$�����j�}E_���,`g�����cMTX����^�2ŇF\,��{�%���Ty/��6C"�s�`�0S�K���0S(H���ڛ�H3�/?���T��N�� z�~�#T��GՆ됼-�M:��s�gSp1��W~Z�i)3���rV�����{�o�x�ݑ������Uz˧�;1�)��##1!�~�m
c0f��٩��^����R]�O����Ϣ|0}>����~�Oշ�������x	G�.P6)�T���G�DnZΏ�������]�6�*q4v���a�[D� _�D�i��j�K2�v��er��W��f�j��mO'�Kq�0~*SI}�&�|չ�������u��̬!��-AF��m\id�������Q942ި"Z{��W/�f�|rŚF��~�VQ֣;ӄ�ո�د���ʨB*��{�i1�CMMp��t������d�O���{8�B�Q�iA�4�u&6tE����(l>JO�E'�E�����\F��yݹ��;�[so�'c�O����e�=�QSUkCY���H�4/[��`�P�5��XE�S���\?Z Vq5Y��x|� ��RyE*,����D�G����䇗r/RE� �Bag�1$ɱ%���\��aU����פ^���Ǐ���[�$���dWK'�G�����L���BK�x�)|J:0;�E+3�?}�\�)���j:�(���ؚ�\Y'1K�>&gYǣ�9>,&��F9��(� ����ap�)�S �IC�*�/2�۔x�����q+��)4\��DcT���G���]<�~-��5�N������V�h��L�;.�X��^��1���źhT��%�Fx�B�<ABGXxk`��u�c�g�z� %�+gSHfO���A �_
D8�eh3���o����,�0k�|^�?D�"Z�3�:d��6]aX�wԏQq(��O�гȷ�CnK����$U��6�H4s?��3�l�$���0�p���V&h���P����z�q�r�0�:g��^����.�Y{V�J�}A�lR-�~Cl�:#*\p:�v�URJP>���(0��Q':L��u�n�'�#p����H��a�M�ɚh�����F��\3D���%���(�Ş@�������
X��F����o9�?�5aT�VfԈ9�^�"4���������/�e^������/y7 �Y�В!��b"���`U�������G~����ef�LK�КT��9��!��]<e���plN:�z �տ9l��Y�k��:'H���=�n���v�����"n�"CZN������Bv���{�ZK��q)-S8�p&qw)b ��}U��q]��o�VN��qwN�׎��`J��N����?�d�[a@�O�1c��8b˻X�� �i�$�D>�X�@�u�����������EA����/|o�z����$��ܘ��gĹ��VKݖ��]͖�_�)%rDT18���&�o�x�v�?��sf���7?9�+��*��i0X�K�/�O�
����'/�t����P�éVHZ���b�ʔಡP}��z,0�T�3���^Kp�o�7\$�T�+$��J�!�b��q��1�h���8aWS9���6qacVK�^����~]�^_����v�
�(�����eO[�(��������5}����=�Y�WF0MP���C�
��L(��P��t����k��c�܅��k]=����hy�^��:�(��q3#��9�m�RA�N��5� �+�HL�2����i_Je������o��[�=an���W��Q�Ϗ��2�\�<N����~�:]곛i�������aU����.νe��s���O��,�Ί��wC�����/"���}Ja|?���dX�S'�'5��!�qᔿ�Z�nq�9t��P���V��Dx������5�(�F/�Pg �v�{Ti�(¦ras�l�tPߤ�G�~������x���%2������9r��_'�CK�{D5eQ���Jh���+�>UϐN�-��	=�ܤ�C&ڣ�}\�+
�j1c�������emo�M�Y�g_�1�"Y�X�C����n�]�hQ�:m�� 3�Wј�
{�F�¤M��"�l�YH�~i��C�� w���S���C�1�!��v ��\��S�oL"����x�q��J�|W�P{��,�&K�@��]�\v׋��7�� �Z�� ٳo�\�
����!-@��?0��0�E�~�����xnˇ��F�x�.��-��A`�mx":_�������}fƫ�R�ޞ�JU���5�{��'"��kAP;'�sG2и������R���W�G];�����	;K�-#�_�z����Z�ڰ��8}��˱�h�����s��`:�����4b�I���[ʐ��� ��a�j%�n􏠒XG/e����7u���6k�;͝�/��,Q$����ds�tpMq��i���k,;�x��Q� F�R;�C+U��tg����N6�X(��UP}��|�r��uk�I9�����U�C����Yy�-��A1�32e�`=��O�1(�;�$:�5dm�+^�I |'c�f��ue�ئ�,��R�C

䷉���+]׶��]��/���/��qȕ�̕2HI�*��2�fem�`�������m�;�q�\�ګRA?��/��%�����ȹ�2��F�*%s��]�I����	t��pt�G�.���채��#�����D�
)7��Q��W��K$�,�]ԍZ�^O	���r�Ec�Lq�||��b��^�����>d�z%`��v�I�ة���u���ڗ������lC<��2��q{^f}*e��f���/e� ����5����[�
��ć4sQ]�qehLW�k,���8�~?=ͫ�!g%^	�b�S��%��̽Mi'����Z���(���t��%�x���'�r��s&�xͪ(K��h2b��z�q�OG�Bj�xB��KWr��u���y��������`���A�
\�v@�S���}�%U���Y�5C�(�^��z�L����k;YsifՔ�\�L��b�)N6N��#�|�0��_�f�ӈAM�W���b������i��2U��AQ`/GFE}���2�.Ս�!�����}^��z&3L��-���^A����,��N9ZM���#\J~�V�rX��9��5����ͧY�:��
��;��O0ތ��ds'�����9�9k���틱��\���4t� �l�I�KH	-P����Îj`<�×�Iו[�0�:�׊x��q���T��b���4�O��[�9D
A�� �EhȎ1i�:����~� Ԙ����c�=��2���m���.u3q�t�	ߓ|}�D:�$����G���vƨ���������:<��Խ���zօ��.g��������+k�9�o����Æ�Rd}p��t "���E	�g��ei�agy�DG�SIxw���S�.�9��e#�gE`��s� U5��B{`�����^����P���<�&�����N[����:$Þ�ն=H�l�
�|�}�f-��a@va�á��a��RG5����qU�#\�Q竎�sc�f�s\�N}�+�$Z�	$��	w�PJNYb�7�M#�������&N�֙d��o�7>�J�f�����Z���h{�E�	Hq�sU��{�֍��d�y y^M�����F�!?���`�������t�%9"~�<�/��=��/(�O�(�N{HM�$�A9�kƺs#��B"�TU�|^�@m;���,oTU=��)�L��&�L1�F�NDi���I�������?'���(m��v�֙-��D�6�\2hG���f���޷�z�a?�\�%�\<.�T|�q� F�c����U�ƹ�
�j�W��.i��bF#�@/F�E�o��QW�^��WL{Y�D�A� �)��	�z��ӃZ���-r�'�\�i�&�i�m��:V���l7�o��DQ���T7B�-Dx����A�k�&d�h>���J��Ĵ��z��C�ǉ�O�z/���@	�An@��_4:`�tP� �s�p�JE1�v��$2Y�S-�%ZSp4l%���-��x�#CV�og`$�HJf��l��ˇ���C������+o���� �
S!��z�92�:��
�E�*�pd�.x%nre7Dʴ�b;[��=J
��.E��.�5v_�b ��0,��߇\�qBie��BM�&�B_}ٳc�8G�G"�l�,�����G�(��"����<��,'٥x�U����H��Y ���Ю���C�{�����uH�v2��� �0r1v:1G7�ER�֌	�L���z�7�ߌ
��Ji[�%�b��\3L֞���˒ݧly��8e�زN�0�_��,o�S��]�4�,�	9��D���8��]���T����}�h��
3�}H��������_�Y���,y�2O�5_���2��F��~����I���F���??��_|�P%��Ǳj�[+ޢg�}G�>PȕU͒i�!o�PF����[���2��Z�3I~zKφ�H���9���$�:����W���L��� Ö����^�L+���q���y6��
6�G�NR;���tB�b��ˉ©JI&�+�|
-c,�7�'�~��z�q��	�6z��Ä8�Y�n�=�H��f 8]�9),�ڼy_�gl tP�@k}y�@{��r�[�!��Uι|q�w� ��]�4{�&~rB�QL�'���98'z��|��e;���;����y�)d�@M��4WJ8���[�_2(3�$�\e�IW��/�0�I(�𔜶z׵Q�ѐh{!���p��{p8������5)�ww�Rte��:/�7ڹifut��"�3� ��=tL�ٲ�RX�G��'�{#U*�0סj���ו�45Ń����}������9���(��H �]!)v���o�r�n�K�(�r(:�N@�g��&Չ@�u�?i�8{`��I!;�Ր�b��a�C1�_���ĺ�������>����5�ƴKpl�Y-��/f��=9�u��}W�U��!���d���d�R��`����&^��1�O�&��񷑮�b�kFVA{�"��4��}EiB�*o"���\�99�-�h_�����'��@�?�+�v>_�"Id�eM���lG@�τm�M�t��^Ƶ��v�Ƀ����?sb7���������E#�i��:?�g� ,9-A����}�L"5�������^�d��L�!4~�u��k�Dլ�EDl�資��\(���R�� F cJ���oNo����i�gh�>#�]�,9�{9�o:�f4W��W�.5�<��U���B��2�aG���B	fƵ�,��0����i���7������u69�7�J�� ����o?�.ǂx��x'�J ͫw�?�~��Hf��r��;3Ek��k� �b��]LM�VG�%��2U��*։W&Sc�w�*�ʒ�g#��	:�c���-�g�.2-1a�ڑ]�tXtK�Jh[���*�A�*��^�A5� �ސ�X�l{9��5�!}Q�:H]�9h+����F��Fu�Y(;}Itrt��03�T��9��Ml��c���E7�n�e&W �I߅=�آ��V�� l�I���_&��Hǈ[��=g�LPXk�q�d.�(m�M[������*��
!)��"*s�`����gc���fpP�N-��iaY�m>i�]��z���+Ao��%R��~2���FVY�Íٮ����wX3���a��{R�W.�$�;��:~������~�?���F����nf�� 3�>��R��Qa�1޲�_�Z��{�D���Ae�٤#�z�l�`����"E��E(���i���<tr�"D[���d�Q�����$!�Ԭb;�@��C"Խ4�Ԫ'9V�n�º��Z��v4��f�~�?E��;~,�����4'��_�B����-�ȗ��V"6�����m�dS�F���?Q%:�"�ܺ�ژc�9��*�|� ��Á�������'^�(-P����.찯y��K� ����$�=]�����Q��x �xC���J��p�����㖆p�]�4jWw��5>אXX^�vd	�� ��PۭI}�'��`��xr\�B-�W�1�m��� ǾN3Zq&<S����^�Lx����yȸ]9<�W�?\�a��*r@�(�O ���&�8��fO!�׈6�������q�Cv]��x�� ��+�����@��L�)�s9K'{1��O�\/ꠀ�����u7V枊IR��h���v�M9��*��^tؒ~^n缸��M��`!�>��ы�$�3��}��i�*��>n���������j����&��,�P�a?��]����_*lpM[.H*�!PH�b�����|��WVn2%�5���\}R��q��/����v]��&F�6ӥSB�V�@Ъ{�r �ﯙN���W%��s��&p��b������c�{!�|���N��Jɨ�WQ�+1��`�kCFh8�O���LT�D��'���+Ui��72�j�\?���%^#']�JwT��D�	�Wo�{:�"����HI����y���D��Tja��/�D[q_�~N����8�H0#����A�2��9d����孊��Y�W0�����b���,�%����;��ղ�2K�EHL�Bx�B�bZلk:hBZ���	�ݝ�ڐ��;0��<�����-��I�ځ�C��;��YM�s<l�Q�Ņ�hV����]��`V�?|͐:����9����Q�S8��P��;�TQ��H���IpQs���C��X�_��q�^�}L"��E.]�[�hG$�~�³��{őn�;N�h�� ���x�����a���Xz�ơj���p��@�)/�EJ������K�m)r��x����$�z8SVDV���V^)e��B��h����y�6��ݞ1+[�u0	� �f+�F��=m�u���R�Ҽt|�RE�RS)��9(\P}ռ����G��t�(jIGƾ58�3���#�l�Z�KY��ɽ�~>AS���;�ް�\^;4�ϗ�k��8��$K��.��g������")K��Og�Dw���G��� bmf�'���@�B-<�3q=���7��£8RC���k��tM�4���A�f�ȄA�	]݃Ե� �����En���Dt	�el8�=w�����c�=��Q6�� %���dj��d�^�߂a��ű��og�k�OR9QI*>h�炞U5O�U��`�X��A��5�5��3<���������*�ۑ%���L�؂�OPK�T%�*T���P���1C�sC�v�ҩ�@�bo0�؄\��38N�B��Mp� �K��L_��Uv�_���G��!�Ш#gҬη�Ծ��cwMQ]��i�.�V�O+�����U�R0\
���C�~	���/���J�k��N����V����R{���KɎD-�!3��xi3�B���Ϋ��mMp�n"�(*�G	�D"�`�vG����%.�
-���Hp���W�\q� �j����ə4�����U��İ��f��=4��9(��Ԝ3�ʕ{���$4X��ל׬t_�~���� ���X�t`p ��s�Ѽ����{%���!��`��uVˍ����w�U�D� �^����R-��C��c�e?q�C�@S� B�9D�����&������y��
vTUI�^�����d[c�|
�ԞA�=s������k�7Ѱ_�t	@{�ApՈÞ^���(�R|�Ǎ,Q���}uF#܆���J�wF9��T�$FjV!��룓p�[�,�c��aJ����s'¹��nd�Џ�9�����I�4)>l��͋�+���w�r�K�ܙ�q��`�^��6��(D��p֐{Nr�w���1�T�2�$l���r�z��;����kU����BPpZW`MϨV�4�(�$M�D7E���!1 W3���=��D����c�ALP�cR�@��@���,���m7�-�x�IZs4��%�g�[#��W�K�9;ɣCM�AP� B��~!/\�,0�?XB�9 �k8Ɉߣ��Z�fIL���>���!�0�F�ƝA�%|��ff׽s���&���m�U�2�׆2�¼ǻ���0)�Ԃ�{����3~-���k�뱘���V�ĺ�a��\Hw��Q`�#��.t�;�	R�]���ovzZ{强;Z��c�w��>*&�?O�gSyj�����$��Ƥ&�V�j��u�C�a��L��t7S����&q<OKJob���xBb�`�������I-b����:t4�Jz��2�١���)��RV
���v��F�qL�c~�b�_��a�J��1M�.eZߑxi2����Ah��{��	[����j��Ŭ����V4V9�K�]Sn���(�\��a�sh?�b<�W�-"R���o��ķ��Y¼��+`�[�y�!,i��l���dq��O냫�/���кNV7�+͌�LB���y�t��z+���8������-����ֲ�)U���/���̀�3	%�N��9���
2ȶ6,33a�B�0�wEBm�;�t�=��~�m�=�M0�asn|�q
�lS  �	�&+b�vO�_����:�>�����4�3�%�6���I5��l�Ï����v��t�?�|��B}��:Ǯ*�k)EY^@�U���2qa�/(�NVr9ѦV8SF�n�L��`�Af�z�$����O��a��Dfl?X��yv��j�n���e���;���6� e�hf �,��p�Qr\��r�^��ӗ�yJ�"F-�Y9���w����s�cu^5D���X
�0:s�u���5�Ǹ���\S�6��+/�l-����ġ,s�p�k⁛'����%�,�l�G�~��c�����
mX^��F:E�ݼ���i�Kǁ�`OP\�|l*�m8H���dv����s{V<�ږ��UC�!D��xt�����Sz8E����K�N੭T �K'�-�7*Q����ճk�j�h�<f�r�����v?{Y�Ey��O֑h�Xs{��X���L����s��(Gf�=AkW��}��Sy�� ����^�M��I�.�{�{yt����A��}Z�Dw@*zJ�#�j�ЦU)z�)X���P�L��(:_,�,L$X���$Ԝ�������h,�ԑ�;�ؽbR��XX�T��$��:��9�����G���3-�Ċ���{��u?5�2�ĵD�9Q 0��(s$���\D��)�B�7�� >f+9ywxՇ;�_��(���T�x���M�U;L�a�Y/zr}
��)�c���7̪(�a��#Kkۇ׈ƪQ{%��Ro�����UtR
�4eO�GX�M1�|v�FY3�!�y_/F�aϱ����7�\���q� �s���p���<�h�z�'iO����l�F��A2j�hn"���?���.���hZ����*���� o�Q�$u�{���7�u�#�i4o�N�yq�N��M�U	s@LQշ���� p� �巋2�F��7b�&�'{���BĄ9(� ���)�%���]���h����m���(H�I�d���C�'#�a�1@!�Pǿ3����^@g(�X�D<� ~H�l[��,j�V.�p4���ā��?�I��Ix���5� yE�θ l�P	 ��Ͼ��	*��H�.��M�9���⺪���Xbk�Z��&�|�KFS�M4Y�9�䖹Ĝ+,����qx}q"��ˆ+��/�		���Q�����q�����$�'�W�x��?8
w1G�E�o���z�)u����-ո�H�VL���HA�&��j"Q��T����2�G�t䮓�K�h�G|c	�JRtk��1`��/9�9���9����&���������D��3�o>0q%��5���=S[�c>�2*��a��D�=�m*�Rc|;��o�P7 7�Jj�fgNANA��������(H]�t��#Z���IX���H(�˅\��7� !��J�^��پ�5C�UƯ&u��G��-�)�RP
]�� �b�W����!#�/��ͦ�`�5�ʇwp�)a�ϱ��t�jN��N<�
�������
N񪐊��L�׉P����E�7�G�v˧~�՚�T�⇜��l��.��[�/�����Q�\�?���	>������-���4p��7������`ׇ������[�ӪWx|4F��o��;/>8��5�}v�qj\xԇVˑ�L���Ȱm-6�i���2H"O2��K��0#<�F���:,�N�(�j��1)D���ϯg�g5(��gkX�M�?Ja&�d:���9���k^���]�����u^ߓ�ާM�?l����7~ǌ|�	肏m2�̵\_�Y����c"k#��4���cU%d��0ꎴ��G��a��ֆ�(L��8�67�-�%��Mda��G$-�!Q�5�_ն����Y��~����/�3:��x���m�[I��*�S��=�sX�Y��+�fE��bYW�H��繫z���:�sx�m��C�N�\�왧�����I�u�K$YD��� �0���r�F�&O�p��ߩ[���i�����㔖O�����"h��JTX䬶tEg U���~nx m*� "z�N1˧���([`�V^���"�"m���޹4Y
'��L�VZU⹦4�u:O.��B�Ŏ &g� К'N��j�-�YK�O6r{�7mA:>1I�b/�VfFBV���h��G�4��L�$���/�]�#�å���	I=�8Q�'?� "��X�
�n���W�j���K�y/g3Cn�����RYFטB�g��>@"�>��SY�>������!SJ���?g pƔn�Z�q�5^��9�����:������BT�����������Ι2	��贯�)��qͯ��cH�06T�S�(�ǻ���/i��r�U�H�Ux��]�A���68��6��~U��iR*��C5F_�7Ѥǀ�{��v�\�;�7���,��?B�S3Q`T�O5k�Ʒ�A����$���}�����O��uݯe�w��9`���D�'����L�{ ��	����n��>���yL6�+P��t�������C��AW�.��-��H��^㪛�s�x�;}M��{������7�vM�uV{����������nV��.���C�g�S�!R7c֧���g�lc��/!^~� {�l!vi��,+�D���%�<���)�/�D��l�mU� m�fQ���/+��~�a��f���q�\��4ךɌ���'����vX���@E�Tѻ��O�R�S]ɦO$�hYYY�89(�3{+	��F���W30��_"9rm��-�z/k�9���WJ�����t� ?�ؚ5�|m6t�3>�
�ͱ�B���.:����|�3���᩟��x������C��Xc-2Ԣ����Ɍ?sY��I�}�#��,׬g=Ew����a��gSnhopZS �Sni�&0^�^CIJU�u��Z�0P˟է����L���sYE��K(g*��إ�(�W]ݜ��"&���k)e���`�q��a���D��&!�N=�w���s��'vW��h�9 ,:J�5�l�X�P���9�����O�_�K3�y��F����P�M",a}6\�Te��L�<��xD��a��f�z,g��3fI ��P�Kg��FW.�+V�)��{���BNT������պu9�ҩ9җu�JY�q��꣫��K]�W� �:r�8�ִZ6���G0�� ��ӊ&
�r.��y+���l�o�A..ޫ裤u���g���5�jH���[�t���=Y�� tzo vW^���w�8���"�⋷֣�$����w��6�b�s��X����_N`<^׉M������U
�PM�8:��B��nA27��0)H��]pƕ`��~���6��*�Z=�?���8~] ����VV,G7��#�1�R/�,�lC�qs��5��5_�e���b}\���At���'�A�� 2�Ʀ�vK�P�H�@���.���)#�k`jI�ȵ���$��̫���o�s)�"D��괱n��X���<�ޯ�=������u�1����Lx�	���~���)�̑��¾�=Z$!uf���ХE��{-W�U�Ή*���1p~-S�{
�P�B��m�g�b�{��n����D����W��K���;*�aP0"�!��jd!�S�y��
Tl)�M	;!@��i�T$�w��W����ͥ�r�x��O%��l+�]x��Z���zz�&!��[���t���,	04MT���]����j%���М�t�/�^#���"Яޯ=QVkX���'�G�R�&m'β�"�;4�ĜR�q�Gz6� �g��j�D?�E
&�}�gpz�IR����f< l���<<b)�\�yDB�Ie�v�^a�=v�0�l��T�[��}�s����{@�/�(J�E�׃~k��`U)�i�k�l�|��XU��Jo,F�^���6�WS�� �n���د�k�<	vt���"�`��y�ك�H��@�� �G���q�ÀzF��F�{�X�}X�u��׮PMs�VV�`���\)&M/�/�:�r��[*7��F~=����r(��=�AJxe\�|)n��.�C�V�]����6����_���7)0���\o��� )�~~�m���j9�q�ʰvNqEh���j���B'�㪈���5h���C[��ry:�7M��ԑoi����j�g���=�i�����_�x�ј���ʼ�(a|��F��n�g��1^�-�C4eޖ�#�\\�/�J�����&�TF	%)�u�������{ 8n`+��7��>L�-|��~���)`�J��-7a�Z��u��%��v{��о1�����.L�&M��D;䔕�rr�=ˋ���3�,Ёz�36��4��ک��E]���Տ���W=����(Ԙ�p`�C�:$�v@8��)*�����21 ���_�J��c�:u�����=���&�-�2�~��P��C!%���0��P.E�*�p�"C���[T1���x�Y�c�&G])(e���*���.�� EiN�e�ֺ	�4cJꙫ����3��<���Q��i���3�?��?0~������S�f7��U#B�!�.���f��� !�Zۣ����Y�i#�R���^C�︡����o!���x�hrw'�c�3du���N_Â����;Т�塴PP	5*�aI�^D:#�ʭ����^���"���	Ea!ܗ�O�ɳJNI�5 V{d��8�5����I�"l�c�\j�������Yr/�ޤ���^���v� 1�R�V�����0�|X!��c�c�J�+~?��EBA��#w��C��8�Yٸ$eBz�� ��Yc��%C ���W#&ׅ$%`
ڝbA8��ků����C�u����Yy:�P��[���T���|�I�N�2�#Gi��"f)\HJ\�x����զ,WSo�l������R�\"���qC�_ �;�X�%Q4o�f��{J��|!.K�kc8&l�Q�'����:VX�~�Y�ɵ 5����xQ@Ɖ�+�(v�Xv�_K��J�Xɍ>�GiO����S���j^����#?��R�#���P%-�W	r��W
�'����T۾��yЯ��Cr��\o�.�2=��Ht��b!�1�QZ-h��]>�&��I��r0nRA9~��K�΁��-0��_AvKl���w�b�}l��6�NXi�x���o��r�%#���1�QK5[��8vU�|��Jq�%�P!yS�q]�j_��]�Jw?ʨ�pC��
�����m������
NU@5�=����$j�lS�^8�>"uk�,� ���T�3�xKa�r\>��Ÿ���qD!"|�~��D�ƕ���|*J���-n!����	g�8«w.k!�Z`�>K|�����j|cs�1�oq���U'#�-FOq;2�ƃ蹫�xL@�JF
��?��_����YO_�����w�]u[�#��e��'gѣ���A�x45h�D�(�Sp]���8�2��R6Q%����7��i.�~ñf�d��1����!���T�B�
F��S�ɴ/�� ���� ���0��A�<��g)��k�b�����j�)�@룓g�XY2���bB��E�5�ȕ^]��w]�����ZI�I9�~$ϒ7��(E�jǐ� �|?������W�+��2ȝ=1��J~H �g�^O8Ťkw��o��1�v�8��oOQ�
.͵�A�i�w��.ս�0i��	����<�Æ���uro�߫噝Y.�ň�\�{�3P)gh����+�5�� ����,MX�;-�u>�y�3� �"�clEK/b�v�E��P4�$�4��>D�sL�6�	9��*ױ��u�e`-Ƃ�im���d�Fh\o����f�U�{b�a>��F���`���o:�D�UG �p�b˶�V�YR²k<8��a>�H�+x��嬀�S�ZL��'�R)`Yt���ά$����1�q��� ���(f�f��I�pOa:���\]x��y�ed��;��׮�pq8V�r�Ǆ`7-������3iV�j�Lvs�f�"��$���l�&�_�-�W���:M��4���e�-W��lO>�=V�VJ'�W�Zu��'���^1�{=��X�]QT֝�z6qdF`@{�%���y�5�Kc��Ha���7����ѹ�����Љm!`�R����ofY��޼�W�Ԅ���[D	{Cg8�B��6T���m!���f���\;/SU�ro	�NpQ��^A�쥐�o-���-������^�e���)3��՘��@Z�ۓ�.,?�?���t�j���0��<�%�h�0�䔷D��,vt���A l��ȱbXk�RR�L[�_�
~۝���8T��[�Kj���:����	Nɍ� *y�M��bdj����ut	��C������;q^~tlw���~b����!$,�� 9C]����dڍ�B���P�܇-���o�t��:�5����.�b�C�6V+w���U=����_��3�^MQ�M��k:E��_��{MY��tjLh�tN#i��V����$���w��b�Yv���Є!�T�A��,�~���.�����ϡ�s`����d1�Z P�u�{��!e'�j�$v�%���H��N8�z��s)B�y�v��#����jW2��t����ȓY*��wpd���!a�)ϻ��}�g�J�h�B����<e�Nx4���؂8����#�/)@e
��6�gl:m!����-TP!��~�^S�:�1�1�Ҍ˼�Ar�$W����F�3�ȏ=p�镼֭�������My�,��A�gd��T٫=�Q�$fb�gE.&Q�87���4df��v5��iB0[Vt�r���,���aA{"�E�a��E�:�Z���
��M%Q�a3ؒf�S���7-B��`D�;�ʦ�"[��ꦱ�&�>hv�8�6��D{,���
���N���+���I����5�s�Z� 7K�K {�t���Y��G&�d��ϲ�����7v�r{�8Ӏm��l�"��s�� ���v���q�h:W4VB�]�̐h4s�Sq0'͊�TŠÝ���m��ߴ�!d�5 $�����w6��BQ�`�S�JC0�� ,Q;ߛ N��hVw_>QpK^��j���2�Г�j���ݲ�����諑)�|ݹ���|�y��GBMY%�`'� F��[	�Wo�f[��wnϧ`�o8�>�=���3=��5Z"�P,s(�I�ϖ=����QBNj�{
B� U� x?���_�W�D��:����2����3����u���� },�:��G �dG�*���B�L���1t�I{K&|^*�9b�W���oS�t�+M��kqbJ�ʢ t��ȿ�E����FV!;*������..�W��הE:��؂�M{�H�4�[!�F���$�+C��n�{$�H�D�֦��w��;��];�9�{%ö�S&�M��i�_��+Oa̅X����hdFFv*N(OA.&k�({#�c���B�$7��<u��HԴG[Q �����ؽ��CE��'_߆�����Ʈ��Ed n7C%$F�t��C�iKf�X�}�`(q�D�<~�⛃������K-�/x-�d2��&�{�j��X+��G!|k�Q���p�1k�l�YJ��A�J�q��g�-7��V}�<YU0y���Ǟ�A�0��a��+"{k��+���:�a��e8��WJgn,=Hf����J���ד4���6 ���.����w8���d˯���0K�tE����F����L
���z��_�P3]�e�e�#�hb��,l�==N�7��W�0E������-�5�f8��i�P.E���Dٵ��'w���i�G�h8�o��6�q����b B=�`hQ�*�n���?�����ʃ�?*|���T{rè���V0���=F���:7ו7���G�
�7�ed���U�^��v3�C����T��lD$�()=���pE4G�K|䉼��_�M�Ž8�սg*Z�\k�ܰN�(�^\�f*�}�@!�m�)���)p@j"�[�>�@ߘpi
��'����yHfqE�Վ��}	(�啇e�uvv(�	�����P�ɒ��xՖ�$}-H5!)�{�#�.�w�8l}���J��|���a|�>][����9
�8�Xs��y:T�9Λ���$�!��F�~�,�xF���|۹��/L"��>|ܬ��6rψ��x�4�⪉6���aZ�t\�<:I[�`[�d��� �9��C���LD��3��+�0j%�%H���j������R����e$0 ����%$�$�������8�M�@���RA<���Hy���>��	�'�r.�N�}�Ia����[l�~+wy��6/��)��*>v]�w�h�+��S�/6p��mV)	��x��ܻx�p�-��^���
�����7Ε2�+iҰ'�xTPY���e��ZA'��;������2����Z�;�dT�|��V1�#�@�20�"�yK\��QR�9==�l�:�!����UsL����zꦞh��"��Y���2��rE}�����"��G��lU`�/@��+ȋ�z<$���2//sba��)-D���AeR��I|���h8�RS�:^�,�@�_�՝Y�v� �Ӯ��8
lQh���3T�wn���gG%���v�{�����њ�_L�h����:����^b�l@B�b��>k���O�;9e4r�y�\��E�UkP}�_LP5��gG�1}A���GJ��r�O�nC��@�:�!����D)�lS`ܷ6�I�m�kӭ�h�aAK��7������2A��*�o9��j�\|M~Y-앷�f���h*���S��� ���9�g$��Sw�Y�*#��C/�*?�6��(\ vvYR�*�en�e�dm���MgZ\��3�}]]�l�y{љ�����O����_@f�v0�ٕ�������VO���r��S-�Rzr��~+��PGx+�ס]�<a��k�kozuvu,�K�Sc�G�y������
��V���ኗ��X������[FX��?g�݋�yk���_3�8Az��g�����U�� [<��:)���Pg�v(q�)��e�I.'��܆U���+(���q���Ն}���ɺ�	p#=Wϒs����B�mĺ�%�ah_���`㸐�#�e<�\$(Mi��:%+# 	ͱ.�KH,�+[��v4�ڄ����Cwz��`rKݱ
L�]C<��7��ʼ�3��x�?a
1�F��4S�ݓ&�w�/9(�L��ۺ	��ҬKy�����r��BZ�D�Ж|����a�=����a���	��~�1��7x����P���w�������\U���/��v|H��Y@(�XS�O`���`asݫB���EU|>�s6|�IDiM�ch ^pJ��M	�lo�[�ˋ�(�?�U���v��HFf��f=��GN���fB�[����5�O�+Q�+U��.W�L�h=��ۘ|;�=�} ���v�W��,l$�:�o|&���&\rC����+$�ۡ�c�z�>Cf�䥓�����P9��_�8����1���Qz�K2��w��v6T$����o�'jO㇠_~�����f<�ukˮ�b�aY*PF��-vP����1C���)89���;�*�3]E�.�u��댘x�����)8R14[m<�.Ԁ?�$ř8]b0)xK���\dC�4/�:�M��֮�7�?⊦㊡�;o^L�_�\���t� ��q�_;���[���r4�>O��!g7�1.Y��)��D�7~�\������(�0'��?sBgH �<^�2�d�����v@F�;a���|Twi~.�Z<zk@
q6�ܨk������!����N��e*L�z��ѩD���mԷ�P<
���^�~���(��n�R�����n�3G[�[I4���e;|�Fۮ�:M���������\X� ��q}9^��گҷ�OId�6<b<�i�O�<�%��"��EL��LR�=ݭA�ݦ������\p�3��y�}�R.�9ˏ���Q;���o���B�'[���l�.�s�^ə�W�6��@�6]�&���O��/l���u;�Vh�r�'�f�w13��������C�?^QY��C�H�uC��o�S�6Ep@��2!��8���d�y��r�aNOCYw��Qj�8� �X�T�.e��
F�{\�O��
��j���KKAUl%n�Vbm�����A �,��#h#��/w�L�5
��VT����K.�<-�2{	�5À�-8Φ�0R��t���c�㵉97E���/��Bz��X{��U^D�dt��]�|�������˻���l�)��F��>�A�Ƹ&3�Mm^B��-$��L�]�B4���8CVqђr	�u�Ї&-H��4�eb#�8X����Y���B��1G ��h�q�>��r�Q���`�8]���K۳uK/�ua�p���|�WK��M�u�>]������7Qs:�]�Qј�Ep��d�.�>�i�^��o��Hz�P�%dun$c
�Am�8/�h���C�y�=����A����\��e�7\{[N�˓��8Z�MW�l�,_C����G���������$j7��p"��׹G��_��c���[��Y� �hrM|zt��H�)d���r�%`1\�I�%u�;��2�ךG�u��K�G��R�́�c�� )eGKc��@�^��_,��%L�R�s~s�C���v+�W��/3�Zs�o�I��R�-{���ޣ�	�I�	�aX�]�B���lJ�Z��~fF��i��Z��i~���f��=`
fo_�ij\����z*�h9�Y�>�E�����8{_U��E�{q3\�
�VH��"W�0��IK;�a#�iJ\ُ_s �T�߿����Ꜵ���}3���� ��#��cE� %y��+5�i�}��F��_��tvڲS�[z>�#x;�:d�j˳��8���c�����ݾ�)��i.����K3�����nw�6V[pG�,��n�V��༿p	���!�_�U[�JN�� �I���S��#-��gS�l�c:�?���I�5_I�}!��J����|�4A8��j�R���������i���"֊��zk���K0�&�Vr�'T��=���ʐ&k�8����Rkz� �2�v�=�ѭ&P�&	�K$�@�����5�:���9s�C6���<�G��9���nSq�ez��5��H3�.��H��]�i(�t7y��}��$�K��V见����W��7��h��òu�������p9��z�$Sc�2Ô��h�� �z�zHN��	�k%&�����Xb���A����jJf�Uk����6mi�>��µ�2	��fE�֥����Q�b�^����uh@m��טth�ڸ�Vs:�`&lwsu�jq�U��k�v���g�q�:ޒ�����C��`ӎ�k6��$�T0�͙:�<���=��H:��Ŗ�'	����ۀa]=��W:hzt�V�Y�'����f�B�x��k����YuQ0S?���F?2h�E��2���C�����*R\C���%11����3�&3�� �~���5i�� *�3�mF#�+ԤY8��:����m�+�VUhd����ٿ�^�𗨷`¸m�=@u�ۮ<�FI��Ǣ���R ���Pm�|��5M�KG-�Ǔ�go!7x�xl闫t���I&�(6m��� ��ʮ籠��W���[�l����-�չ�$h�+K�K���R����ħ���"'&�,��GkK7��׮y���r(v9x�/�_j;�)�Q�0����lZ�j!�'l�6##�@&�_^�z�+�'���;�z����1�����g��ﱨ����qQG����fG'���L�Dӂ�"�!��|�v�?��)�`z��Fx�(���#T[�f�&��6�A��XT��1�ˣ݋�њOˍU��ٹTq�:�5�%+�c��*T<����cU�"��C:���e�%�3Z_��}�b�j���[�9��"-Ԓ�øu�O�>Կs��yr�����)[�x}�<���A-Z6]��V�|TJ���c�D�(�"N�bṾ�1t��{����ʁS�-	Gy��MsZ���Ŀ%#���B�h��&���]�X��*�u��G`_Sc��]��K��.[�ӋØ(���3�X��3*�|
g�>5�����R�7���S���6
{��o颲��m�}��͒�eUw��>���D_�ڮ�ͼ�_Z���t���rs�z��Z�*uZ�p��ɰ��F?�9�Sz��&f����~`��Hj��(�[�2T�
md�L�<�Q�}��3�k�&*�7����s�T���݅d	�|�g>K�YQF]�M�3��+r9�I����KN��^�A5��L�d��%�{n��.1=���$������N=�AJ�9]�EG��;l�)�sq��� c��W���e��"KLC�jN�D�e�K��x��@���\@�uX���X1�U�.�V�Cb�B-�ذt�PS�X"(qcʹ�N��h�4���� b���ϣ4x8]�Tyi�MV��~��)�vC�Wx�W�0�U�S��TAE��9�;n7����{Ӛ6`�B���.���!�އR�P���ې�)m�q�Goܑ~�Ujd���e�"�4%����6/9O�.ٞ�w�Ɍnw7x�j����A��H�ꡂt��+ �h���AJPu���aѾzПH;�2�j�#z��J�� ��^�}E�{�% �����h���?��%W>:���l�}�Sc����::THhm�O=T�'�jB@���ϡ��	g;�r�ōV�`yN���v�|c��>�� �,H.Im���݂���[�f'�J�ڊ���-���yszT~籦� �J+��1fj֊�[�mwl��qH��>�B �!z#����u�5m�o�����|#���̱N�T]�u��n���ʧ*�c��7q}�JYI����'�ӑ�N�Oc2��K��QNHR.\�e�J�M�uMk)�2D3Q�[���VAq��D��ф�F���hA/��m�Q���fw�"vUmm�
j]B��)�2{N�^_�s��$���?�h~l����뱒ZU�KoWT�躽(�
��fӯȐ�b�� �Q�b�v�R��WI�>縮w��*��Pl�&YEg����>�Xﶢ��x �h�:��;���9��QF���!��5��S���W���b�#�l�v��B���?s�<�/Ĺ����ZA�i��^$��2%�hm��3������
�,��z��\SH���m�E�'���/Ш	h�}�����
V�;L&E��rUg��K�d��n��0b���s�k�?�����I�`[�t?=�����,��L���������ع�٤2j��X��N�U"|��i3)���5�J�PKn}&�Giƒz;Q�7�88<b���i,HO�\�4�U�֐Ao}M�| Y������0m}ZR���Z��:2S�ߡnj`O��cf��X�J������]�u�3� �$�Wa����=
���7�G���n��B��,N�G=��0S�3���6P��|����z�ɠ�{�K	����W���C�"��˔#����9����$F��X���Q)�Iyf߰�wK��9E�<:��({��i�KoO���Z�w���t΋T��wQ��Ї��3+`Sߨ���i3��0XtB�BJ$so�%1�B꾤��Z2�Ȅ]��"rҡÅ��Ӛ�˜��"��O�[wTT�����*�;& *p��1&L�q՟w-[A������,��Ax�V��(��܊D�6�Cy�Ki�gܹG ֮��h"+��
�$�Ȏe�Q@P=�$������!�ڍr��؍��F��"�̉��ۮǂ��{ip��K�5"�/�X����N�8O��MP%���o�.�K���������e�~j�XJX��:(!!P�=�%4Yn518��n#�8a�c���8x�:E��}�dB�,�#y�c�אp�>�r2���{�hLy�V�4�L-d��p��Aߢ��Bҵ7Wl�]�v����­��M�������i	"_;�@�K������m��7VU��3E��x�L:���kL$��U��i/Nl��(�Ig����Q��
d��cQT#��o�����9��H=�1�t_���{�p����� ��4�윜�>v�^U��	����Q7�|��:3�E�43i�8c��c�8ӣK̥�(</?7��F/����[����\Y<���X&sf7��'�(��f��b�0���pV�V��л*j�"����!��+>�k�%u��� h*�b<��R�Z�ŀJ���m��"إ��`�r����"D�3N��E��9ឌ���!��})A��k����5��D��x����.����6���
T�!�$*�֡�^<*��tyS��D��1�I2XFݯL~�{�r������RD?���5��ZI��0���H 2�����@��(�zwi3O	�kBXA����%7)���X���t8AM��;��A��E!�f�e:�D�}5Ʈi���2�7� Yw�GQ�5(��	T,j�����>����F˳ ���~�2��!e�t��q�g��20�Ъ3��_�奬`"<K8��c=˫9����U�{V�8wq��EJa@���q�v���hPf�ڌ�����C��p���8�v���^�| �
���$r9�c�}� �&>�����$�=:��c@j�-q'��`�ܼ�ƿ��!�Ϩ�3��2�
^���oSa�:"�]�%(#�Z=���L�(�c�F1��K���2�Kp�����m�1���G|l}�w,4Âґ
?�ݘ�7��k�7����dR?�~L�.ĈY�)dT���H~K��pT\V���շ7�m׭O����6��A�N>/�+&��tFp¾�b,d~d�&ƍ�X�ʙ0K=��n?�X
K�14���#�� �[w�A�0E�v����sh�Mn#N��P�Ԧư��H���B�*�J40%t �Z~���Z�!��gn�>pT�9�����8��~�}�:�l����h=o,����4��d�YAM��>l�o
fؘ��0�>+-ݸ���>-Ã<n����FIK��޿�LXw�\�������QʁH9��\���n0/3�Z�3_��KaX�������o�`��_�[0-E4�?
�ʑ��5yw.H����f[n�or�?�WtW�wڇ΋O���N�Z��v~4�	%����)��?��tPv��`����/X�	o���Ά-�)A�Դ\|��!���v��V��t�q��5���"jD�rX�Y�h���R�|=�f҂���ƊYOD#KY��'J���9
�q�����l���+������M�^Xh��ST_��*��I��Mtj��=��T�Lu['�Z����,梃�C��x?I�7�jӋ�r�������Ua�;P5���}�P��3|������AJ ]�2:bU;�-q�v�������-*s<���k�q�U�|ȼίp�w�5v��,��,9��"T���B�W�,_��E�D�.�E��F�֘�؈��R���/��2T4��Oj{���?Z���@9�q���8qpm|��H�af��Լe�f47dAu�b���Rߛ�Y��Y�b�N� ��C3<�����u;"HM��"|�C��3�)C��@-^r��/[�O��<����8��5�e�� h^�Ӄ��"�s�ߗ�Lze����"^{�;]�~DU��������A�E!N%�E�R��Bj"�c����{�꾊��t����Q)0UBX5��dȯM0 ;1������/W�����O�����q�����Ĥ�'�چ����D�T��}N�I�'�^��2C����8��+^F� �u6�􎯮���l̋
%]CΈ(`���[q��7��Rk�c(�s��X�*�6��\.*x�7�!<�8�y��f�|2xF�vz�V7c�q+0�ؤ7KT���
��b�����oJ�J�*>�����s�U�< �� j�x�+��g�+4�9�*K�m�X�oZ���>}�͐_���f��t�I1Q-3�����c�:����İb߰�Ӌ��M�į�-�+�v��8�(w��:)⣄E���f/T�G� �AK��=�B�36!V�|���+>Ɓچ��i�6�ˊ!b��Q�P�߁����u�`&hޞ�<��~c��o��7�v���%7P^sWcf���#�X?2�u�.L�������Ɔ���L��	j>-*�\U�b-Cq�����#�*j&�|'S�˽��a�j%F����r$�@�Uk�)|��V���&	�.������Q<0�);4��ΰu?|nY�K���s�T	3aǎ�V�@ϫ��+��N�Q%��宰5��#�,7�N;_��l*>߷z�L]�p�[]�J0�p��뜂����� �'I�m4��慪�ƯD{�$%��?M�d���/L�=<�-(M�����(<��<{�{�Pa���yK��%C$C�8x&��㓈a��͎+h���[���������В�-l��O����¾���4OR[�眩����:)�G_�� >��AvJ��l���K�I\���c[$[:۸O�%�.H�2 �,�.�\�ò� V�[�U���u��r��E��D�F��A㴼h�oq�~�kA��Y�ǋ�5l���\WV���XD|>vTЗ�=r?��G�����28�!��.@Ŗ{��>}�-Qlwų}3[F��<X���:Ӊ{I�����.S0��W@�Z���M�̲�8l,Fs롺]���Y4D������=Ҵ��!��Q}\F�hdGY��[�T�s����h��ߋ[�]��T;��2.��-<�q�Wk�Z?]M��,h�CT�D搇���[x���}��x�5ߴey�@���?�wL���q:��( ����Wj����9<[�=a�����9c�����ט�Ü�N!��Щ��cO�W\�y�-f�:=��k�(/>�v#f/���.6�;�2f����-�+Ό�ʇ�W�}=޴��mkB���-u�y��*���.�M�l�����y_S��^k��?^e�r���'��˸�ˤ��_��+*�T*qA{��C&+\�%h^3@�Pd��]�|���k�o;�k�r�IIi'2h�W�7�`��A��N���K�lS���-�&��"��H�����L�֝�jY�E,*��|q��<qZ�W942�� ��}���A9h����ZG���r�m��i۸��"�7!XltIV��eX�mf]aMNS���,��G���B��qY@�F�(�¹}ct�L��2��gZ%�瞏U���l#x���;$u�܇�5N'�M���|)�<������ޕ�]�;��*�E�͸i�"hŝ�t��K�QΡ���OT2�o�J&