��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K�&	UT.y�J6��}԰�c�"�� �.ŞtG%��\�&l�@%[(q��
�-Ћ3�E���_'�0���RqVw�{�v{D�|��*��C�HP����h�����+�>����6S�>'��]��U�7!���Q+~p�xʒ��2H-}�z�(��h\7����@|/D�͡n��!�h��e!;�<��8� ~YL�@�S�u	@�ܚ�Wmer�P���J٣)V�)���ه�����:�6ZtY���'��@�p���׺V9�9��/e=�>��`0�H�[�
���xi�ZcZ��ka�A�ϛ���.r��ş|��0U�L���܄@�`��o�J|>�~�����-E�ύ����S�֚��Sy�S�+�y]�P+_���Q���r�ޜK*($\�ᨰ>����0�P*6�f-d�9�&�&6�����c|f�w�P�Vq��k�R�PtJ�\;���p�'�o�� o�����A��8Wt�O�j�Y �]� ��l/n���E�h7���)o�Y*Ѵ�������$M�.\��"�X�i����l'��R<��#9Qϛ�We�c�k���b@��'�/��B�1�n0���u���_�N§[�t�Z��W�v��F��eg	/S-�1όQ[�4���<w)[�	� �k�N��jٯ�A�}��eb�#槛v=�:9��g�g����*g�# �T���~����'^�-\�Y��8����K��қވ�_�^E�*{�A�=��%�5*�X�3>a���UuG��KT��>�G��W�D���p��
��d��
w�xj:1��%l�i�5k�}x�Wץ�AhA�f�-<�d_u�e�*� !=f�/@�q�GY��4�l��V��-]��7k�e^{ z�O�3�kPI��ۊ�8��I(�G�ȕ�3J$`ۭ����GCq�j�� ���vWBR�u6A��3_/�G�+ �,���/ w{��[˂�<r7P���]"Ft�����A|�OT̯N��I���М���4Â˼�C\�Z� ��uumD�9n��:9FS��c��9X�vٴsO�e�,y��W>��T��/S�e�=�D��Zq�i0��ւ��C�?�㬣<�@^��ܛd�N�T~�	u9����'Y��%b��K��8��)1C��h���\S���4g��@��1����GI�/��xdF������UM=g��~��c��2� �:@6/����X�R�37[���s�^����كّ�	o�<�V��0��	Th?��k��u��{�J̢�v<C��͇
3ܗyj��}���|&g�'���4�W��i&Ȧf�Nx!��>�X+��9���MW���a�dq��_����v����M��%be�i��w0R�}��z���Q8���!�2��R�x�BN�R�tKf�]�;�e0��~��5 �ż���B��<�Ǆ���TO�����`N!��~�8u��S�KZ����/Iʝ;�(�s�s]�l�H�܉q97ȬC1ۥ�+X���Ƹ���b[�gQoSa�U� �1��OJ�
��7��v2�	 �M�[ ʐ�}�&���m;OP-dA��6�=B&N终�,^QcN���]U��U�ǩE�p�^s:������0m�,�c	5�I��48)���t�R�\X�h��1GU:m_���A41H�3MMpң���.|L�Sc��LP�nK֨o1��.0}Ϝ��8������'�L��*H�M�jB��7�5�?�������<q{�N��z2
?�D���F�g'SO�7%���v!��ؼ�*�4t0)ij�����M���&C��F��f|�T��O�L�بۻ���LA�I
'�(�g��X�Q����m��7�����z����_�8���ዙ��kA*��B3�kQ��<X�%���AO%��،�'FL zy�i�<�)�~w{5̂G;4����'2�@i�`�a�j�m2.Y[�w=�QX�Rc^�����a} h�������J9q�dj����O�
�ү��]R#l=���f%�E��J(�h�Z�j�S��#A���{��UJo<G�mv,�uU�ۋ�s꼗�FG٥u��|������]�I2��7��W?A��̠�����Ǆ� ���7*Yy�J_{�İ��I:{s��?d���@J����xD��-S�H��5��0q�yvst�1OW�O�l�#�6�&ʂM^�lM�UA���
3�|e�&,<���gL��K�[5tFF����p�k�1?���䀈���ş��b`�I �X79Є���k�������c؅�K`x���>i��2��<{�(�5�Q��cn� 9?�o=��oH~c6����P_WyЊ/�F���D���d٢9�8�i.6 :LV��ɰ��t��T�/<[�p�tL�wr��1*+<�G�DB,�ۈ!9媷[9�����S�->�p��``���˿E0a�����2�څ)�ԡ�2����5�~��J��q|bO��5�LIՕ
9O����FL���C�����[�}c�Ҁ�K��۩Kl$���og�b9`�x^�G��Au	�*I��`G����>ЩN�Y�����9�C��!�>��Hh0;ޗ�@�{��m�j��� �l���:���.g��!�@�Hg>����o�	�t�D%�lZg�G�
�4����(��Os��["�jH�B�8jx����ڝ�5�L��t��H���l=_�+�݇��u}�w�s"E�%�V-�:��#���K6K6n^O���
�Op�~�J�Ġ��n��xEڧ��T�Y%Y���h�R��D|�v����+�8���L_H=B)���uO�%R4en]qGjμ��2��<zD�	���jaՂ0F�K�|j[Š{�K:��̈́���N�S{��C|�lr�&���R�r��%-B؅dۆl�W��Q�Plq�}�FSJ`V�ŖBvg�A�	����y�@�x��g��wyv�t|$�}8T[l�v��d��5i|&uϾt���_�k3�ny�jA}�1����n)3|��qm�$������r�2p�n١�e�c����eQ#��KY^�t�	�^��-���� ��;H�jH�
?z|p�4���ZIh��a
�X����@��L?�?��c�J�[5x�۲��$5�R~�mH�}ĄhS���������`��E�ʦ��U��h�:��O�r��sJ���^�M��_�,?G�6��j�ꓒ��!{�1���XuRq�(}�����l\��zp;�5ykC�A�Aޢ�LS�H��X+�:H#3�<~7���,wF��JlZ��z�������A�;c3�h��)O���9�k|���7@���^ƙ�7;.S��oT��}��S�3a\iQ����P�'$�����<$�ڽ�:g����t��V��]��|�=;��O�B�J�D�rѿLֱe��#R�@�� gv�������A�B6(`�[KtRT�	����aB�]wq����l���>��V�����r"OL��_:(}��ՍJ�"�fM!� Y�h�3��{���"L�&�J0�N��V�LM��_?�M
�Q�����:��3 G�8�Ȣ�
� �	�0D����L�qw��b��R�B-���A(�H:�9��|@�ܑ=JB������W��}����A�1iZ*Wm�]i�����^�mQ�w�ũQ�V���}j�ai���6>���>���uH�T�ߘVN�2O�4���m¶�ֺ��5��焄�'�ti竐]��O�����w�$�M�.�������0���n2�2o�<0�}�3*��s#�neI�]���@�v�y���OP��r�xZ?�Y@\�T3C�<��I̸8��U�s�TF�$�r= �v��MwN�n��@�P���ϙs��t�;�"-�D1 G؈eZZq�.8c������$�A`�ZU��@�jOl��Z����ںv3����Yq̅k�1)�%q�.��S��և�j.�+=�����Ug���F�@T$���v�
�#[���v-�C�isЊA� �������*�
��ؕ\����m��2k[� `��/F��(�4��Y�<l�8Q`�2~�jM�~��ƈ��|��Z�8���s=�S ��&|D�������z�`��c�6�=�vq��6�rh�yY����{-�����UQ9s���E�寅�������.#Y���`k}���	���Ͱ�����$D���DrmNu���ΰ��M�!�Ook9�_>R(��̻:������y�坧�!�*L�~Q���͒RF��"GY�6~��8����vF�sZ�ϧS �9ϫ2�ӇB������Tga/��_���i��^����Z+`��(?1p�?Yt&�錵��Y<v�yW�W,M��u���f胈6�+a�˯	��_GF�mn�[%�0i,!�˦���=D�Z��,ew�L;���a���\��oJ��<sm<���4�ʗ�IO�dgVY��d�C�4վ8�ܸ����Sڶ���p6���S݂�+s&��4�:�4n�k�����l��:t(q{��� ���)Rg�[kE���A��6���J=��b���f�Tl6��zHn��i���6��k�<?4�V�N�.J�J�v�^Hc@���K�~U�Ko����e������kܫ�G�#mh��;��%aL���H�,�N�H��@�	Q��Ok;�A��u���F���>�T
���o����S�|(�ܦ]�HV��[������$�g,;tY�킺��ΈQ�s�� 3g��K�ѷ@�����o�ōG�sb�@�X�N~�?*������\���u�;JA�(����uS=����;L�����Z�\�p�Km���IV�k-h��M�}����4'�4ĖW 
��R}��Φ%VJ�Q���¨fp���CJ�J��>3��kH�li
�iW�q_�C�<����9�t�R%JƮ�gm���H>/���A]��Nx���IUs��K�qga���,��;��-MQH�+m�N�>��a
੠3!�E�
m�r�o��m"C�hF��֗{��@��/���'V�jq����S6���O��@N�lUi���J\c%��Km�J�3�&��xL+��� �[xfW�F��A�#́e�A��A)rYj$StN�M�\f��p�&���-���S��-�:����b7�^p'�7S_9;���X��W6�6{����x���w�����U�{�;���P��?Ȩ-�� �O>�~��2����t{(hH�߳���i��q����c�!0����w��P�h��u���\�������5_���Ҙ0��3�)����e�)f'�G�S\���.�������`(v����x��7(+�1����@�BA�=�"��V��b��<s/����Ļ�7N������ь�F���%x�'�T���T��r���!���=����G�4b��7c��
�Z`��	�,�T+�p\���R�oi��J�<��4�4�����}�Ӻ(�h�b=�P�v.��{�[L<��s���bB)7�ܳ	fj�7 �65�"�T��<g��V�K�q¹y"e�0���J� �� ��|�r{ZtƗ}�s��%F���W]y�<��p>Z 
qTJw�Nє���3"��M�q�K���GnhQ�+H�p@Փ\�0L��5�&�Mev���?Q�`��'&J��Fm D1k���xk��t!f5M=lF<'�����������+�剳�+�]W�I���$B�_�Ղ;��Q�ht���i q�y��������e�z�6��s��{�f�9������8k34 �:Y�6(��-G%;8���8*ͩ�� 1�gH����_����(��ye�!��wn���z	�u老��ۚ�樿�a��  `I	��?���L*���;�nbT�S�������j�
�yh������1�ֱ�SW9z,;��kK���:H�|�xj��+��>"�i`�<�m�h'cVPnvo�A8�#�#�8��n��=U��1��7�IC�Ky����	���h�t0��\C���Q�\}o��T3�nf��H��V^Et�������O{3��,��>9���a�h��
�Ѧ.����~�����ȼ��_4 Ǉ��Ozߒ��n�&�v��X��2gD�z:S�5��n	�>>��i?���i�)�F<(_��ՇK��a/�cR,�g�z��,A�?�4+u�")1���q�uw�����:�w)��q%ro�V�i�8It��1g%'����=Iz�3C�L����ҕ�K�ed3�����M.[n��{�	2G՞�1j]V�~o����F�@[!gnN�~~(��r{)�2�2لoUqd
�^H��EBZ����*�w�uv�����\ 򐃲Cm1��䦌WMi�HO$�9C��J�Pmu-2�	m�?f"y�!O�)�d{(Ս����	�;FB��'�łJi~��A��~��0���6g�д���o��kT���70[�
����f/s�b�>d8B������Z,ҡ���s�H�V�sc�<x��FA���p������Щ�eUU��gĜ�b0Cȗ����4s���{�kӱ��V�IO}�������X�K~Q�忖�A�����_hW���D�ލ����5�&g�N��FJ�eu��pUr���GD���m�Cfʍ�(27�F�0�n�=��k孭��?8M|+W�w��FЌۢ�oL����KWY�xx�e`�K�V�{����BY�ʲp����Պ��ȇ3����/��#S����iM|��t�,�GQ~���rPľIGd�%= �Uɹy�+`�y%7�����c���f"�N������[D�Y١�^Hk�*֞׋B���jh}����ț'�r������Ob����F/��k��qB��[2�1"���#��)��=e�����Uf���߰·c�tbw�4�It���×#�Z�vDn�2K��k3)___��j����� �Z�����#�;�}�/�����Cb�)ܢ_�l�!�ێW�]j���� Ϙ�jīT�K"�YDc��c�Vw_�� ��˪����zP��c�)��Q�C	�bNѿ�4t���z����<�ǣ�Џ�� X����C+�36D��"膮=$�v�WNϐ`adN6x�\2k�R���b/����LH6=����� 0,cNA��bS��~}�!�<�j=oA��MДE��.����v�6�����<p��-�W��d��o|147l��j��2������6�i�>�97��+����ܛ+Sl����ՠ޽�p����Y+�dU�FuVkE|�?�� *P
����"s;�Z9}x39�Ȧ 0�����'���Hy}ð�8��-�}	��ţ���J������! y�&)�d܀K3ZI�'
/SȈ�L��zy��p���ߩB/�f��&/��w�m4�;�x������b:'�u�&�x�7o�<��-~��9��b�F5���z��2~��>"�"����X�y��� �&	2���t��%ݭQ�������i�;��1\��a"D��=�g�Uc$��i �)e���LN���B�9t���C*�}Z�]s$B�,�N`St��?#��'xgW厦u���{��3 �u	I�X\�>մ�<M���e���@:�Wu�{�Z��{���1��E����1�������т���,��5��JA���R>RV������{6��_E�M���ev?&�x��f�m�رS�o���DRro t�o�]��ǲ�IQk�Y��^a��8
�&<�
�jD}�VH'y ��E;``V���L�1%��owV� �SK�����͢�ؿs�2�Z:��T(��Ä�.� ��GRJ�Y�. X�_cߟW^ �,�5$� �A���n��j��}/��[�-���W�o	����A&�ߓx{��Y��8a��A���+�Hq�@�5������p ��dݱLé:?zI��a l� ��v�b���[ ��x�����,����w����;[�G'�]AךEr�K�Tj�Z3pm�-�̹C2�~PE]����ьJp�̡t���w���B���FG:�"T�^5a������c���.��ٞ�Mz�q�`
'y��}�i�����3�Tա�#{9?^������sE����d�$�#�� <y�lv��X��q��f�U�%�?U�'���P�T�@gh%�9IC����D��2��.)4=�0�⦞ƻx�l��r�j
��.����:��M����GrL9����c�W����!�P��������'��n�-���/r���f�>(d�+.H�!<���s�`��Jd���þ��E��h���O�� @6Ȥ �n���������Z]��(�J��bǨ���^����_v�'IP�0ZFRH�q1�
��YA21U�Wd�,��^��Y��Rn�04�He|���B��p�$%6A��Jm3��e��T.:��y�a���������C��Ic�_?�0�l&���?A8����`h���Z�_5M~��������.�z��y�e~�OA�ܾ������vn��Y-�苋��]������"�ΏuF��1��g�ٟ����ě���7s�����m�� %Ҿ��A��c#�w.����S;Fo