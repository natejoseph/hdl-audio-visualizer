��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��i�X��}��ϥZ)��eD�De�Ůᒹ��7_����?A�;�����#o�[m���sAٌP�*V�<��;R#�m�[���)?M\����,@��;XV~s�c�״G΂8��^%�TY��������0�U/�铯.�g/��ۍ�P&܎ck�1��Ѣ�MЦ���f�W������'9��&��3�G�y��LI�����~`���y`h��35Z|��Z:���i�K2$�P᩻���3�KQ�4Qn*������J��%	uI@۱l/O�xo7lD��K\����F�D�W����78J�l:(�/D�E�4a��GW�j!u�N����:y�rOwP��>�'KJ8Q�5����O���+�>ԲcT�_��l[q�;���:;L`�0�H��jE"��řIŠ��+dU�ǌ|h���T��P��{6�>��>e}�����!�����#*�S�pDM1�E�-�j��ֳ�QC�
��*�>�(���*�0T�3u����<|�GD��oޣ��*��i9��i�%h^��������D��}~ �úBq���[Uw?q�=��i&�2����l6�}��vq���n�x@<[��4S�.Y�}�@?��4����Z�)[c�Y�%�9{l�H������|f�S��4����3�-?U	U";�7W��o����3��6S� ��}?�H�(�J�;�i����m�"��'h����|�������d��0�+�0�E�1�2@��
}�c#�KGCMv aA�듅Q8t:`p����"hvLh��즯��1���$�a֑&u�;S�������p�uߕթ$�ɾ'�'��Q��pO���͂�"L�	�zF�}�� ϱ��L��E;��x^�c�>������3��J��C�#L�03�jƄum��s�v��?�qX�Јʗ�G���J����5��T0v�Դkwg�����k��f�O��� c�dW��s;X+�3��cCؚ�&���A�?���'�ҺwXۦ:��85ї*WKQ?�F���w�`̃؍^�,RLv'�a�t:���8�� +���e	
��)^��ӌ�������Y�i����%ny6��5���AA�3�zOoxre�7b���N�f���.�l�-Y����JE�AW��ؽq��
��W"`�C?�?�؛_(V����P�!���9cAo�+
'�?����B�0���@b,��M�ͼ�@���m��Ԓ���(@6�ӏ�N��#�`�c��s�"$Xp���#�RM���3� �q�]sT�EsE|_�U7k��Qu��l�fif�e��#G��;�V��ͧi�f}�g����P��g`�����H���ٌ��¤c%οʐ��em$��ē�z���
�n��G�i1�vF��J�k�b�w�kw��!	wл"�S�d�Vy��2Q�_�n�Ҷ���-v�b�ht���P� �֕��\,��^{�v��*{,���_��B;�~�T��SlH��F�Y���\|��o �X��UΡs�R�������f~H�D\>�����ﮗ5>��1�Jz�ً���v#����]�Nh���2�r�ٰ�5�֝)|��38k/��2.d�����[�E�zI˲_�5���Ҳid���/�na���2�[d:y�YA,������b��L �q��L�B�U��x�w��"�lYG�*����̨�u�y)���kR�I4i��x�E�y�]~���v���%��NZ�S�?q@}����z��r��=I	-�D�;?]��Zae!Ι�Zh_S�r�a�M]�%- J����kA9|KĀ�$��F�ɠ���s�:!�� ��i�'��^�[)"�]Y~;9:��Ƹi���-�ȡuթ��vܿ>˨�.h�ҴY��1)�9R9��$\  ծ��մ�E�-���:�"�R�c��r+\b{�^c+r�)��vvK��yS��Q�N�G�)B��>$%�A�x��h���Q��	��* n!di���\d�7r�=x���������l{�N��q�� ���\{+K���ӟϥ�-��_9������l>��uчU<�}g��Jx�X�ņBx$�>6h�^ut��pq��u��y�"KRp#�oE'K�\���s7�����ϯ�,�֜��)��0�l���M&t a�K��GPS�d���.���T��S��>�
��=�`���D��j�mw��;U�V� ��B2E���_-U`�U�7_��Wa��qM+6��O��L�|�|v�W��Ε"<#{ŉn5vF8�1=�����pz89V���ۘ�a���_9�_��hb�����۵��u�M�����4�QfGݶ�ln\l *��ތN�҈�F�
iD���x]�B,��8!W۸����ip���X�T��L��*�]8������O�S3��d��݃v6r�4 p�n/Ɍ~>���Dr���6�q���5]�iV���4��bSAƀ����Mb��+e�.��i|������������K���6Kthk����}�>b�K.wt"ܶY}��h��r5.`�ah�7��f�Bf9�wG7>7�&�� �Z�P���,ޛT,o��������C��1�	ȢG�*�]!2e�,B%����	cﭿ?� �@]�D�
-��u���Wl�xO����Y#�\��Ua=���NA����*d����w�Y���W��S�i](�Lh�W���r�'�/�����9��s��)q�����U�3���t��1Y��XtU��r$�
श(X�QX
�D^��דn���2pZ�C�*�
�03��V�lS[�.E�^M�Pj��Ar~��)�a[��6~�=[����?��2ɀ�=��dM @7�R���"��8lND�Gf�҆3u�!
�G��4��8�����DK�����f�0�T��ɣ1"����P|Ȍ�0��I�\��S��r]Y�����Gu=��"ݷa���:�I�qt}]M�����5��K%�Y0� /U����x�{x�y�]jp�LZ�^E'Y6�%����w���j���z��o�k�L�k��;Ӳ��6/���~j!;S���B@KOTy,�D��y儞5>����J�Уܬ�W���fX)tLw��g/��`X�h�24�dL�|#�GRa�y!�˾��u�R���nv������f>ֽB���YܰJG}4$L��מ�p�\\d�4���n�-�:�,�EN�N,ymZ���"Ha�8�m���l ���h�� �J�`x��ab�񞊅� �m�����v�k�/`��G<9ސ��7�Ǝf��g�Ѳ� ��>�e����G,&G���qMvj�x/m��^Ԃ�Il��cÐj�����9,s_b�2jB��ߑ�a�7Cc��E��ͯ�;e�1�����>���5<+F�](�^t�+P�BȟX�-����̲�C&�׌h��(1J�
t��kN|ʠ`�p�ĉ�6f<�)[#�<��8�j~���gt�sEt�c`�]ODD�޴��j��;�*�?.>Ù�|�]ɇq��VI�W��z���f�=�-��3{G��.���z�]�^g>�^/��������J�_�)�@	�ӯ|�  4�c~�PM������a�JI��W�S�w�Z �];�#�!��p̻iD`UB1O�1�*\ur��:��7o���x��v���iyR�<�g�a-Y�Iu|��_�Uͭ�*ԍ��@o�yQ����Ͷ�vR�i}�TN�**�QW��&�JݚS��W�oں�xEԌ�I_
ҁ�gv���oۭ	7�ƛT:��c~pʙ3VPg�"K�7~����^��u��̏-�3���w�S@���dia�rP_���tܿ ��\����(�Sѳk�n\g���Ƞ�����ڬ�{֔�%Z�ٜ3���H:"����ԙ����ʴ�L~nǞ���L�s�"����&�fwH?S̺}�8p�B���]�H�&�~띶=����GKr�1��0�Ļp���5;��������l�`rMhƭ!Q�#7�<Ɣa��mu[{����Cif/�Ls�ec &&���յ��#��'*ǁ�������=��K� p�ev���z6�X������3aJ����nŻ��0�a�M��84�oFG�w�ڧ�L���vl�K_6k^]�1t|sR
�+aܴx�/y��/�^qH��i�9�*qȈ��N\ǻ_����"��g����zŵ�gZ}*"=[�pno���*\䑰���qFFn�Ð5'9�-O�5|6,d�_��?Q���1&̙ի�%��$�E�Wn�K�_���бF��ꉠ�±�qnmG��U��R�G�U2v�ۿ��v�R�8Ҍ^�t�f�BB˞��i�A��!���,���~�z�@��8�$�b�<Sp�C�^4��g9E����F2V�Bj9Y>��۵�:�����Y�y���>P���j�����-�Dm���g� �ww^��0���d!еv]80���ӧ ts&}{�����D�ǡ�9}l.."ނ���3;Y�(�o�2ȞJN�@^_�H����R؁�\4^f���2}���~#��a�X5��j .�TK��V�J�3��^��J�������7��x&�`��?KT��?��/k6��7�e��l��ԅ�/�Z̔B��滋�s���]��;�z��h�5�D7NÄ/�Ո�<j���X~�U����Z�#47�!_�[��5�s Z/��q����m�Qn�7��A�׋V���I�P�%�AcS"C}}�2۶_<Sx\�gY'VL��ұM��O�
R�@��V�B�@��
3��HQ�b�'X�E������ rd��hZ��#R��*��	&F=�o��8�Bx�/i�R�Yq�*GB�.����i��NQ�-�)F��{  ����؂� `ӡ>E�c}�5X4B���V�q�|���8�ˈ�c*;�,J���'��?�5M.L���Y�ڃ�,j�"�p���8��}{j:���4)����sQj����wT$�([5�8�H�+�e
�����<�9V����`�v. �}��L%��`.6S�yf_.����B�VrgQ�o��LCSɒO���N�%e�hlO����إ
&9G%���³.uQ�^�-&�i-X�@�xҠS�g��1�W���ٷ#�����؞a�)(Oj(�@�m�:V]xVOf#k�bs��:�ގ%S-�Di�/�k��qy�'�f>ſ�����zB���n��U�?�C�^O���T��)���Np��hl��Z�I�8�� �zT0��3sɜj|�C�@E_�<�B����+	n D�!�GeV��B,j���P��|��#�(�~J���p�MP~ڲ]���#�__�|¼R����;b�3�-j���;��+�d^�.8�+r!F>�i�ӻ��16� w�����Ip�����l&�9�C�F���!�#����>ȉ"�%��K7eGu��g�RM��ր��E�½�JLh�A屹�E]6��ދ[' <ޓ�<y�@��<��X�5����<�Ҿ x$�>I�O�%�JV����-�i�y�f��q�r��NIѝ�+�`D� 2{~8�:Xu������\5C���¿�mi~\D��cq�m�(����y���G"{m����G��_9ǋp�ԣ�_C��Ҝ3&�axkW�n�g�SʟY��h�A{�ء+� o,m�I�j�=d@#��4�pt�oх��_w��Vu���@u�`;��2���_��[%�]���c���o��
��t4D߫어Y%�u/\$$���$V���IN��]y�jIl��:�?06066�(���g�%r���]�8�!S4�%��ŲL��q��9����Nb�f��2���p@#޶�r�}�ėZ�h�3^k�x#c8u���.�6�N���D�Nyʷ�U����\t�uHD\;'r�Lc��Q_>�w�n��VG_���c��-�8�D�`W7�ܺ�m���f�=lM�{���4�!U�2��K�y	��\��������H�n�v��R�?0�L��G՛c���N
���O�S�������&�>ZϭdН$Q�@��p���d^��<�S!p�lpD��M� �[.6���&֋��~�������G������ڦt�>:�&H͚���G:��߇�^>����s~����MJs�ѝĵx�����S���u�aF�5�K&]�dX�����/�A"������%�d����H����M�Rb&���
x���ުr0�]^���ͼ����~�o'J�ԇ�f�ցq!|4Jz�J��W9T�>��^t	����B��'ُz�_�!^M��d;E\X�6���%	�M):]�E�т��(��@=D��'Ԋx]�K��-�*���~4+�AK>��60��9h�i@s�j��"��T�t����`�'�m?�9�TxO�wrt�l����^����U�N68F���Sh�~�o$�h�٥�z�r4P��{�^d�!v�3�oO��IeDY��iW0}��L������hl$差����T'N-Py�c�Ԧ/u�.��_��/�rhB�Uoe��{�%���O�팚���i/��4𳑒,��/F�?��c�E3�f:��ts�������q�������λ�I{"Y��"H!'r����N�eF_����x�74����xXas�<p��i+�y�I>�����v���g'ss��;F{����ǁ�>XU@&���}�ζ�e:P��,<��HJ0�`o�Q<<��~lq0u�����:Q�r7�D6�Q�F�X�pR��.TڌQ{d�1x��?.�� ��g�6d�h�;���r�H�{���F��
=���YsS<U�[����BFn�,nm!Le��,ʝ��a$��-���Q$v6�y2�֊0��~�f#7g�Mn2<���%@;��Mx�[����/�ڒ�;O��iX�%rE���C����*\'�M����Z|�����z令�k��E��!��qX�#��"��˚a�o��MMN�y���O��Y��'_�Tyb��D��;z��Q�3��G�?n�o��,S.ןTNL�2��o1.��O��"�r%�1�P���L�����D�7� 8Ycg��e=�x^[��E<���6 �4�	��g�Voݮ�s����kz3��#&����2�Sp)�(*�u�N�}�r�E�B��x��/m5{�aLp E8MD��d�J�)����YvS��3(QJ�8Q�m����V�������	��/x�-�,US7wV�Ƚ��L�œ���3�\"ie�u`�&73x��Gj�;vӷ��\���j�#,�ប�:�܋��`���[lb�^�D���3}+XzY�����E;����A�:�ERM0�6�C.Go'(ѓ(��͎@ͩo���Jz0�z��ukm�:��߅��tE5|L��}4��M�&�7_�/Kk�/�':ͦ�"�����h�������q\��^���M�{�<����OVZ~{�.��q+���=B���n��u��-V�r*4l+Ϗ[y^�e~�9^�ܢ+h̆"J|	>6�cP'�)̯E��!�.,�M�ut��]�݆�� j��"��V@�i�Y�ΜsUM�&�*�QJFk��$���@F>��������e�&�!s�q���d0�<���|�Xta��\�%��N���x��bՈT�h4�C-
�+�i �MA�)N��5�螼��Dj(�E^�D��p���	�[Hj<�BJy(s�̱�zT#�����>���� ��0��4��%Q��a5���Y<��R�<qnl��'�9WB/�Z�j���x��m��n"g��j�?�P�������Q:�@П�bFҹ�b7/�S
��`���o$�������24+>ҭ��غ�4��Vl�g�dr��3���-���=15^ͯoJ"J�I�g1*��(
�_�mݧz�u�{!=�.�OԛIf��78k��|6+�2�jo��!���x�уn(�3��nC���N;�g����y)��y�#����|O&7��,��g��"�2�Q����> L����R}���ۼ^���v)0�=�\��CR\��#�aD�\�z����DB��S�7���,�+q9��:ųɖ�Uv]S1H&���҉�RM���Y"V��F���9���͐PޚM|/BS�J���*��4�I�قUH��9�饖�Y�s�i6Ӏ� r;3@G\��;��y j��$'�F)�8��+p�~�\]�O ����M�k�I��G���-kl�	&O8,�~�ձ�5�n����s'p9Z�����!��
~�8B?��k2��Rm�����iF�s0��8�FS^n���X��q����mw�[&Z��{���V�8ɫ����̀0�9�H��?׼�^��Hi`��%��hsH,2��OC
�ݤn����0V���Z}��i�j���4��t1D�Y�P|³E'�}s���p�*���'t$��M�������j)rf^��;"PiF`j¸�%}o�nw~̡�Xz.��ίsO���[Ď���h�V�^�r�v3L�<DjV��b�	C�ڦ�(zS���a�Ǝ����C�W�xZ;q��&�{��6�Mq(D=����h������Ӌ4-�`XX���XT5䮴m�	���9�s�">�v�>)\/ZM��0xݛ�/����*��A���ĿC����T���c� ӈ����(�E���/߿���c�������NՉ�5�Mд�&��K:#-���w���ȽO�?��{�o3���h&��h�+��W�
�S{[��X�Eq��X[��A�˛�]��)�a�Q����`�A�H@^���|�>�@���?�r��q��9(*�m�������0���#�0��qb���Y��J2�s`孖�\��P��	S�>a�\�S7e<ܕG��,�IJ$f�e6KQ�X��4�P �l �	ltn����/B���ę�"�8ϲ:��a�.�c�_�l$�(��8������7|�<*�Y�$����(}���6b�,���j�6f�6��ɢϋD�����O��81�I��ڒ�����;Z�t ���X��30�1$���j���壾st$��&ì�7f�!����#pkI���Ț�jU���#���ۍ�_מ��Q�u�o	aI��i~��N�k���'H!tt����=��DU��%Ň������ޭ�Yg��$������o�����L[*�ўyR�f�M�u�*��G ����{��f���q�ÓUx�{*��������_Y�R�� ������er�`9}t��=�����EqO��[&��͡	 +	{��(�j`I�m�g�=��
Sr)��h#��[�/r��b���t5�������uΥ:�i[@9��>�$�p�/�]���	�OV��%nIa�{Z[T�4xQ�H���b3p��y�Q�t�sϦ%��r���:��z��Ä����	�ܬ�)��K������|�ҹ�����2�K��c|$ɸ���	]�j��ֆ�4q�M,+��Y��֬���mK`�_��q�'ޡ�$�:����.�&E�ƥ�����5�'����q`@Ϗu�"�m�JL��ke�D�`��cu7���bH�(۹��ݼj���_:����udI<z���}�`h��8�:-!���v��%��������b���|�%�+�A�	1��hb@�!,YL��Kjϑ�]f QZm��8c=��+�eRX�:�fx��[���M k$.^��؆<u�F:���}ݮP���tLR�>T9�;�G�ۺϗ�{�yvV(��Զ�<��R47�s�Y࠘O{p�`�fC��>k�A��*�P�VY{�߰�S��;��m��#L�3�}{���߂l���4:e�5�CFBB���ʺ����1������?t�d�YQ�䶢�@Sw���SӐIVgP������v���1�SM���?���59_�;�g�!}���e48jH�����Z��.Z#6� �WQ�D\��xO9"Tj���x���J��b4���B.<0�����#ˉ�o�q+,���I��dL*������aH/����@$�e����8JR;�0�?���(�#����{�O�%˕��������F�!��K�E��ʮI����
�/
�[z�3EB7@[SHp�V��o���B�B
s���lSa��f�@��.�A��� �Yi�u�:�`�i����]s�p��<Z�U>�OĪ�
{-�<�cȭ�O�.�X�/C���&
#���e��o����\��pu�Q��̦E���(Z����.�R��� s@��u�&�S����CU�9����H�g�&����a����r�\)!tɎ�����ŎB�ƻK�Z��r!�����հό��Z*D��y,7�H�9] O�v3^j�A&�ȋi�ֱ@?M	��uށ"$Z�Ilt~�J������E��_��v˸�+�f�U�Ҵ��mcd`0���%)�oW����	����d)VW�+8(Zb,�����.o4qo`"ܥ`0(�0���Z�c��s�IxF���@욃ˉV��ghZ������+�D��$	��ђ�L�DI�h	D�-n����H,��r@2 �9��;��o#��&t���(�H�Nࡣ��):� y&r���%�Dxt�Da�Fp6"
8ݜ�X7(�ԕa,�o�B1. ]�Z,�z���9�j����)k�Q]��Q�����LP$�a�u���W�Ɵ���W*F�� K -�&;y�R�!��y�?(�lT�=ҥ���>��P�&��EFi�`��ī���/O]F�cce�J������@�9%�/�l�q=�Ɏ�N���5���,��*��	���Z��!1qj�D�ŨK�� vX�����#ze����2�<yٝ#�O6cXj���Ui�LՕm����00v�L�����T�"�(E�k̯qo���8�dwlS�$������r�#���S)"�}q����kX��%�$z����R�(/�P�u-X���F��oZ�!@��=����$ �=��/��}x�u�w=�C����U{�<.�i6V�b�J�^>�=�s ��p�BY��޶l�;�=m�t2?�-mp'l_��Q�i�P�-_tn�4��NyϷRq�^��Y��'���_�W�@b����R ۼ���<~�b�ٖ�s�/���%���#�5�<6�]�+��%�&v���)�
�^��
�r���5�\��؀��[$ˌ��%������й��%m��V"?�5�G���=ފ��˾Ƒ5ׯ��8�)�Y%�l�x$s��P}4z_Z�2���u���̦q6��Y쒅m%�C�odRg�d�����YzX�?�Ӯ	P����G�eD��v���8�؃���ƜS�p�w��wNn����Za��k��]XKrn�+�f��nbQT��9�v3+EUfKN+&��M�!Ol�� �!z�ɭwʄv"t��l:�I�3��+�n
GbdT�6��5���!����d<ʧ��}�����}���ײ-���e�T�7^�g�j�dw���C�σ~a$�YT�q ���@~�� �ϙƄ���h>l./u�e�5_�