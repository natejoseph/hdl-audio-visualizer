��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��S3x�K����c~��ln\ah@ד�/ș���3d�?>������\�5����@�H\o��\s7w����0��K��#F8��o} V����\� �\IDjVs�']����0�ŨA�'��8<_V><&fmCt���0Հ�f~���=z!D��V�:��a�_n�	�\0k�4���[����P<|��QB�Q�CϣP�=���@s�%6��[��o����0��wnJ�W��hî�K=ӺdԚ-��qkNO6�h�p�O�U���'�k�3)L! ^d��%=� Hg�#�vU6�k~Xw&b�*�0>����9[<���o/$!���"�0Q��	���N��F���܆7e�H�a\�S=I�'=
#��D�qu�fO}�q��xkz���Bw��ː�����R����f�T�R�O�,�U���4�$�h!��P\�K����vU�q�j�Z��2��;�|���ܭ�R�H5��!nѯyί���6嶄g�C����Y��oc���k�3��c+����IB���R:N�TG��WF!����z�.Rg��U\y�����r�(:��H�a�%=K�C

��k`��� �A.�}B0��� ��A��(��߲���tvjW����-J�4m�+X�����U�f��"�T�穪��^�2�{����o2��߮3�5�tD�UP�e�jm�a��b��������bt�C�c}���l�9� n��wG�5�����j��fv����k�F�~��Yk�ϴ�a���]�$eک��c�q�0���6z��$��}S"���}2�a�M�E�����|�F�a�%%"�I�⥦�$�s�9ot��^�y�w*���
oaz�������	r!E�_��^����F�־\�Q�h�fP���C�yW9nϷW��Sden���d"AE��J�CΡ���U
#�*!\�B�"a�_�q�VZ�۱�iOK��6�fD�<(��r�z���u+h�CfZ���i�%��ġ�yX�f �x��O3�&�\�s��U<L��%D���E4��)�U�k���\���8�����
9*8�ȗ�������c\W`�6@ͣ�G��Ҙ�jހ���~ύ=�'>��1o��D<����Z����
2泚�f����3�ӞX�+׋����p��ף5i�UY���G`��䙛 ��Ks�	�!��,��a%l�d�i�5��``m�����؜��Xc�+l��5�$U>�?6;bJ�|9����D�w0)Y�`����
�!W�,q$ٺʴ"����m�a-2��Khlh��U����B+�F�����h���<3S@@��N"53��hC9z/�1���ȃ�-n�o�"$<�5l��"��l��Oӯ ��3��)�8k�����9�������8�Vej<��(t�)�������λ�<����S���+Ɯ� �
u�^�4v/��(&�[��>��g