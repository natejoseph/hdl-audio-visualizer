��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��S3x�K�F/N�B�;����[���3�v��������tt�C���	��%�o$�-g��X"�cNg�KN�R�am|������P�BZ�_oM==>�|īR����n��;����Q����_��^TB:Y�DQy���������늊��VjTd���v���ࣉ@�ra���_'������ЦB���#sQ�FKi�d_E�9^�Y�� Q��V~���>� ��!b��>������.�}"~y�%��UP�ܯ�UN�UT�\"V֪M��\�}�`1��Z'ȷ��o�ѷ*ёD��7�/R
_2s׉(p�Ǹ��{U�8[��Q'5��5':� ��z#���K����j��k���\6b��2�Ε��.%���U�OCH�ڛ���S`��(��L��Fe���V�4����;��&e�s����9�r0�%�H�1��+�3���N��x�����i�[�\�:��_�S#E͌��{��*^�\0��U��&�:�*����b�I�*���u�.�����e�/X_���<\�qu�:	���{���rg���{9J1D���%�A4�@��ڌ]�X^�/Aa;���ɼ�5��\e;X;��G�쎳+�����:��!#�<=��ݹ�z��3=�����HC{Uk�=2�8�0/R��R%�Ø��u���l�'�3&Kְ�΍X�F	�e���~�Q-7�X8 �Wy�~�-�*�ė}��t���ç�:�OĊ�X�jU��㸨��L�Դ
�6�H�j粎&�]�:�����ښ�ʄye��30|�V�&���w*��?+!�
/n�p�շ�Hgs'�[	��l�4�_\rM���Xԙ��EVl�P��3mpɛh��~�"dN�?�@��*�F�(W����M��5Hq��HT����v��x��;�*�x�15���{T"qP�u�l�wQ\&���o* +�%87'5W�dD�s ӕ������)�GF.�;ǩ�����ZjE��hC��3_����ބ������A�vnhH�N��v�F�cq�qM�)(��Aq��s��)����Q�п�i"�d��F���b�A*�0�DoԴ���:"aW�υ��A�K�����t�"�Z���xBʳ�h�f�����Z>%��=~1c�Ŧ�.��=��-��يM^vD��F�v|g��rZ��K*��ׄCwO{�����m�X �Q��n�\K�5�N���Y.�U�!2�7�&����*[�g�	֎��m�t��&�bd8�a3?l�Sl�IBK�<�WOEl�b^�(��ol��?�=���.87�F�z��ҡ�Ʋ��B'"��C���0-��	/K�$�N��1H�4��q{��<�?�������4g�8���k�Y��Ĩ�
cZHGDw>]YR�N����5t2 ���'^�:-�4�̲+���-�b�+77N���h��n�P��F"'����]�Yp㞌��{�i��@#.����uZ����W44jgaO�S�t���z���n