��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��=HAW�dn���"���1G�V��K��{r�4�t�?����@7�ē�t�}P�?��l����C Lx����k\�����KԎ������Z����ȵ�`V�0�HW��)}�P�ӉE! 8��DOjpx�٠�~����J�	��h��vs�wu�0ZuA���;�<~�s�%ݜ���mM����/$4�-!ɓ~�$cY=�p�K��M���&�r��'r0��sH��3~M�:ťę��C��ק!LsW���u"��.R�IT�и������������·J�a��Җ��*K�r9�Rw� Z�n��`�U��/�^p6.���TtTw+O�6*2Xq`D}$�j���ZsK�{���S���j-����3ޤ�Y��䕝�+-�qhJ=�Bܩ\j��R�K�F�|L':���^��X%�SU�����/���}+�_���{��o��\^�'�P�-��l�rC�[�]�T��CE?.��N
T.@r���C���I���vU��!0�Q�y�����9����~�|�׫����\��*���g��_n]4GV_Pc���
��*��U��14ϧ؁ۄX}���J�	�^�Y�R���㋌wa۵����)����al({�3/1�f�A)�C��Ӭ�3�s1�D�pᡛ�]$�rŔ��ճ�Q��I7����s�a^����^~Kږ�A�%W�OQ�f���4F�����X.\�zPjP�D��Un�*O|�-'�j{����5~N�f���\��|%cmS佼�ѧ���>)e�g�':J�T��|���t22���[����a���Fx�ǖ?qڊ;��w�30�	)�b���!�.N^� P�F��X��bfC+o���ޢK|kU~����+dG�(��̗l����ÎM�O-��ECkqZ�l!����&o.o�t�}w���R�`�|�_��(93N#���e38�\�Q��E��ʪ�
�(�ﾌ���PV�8��� ��o��r=PQ�(r�}�`,]e�9��g�v2���\W��=�N�Q���y�[į�v��?P�:��K�8�z��4�$�M��d���&2_�����Vu��$�	�S�^Hk��5�����_�ϊ�d$��R�^�M�6�Ɣ�5f60��>���>��֔E���Ӗ-u2�]�����gYÙ%�6k~�?��`��-[i���J9\���i~J�_�Y�s�-i��Б��E?Y4��u�ۏ��D�Ң����%�ė;�4���?��P:�]�:p�jviaIdG�C!�2��}W؞
J�j�3��L�B,�C^��pX=Oj��,h仃�	b���q�Y��c�;�Wd�(� �Mm���jKQp��RR��O/:�t�qo����v��5R��p==[��׆��D�zQ{I}q�,kO�6BrC%�;�pGH��o ����S�u���w���v�0d�I�\�(��Ȕ���<�y�e��R߼���$s�tf��Y��U'ۨ�Ŏ��CL��\���@����`��V�}J���M�|j��I�S�r�� ��V�y��s���1T�փH�A�!�eOе��; �u-o9c�A��'�X*�H[����;w����ӯ�z::Lu<<�c��)�(ڨ8|���G��E�F�[,�v�K%O^K�bg��|�޼�,��5Q�����<%(L�!��/���$��X�9,t�8�����`��F�m���(�;=�YEnp�@�V1
��!�[����qf��wI�@12o?�j�D^�ߐ���6��l?2�SVs;�hJ�@�E��v_�++������?y�đ�\&t�;�{����.��P��sP��k�����V���m��g�dM�r�|C7���<�[%�A�09��;�~hp\m$��8~%H?�DY1���g�P��lޖ++0(����E̢�{e.U_��
���&'�.�����Evi�U�j��+?���g�����;:��V��?�ra�{Z*O7`��B��W2M	�u6�>�����+G��%�D�e�z��ß���g�[���,2i�e�tZ�|�����O�j �2�F��"/Mm,Dh�x�:��|a����󝿏�6}L#�&Y��ߐB�F�ɅKR�alȥ��5�G:7	�u�h�-�*����/[C�Y�-��/q*ޱ��$܇F�܇4��AtW��y_�Ic�0ՠT�� .ޥ�ek�T��O?������l��b���S*w��|s'�y̤Y��]jn�}-��r�?��AX���A������t״�p����5>1IX8�m��rʗ�)�ʍ�i�����b�F	#�5\��9�7�)�j;�8M|'A�6qa�_��P��}����;D>X�8 G밟����o����+ĕ�xx��#�cg�#{j8$:� ��Z��L+K�͙
K��Ñ��7������;O�Łh�n�3�,�N�/\�P��
���%&z�FQE}#]h����p�Ta-$q�S��`C-�\���w;� �Y8�<\Ƙ�Q4[D���_��� �ȦJO ���mbB�bC$v�C�e�Ĩ��~�	 Jb��0{ @���To�5a{-pL��4�f�1}rk/�Q�����l#�ڪ�8�h"KiU�%*ln�;J���`���B1�gD�e�;%A(�g����MrX'{� k��%�*'�S퀐=gљ?��̨�!Y�,[(K�v�;���_�ɬ��1��Cڣ9����$P�sM.�o`�磖��e���^�n|+�8��Rj��3����-��h��lo���A����9l;��Գ�C�f#e����lӐ�۳�&h:�{s��/bFޚ�������M�l�d��9A���G��wү� !�?[g�y��J�5�##�<$�&�o�(��R#=���~3$񌭗���G�3J��UiB�#�`��}ĸ>=�g2��н(@i���t���w������֕����|��TS3�F��lS|�z��/q6ؠփ��g=7��.��ʵb6.�UA���:}�Q��w�O:�uߴ$i�6���\�p;�� �]GP��z]r#�%�RVo�x��5���72O��A���}������f)^֗s�P�_�mF�{_DqO`�$G<��۱���O��D�2�C�<&�p�ivj.��b�"͓��X +���$�i��t[ہ�$�� �DQ�����>�%��Qp=Z�|Y����H��vIUB�����0
��` ��o��d��Ip���n�܏� ��P�E���S�U���fJ4Y�Ɉ�%�=����0���v�_T[��&��9�q���\��lE�
R��rw$���N��$=�T���H3�BV����\�ZD�P	����1k�Y��^�Թb�*x6
���F���j6}�[��c�+Y��&���+��0�YF4��R��zE�[���t���X�b�Y)���h��T�����*&�tڮ�z�ޱYq�W�]��I��#���/m�������ZwM�L�I1rt�[^>��CY�PHH�б|���q$/�к�"�TM��|�2/Kw&��T�c,�^ӈ���;��V�����GJ �����x��o̬F�H��v�#��`���5]C7�6�y���#cTx�FW�<�6��� �RN叅��@�p��0G�,�t�3�S�o@|��r�#}�֡�/���\��_B�	���tõ�jԛD�Z�k'�cc~(���م��klg�+�v!��*X@F��S\B�T��ͿW��"��X�o�go�ڲڟS?2g� -J�	 ϖ7�kF��U�?�E$��vt<�p[L5̝�J����P��H����p2xQ���t{@L�$�Oo*�/��;�f��D�,��e��5ݍČ��_9H�G���N�A�WxQ�zM�#~k����οC�Ӎ�w��!����U�qu��d��	&�n�L�3r��+�zZ/FJ S�bNG0��R����R����W�x�)<B8��������4�����w�Fӹ�{��4x�k�-*����0(�trt��?u���2sN|�߬��A�/7�ѥ�Q'D�+<��[�7�D|v�r��H���\�����eHu��9MRU�k��-B�4�t�qiڤ�J�c��	J�$܏
�_���1��pF�T�/[��J#oM�)�]���B�ˎRh�:K^��w�����'�cZ��&ש���~�*�$�q�c��v�W��ٰ@�z�ɤ��B�5��aK���Z�-�ڥcHa!�ɺ����h�I��X�%y��<�pߩi!?�|X�{���+��]m�D��ۈ q�����F'�gZ��<���3h�iJ��M�]__|Wg��f��3�T�������B%�����&�+<�wY�ڵJ�MA�İ3:s���Jz[�*>�^�ކ?BD�	-��XV�֓��K��<u�K���<��D��:�<<B!�p����ӌ�}���i5e��C���C	E�.ǫ��B[��=�[/@g��Y(?�ARN��#����+�\�۬�O�����ޫT�ȅ��8���)��!A���k��7P�����!�˔���R�W8U�zj#��PQ�Ȱӑ�q 7�HLG7޸���&l��W~4�������m���r����I���ў)�F�S�E��9�L�. e��S�Q�G���"�ҙoF��u��$>�� �>\�[����p���&�N;!hjK�����H�y��5�T�->|��)U�ɝ�7	 ^��0��-�UE��'nK^b�d�zN��)�h��g%�:�\���`6eV��i `�Rx�ug��|�5�pɴ74��L�R'��M���a�_ �c�Q~���� H'����9D�EQb.�M�E�����˵+�6��ht�{oyRr0�����H.Q��x_�"w]y tHfpA:�s�]�0a�%|�\����H�c��B��Zb�aT�k?WC��2p-R�F�H��Q/f�~5�>^	2-z����rsK5;���'+!�o�
�X���0��b1<�\�xx�@������AW^帊S��H����Pu�C1(�<ń> <>����?`�p����|��%��v�#Yi��J�4p�ey��_��<��j�&}t(��MHo\lA[|v��il�܂�¤an;�)��;�l�W��2�,h5�֛�z���iprSu��S�W��]�̤��բmJ�	85���SХ4n%� ������xzjV���Ijh/6������Tv����ʆ$���K�D,�3���@�KnJlS���k����p^+�֋��}�O���p���f�Z�߿�o�Yd�7���ph�[M�z��Gs���:�ͶIE���<^T��2�2�Ny�L�p7x�D�9�XX��+^�ƃ`�L����Ȏ��ֹ�����ԥ�����}��u�����$�jw��w�_!�<C���gj��U�m�ߐ��m���C�`�0�Ge��x}>Y�l��ɿ�U�b��*/���������jL����5<4��]u�mZ���)O�@�K�YD_����.�_�fv)�d�w�>9A�3M�,���2o��Q��Rl�hw#J� '�Xq����?�e|ߩ,.�*+,�j��/\Çߠ�hn�@0��#InDB}cS:`��$��B!�# gג{i�rh���16�^�s5�v���c��i��:<>H@�M�+_�]#�4`�;Hp�	�DY�._�Cv�m�/�j�ĹH�~����3���hx�6�/�.x�A��� �@�R�q���\_�D]/R��`��#+&�i��Fv�/���.��v.޾�����L���GM;���f�'�n،w��p�Z�x~������
z(L��t	�Wʝ�����瑹�8��Ҫ7���j�F��܃q������^
Xg��R3ف��Z��!Э�SdUI�_��0=��ԃ��/H�㶷p���޸h�U 0a��E�9���.�n櫷��D�h��7��m�<��aA!��z�rW@{��F�3�NXS��@��Ҋ�޹G�}�k��7�X���È����S�jG56��}T!�uma��[�Mđ��¤a3����Y\�5P��g鴭�
Bj�)Aj�:,I$w9��V�Z�_��z�e
1
��I)>�@CdS= �g�[�!9޼\fM2�ئLfu� �ƈQ��㽔���+���8�K�g�֟:� y��B�ѣ��J	8N�Q�X�������\��G�����'ț��hBD��%���Ys)�ze���G���C�R"3b�z|���;��'�Ʒ�)�h[�7�Z.�-=�5F���M"h���3�xj�`��D���`���\�FЫ*�)�
T��M����f���p���84r�S ��me'���n�w�߼���k����zR��P�4*#Du��P���]��
!i���F�Vd��3j}<O����FZoҗ/ �AmU�p�H�[���x�G��DD��xT�R��=z $�E�C�T�S�=M���h��XKl�C�ށV:@W�{���W>��
���)xq4�U�г�6�*n������~�Ɲ?&e�2l�*a�)I*B�=Vࠦ�gG��$SE�d]�|�D��9$,B�.QF��S'V����J�K�ꗦ���˗��/]��P��Nj�w�W��a��f�f������20q���K2 	�Js:d��x?�����\l%#�Wm�[v�i'5T�bN�'C��[G�-�4Lp}��+OI=��K���t�ڣ��@$Tb�a���iVf�.\ŨO&*aMJ�vN%�opC��i�R?��1apa�b�-yYoeAN�Q�,�D��inKN�{�@:U���饴�1q9(�����3B�8�5��:�@?�!S�H]tYD|��	g�T�	Ql���ڲ���n��W}���2��;ꃉ\��Z��O�Y���NԷ$R[:.���L��|���iپ�kϣL��I�[~���'DG?d��qm�����,�m�����=��d�q�D-��ުy���l���5�����IV/���� ܌vx��Ì�lu����wI����	�a���CB��0� �H{PL�$��~
��t.����G,�	1�k�LEA�	�Y/�63���J��xܭ�t@
\~���`�iӍ���)�Ph!ܮ�x�;@-��(�Y$�H�%.�CaY�ݝQ�\@�pk�����VŮܣ��~�C6��5XD6&�(t=�j3
��FC$�7)ˍ���[?��y�!���{�ĥ ؐ�u�E�B�����6"���y�����Y1�3uG
��pRL�ug	��������Y��4���v����O�r{�"���@��.����e-��I)� 54�T�N��'����ci�q,5���p�[�\-�=��2��z(%�Ԣ H7�����W��Fwu���F���X}ܫ��h��9̚v�� ��N�����!LYsO��5bD�C&�Ղ^�e�fX�����k!���i��7�<����G!��ָ$����D�r��D��G p��M|��]۰��gO:F��U��ꏠѩ6�U�g�'�#�濛I��>o�r��[�`����0����+��w��5�&[�&����g��71"/�e��R��\�Xx��\}7�
�Ii
M�
x/�7�\9	|�k�-����8�@ҳLVU���Z�m�$����Q� :�3��E0[�z2[�g�����+
��6�:�mџ@!��+�Z����<hS��Z�,(�,ٝ�:��v��,�D��bFe�c�~�|y4I�K J�0�e��{���?�a��il�`��o�\�L�����Bw��˘��� _��4���
2hzS���1�3�`�A�ԭ:��l؎����#��
�8(kb���i���0���@iT垿�&�����g���_M 
8)�c�XG��.�pBP���9�ߑ��s�%5΀�[�$�U��������>�hn�1�Jx{KG�"OM::/Q�M���H�O�q�63谿�Eg���M�+Z �l����8��q�}=��r�f-{O}4�-���qt�� �VS������?DRY�c6s�vl|����V�����{��6JzML�)�ޯ2�I��Rv����V�o� z&����\��i���$A-g�����-n�(�"�6�1~,gq٫�,O�.��������M]���t:�r�����!O47Wx�'ѫ��{?;�FN�4ɢ�Μ8[ε9^��5$y�w�O�����a �8?�Pc �n �(g�T`�P�+�:jS�uG��j�S7+
:�hU��oF7�@ڶ�e��9���S�3����g�d���/p�PV���&�Y��· s7�|o���7n��?�v�;v�s ��=6����{�yoT�n��fc҆$*�LM�
��r_���ԇ���㘲�}�b����8]�t��PB��':��W�r2�T��𠃣�Fo1�}��ƴ���\nD�[ce��*K>~*�֟XC�7̑�k���6C6)K�um��_����V����%	�`�$b,���
���hO�2�� x/�AR43�Kb�eF�M��M�J��*���t�H-�К6uj�^���P|���A���0��z��[�N�7��'�U_��r��^*B~)�	����FWH��{�
����>�3�I��Ñ>��MGl;��rN�#��Q_r���RQ��T'5Z0�@󄞼��	��ě�F��@%pZP�P[ʑ�
��K�Q��bEV:�!ߵ}����vf���-�K0��e��d���2�2����	{F��Ѽ�J�0:���������|����3��L^����e�(|�+�:��h��( NXҧZiBG��;�%��RE������a!�;�8%