��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�t�]m���moK�����.ER�����7��y����,���1����F��%o��yM������L���!Ra�D���6S�����ǡY�Uƿ��1�r� �� Ig��3Cݘ���m�)
s�k��B;ݗsΌ�iKys2���G��L������������ꕕ�,]D���`�ƀ����0�4�jK����K�i�nz!>������a �*��8� �Q?��g,ݟ�+����y���`�k����6�#��R�\eK8�P�Ȧ.�用�ҡ­����^���5���-���Hg�^&o�hz}��7ܕ��;����`���^��
w�5�2[`!�w�� +xv(�K����z�Vs�T�EwҌ$	��q�c;����jU���r�P��(�����o�r~ �c�8��r���o*�_�U��j1E��aAe}��
�
�L��V(�}�z񕶶���M���'#��sU��4Rf�.�46B���x�E˶W��FwR��w�ܳLJ-w�/tRrPr���"�x��R��8d3��e�p�E��-־�~9N�$Dr���A��1��|v�E��n�w��v�euQ.X�{�Y_q$U�Q�]�O�m�1+�81�6��E�+��j#͇P���BNg���ъ0�2��-��Д�E\���{��4���Z)�0��ԝ���v�@��
�!
M=!��%`�Y������Qֺ�H�@ٯ��.�+|�ډ"ɨYA��==�v�3)�����-Jw���h���MZK��$��<�ʧD��Ə����>$�[ʭ��ɷ�'v(��[�^ݲ���:!��z�g���_ltWY����ҟQ�>�iGn����n�	���s���4 	��&"<���A+����}PIJk�U ��m�4B�_�0����pm�x"��D��Vk�}
�Z1P�3���7>�]��v��X�2t>�zP��l�b���e�9"J@�MY�1�{+�.��1b1i5�0DVא�D9YM����P���	�=�W>��v}U,D߆�8w���Sdt��x�S�i�&���oܑs	V���*p���b_6+b�AZ��ͷ��cP�#9�����Mc����.��H�P��>:�h�6dЛ�ӱ��#�M����@����T��N��L����]rx�3%՛;�lv�j��sar�\��s�;˧��R����6�_E��t�Jw#��j5���~��$2 �j�0@�v�T-�!S�osV�Zn��`H<�x��lT$v����	�x��n�9�08B����\Kg�����k�Jnz]~>{&�bB�y�<��F���,	�Nk����~�U4��M�n�H������ŪC2�ׄ�t�����zPx��1���vh{R{�\��3F����<ɚ>p?��c�o6Ӎ��;�Z�?���rĬV�
rϚSeX=���W�PV�D��MD�/D�sNf�3�-Eߖf�tQ|R�1g|(��	E�!�<�(����ua�:�!<�崄w�S<��F8c�ё	K��t��Qi��O��!����a&����[�%H�A��@kɂ;<�	����;fˤ[k��ې1�!�݆J��Q>�2[���A����R11���ؐ�ۅ�v1�������+�1B��.�j:���:���L��}���9�>˯��ݽExS�k�-��%�aQj,(���\g���G;��hc�� �ޥI�\d����p;�T�K�-�n
F=�ٍ$�p�7�֡�g�l�Tu�Vn���w�CWvpZ�2o��5-w�O��d�(�D۶�<�dGJ�!��|����$�ƦJ��`�e���-	/����D"(F���M���~�g{d�R:`5+I�;��V�$��}�����D�@%�ş{���-/���$')�G�FiQD�(�B�i�&o���Ü.�Xjt��9.��,N��'���@��NNʪ*U��|L���U�Q𮥵��j'��P��������w��z�sX{,8�	T�C�D,*�"ˢ,/��p�VD}�,[�aރ�d��Gr��!�L��G��/��Vu�G+y�;�\���ɭ��W�˳���X�|<*k��HJ���e�Uh�_�����*n/'up��xٳ�khQ4>kZ�H�TL�v)WI�zjJ�U��u��Q��99�ؖ
���S7����pr����9��������6~#CK�a����d�@4d����,F�X4	��Ș
�j�n9������-�$������5dT��i;�0#�Y5���3%	V��gt��!��@�xf�z������	�x�+d�?=(z���2'��A���Z�/��'����Xw߅V��HN�Fv�B�Xb������vE�D�p��n��}�Q���s�l�O0ː���[�[l�U �Vi��f)�@�J �dv����`�i{� |��28h>Ｇ�����N�m�A��^R�@kuP�{���"S\=��qx�ƒU���]���j� ������F2�τ�ʹ��i��s��B��$���A���3���p�P���UDx���Zظ�{yf�yGΊ|C�x�gͳ22�q^U1�YC��5��-���<��ʏNq����rʤ�%��̵t/b�����E=��[��`�'e@Ô�O��$��ɮ��l9������_��<6���sE��t'��,E���:pqV[�~5��,-ȅ�T��_E���@閈V.K0a1).��8�?R �<߃�|�3(���g�F�h!JK�����_�ZE�ZZ��*�"A$gH;�6�a�5B���1��{`ht��H�c�q�Anv
&j���!-=U�<ߥ���wǹHR�2���\C��W.�uC�n-��ʥ&s�J�y�f���h-M�����j��2E��
����SJ5��`v�Q����4V��1��t��O� fN�\�FIDy�=��:�#����_�?л�v=iH�n�� �u>
�x�q}M&r�d�iC���$BAV1�h~q��C���3��g`ZY�$���o%=K�������f	"�9	u�!-]r y֘��|gyx���!�@�Y*t����〮�O�xl�fs�'��������2��r���oSΏߖ�S��TU�Q<�+��N]�NZM�m{�t�
��Q��c��~_����� &G#%���)��z�y�;��L����YN	��\C���T()ƀwO0��\h�K�L�' �=���v%�q-�*��}�DRp�y���`�SD[]�K���@����B�)�V������p��c���p`�����`�>*���^aty]{(�O-�k�*1��wu�Ah�.�������<o�YAf��#r�b�4k����)m���1������H�,"����f=��+�Zr?Fˬ�Zt���_��:V�m�E��h�����U�0&���VugNbv�}M�2�I%�ƺ_ae#�̬L8ҁS�}ӭ&Iz[�J���T�ѣ,�����kGі�DG� ���x�7�T 	A����f�,��ć#�����6�)��,���z���/U��$'M� s����K��[$;�_����O�<d#�vݜ���L�~���m2_��N<��*�X��%�����1Ju�����Me�J%l��B�)!��d/#�?��1��P5+8���W�)��4p*�؋�����{�0Z�	<ZAU	Y��Wd�䕻��`��=�{�������srZ�^� DL��r���/˲�����c!G���(>�a$ep���@9w0�%�9� ��� ��Y��8��Ud
rY�Il&�a=�)��t�ԣQI�	�~Y���8��KCP�/��6���>�^ū��Q|�A���U�)��F<���ú�>��gI�$����i�Ž�6_&- }�M��^���a��H�H���?���:��\#X	KM7!s?�J��J@q7l���Gedfնn�BRZ�Z����s���GɫY�-F��|520��Af���I�)�s���s�*���Sď�����֣ɫ��.�P�@���󉔿Wt[�  6N�P�����y�exl�D�P��l�(��H���Ї@�.��`x��Tk&�YX���Ï�T*`�+��i]�b��IՀ�P|���X��S�Z�2M��cis�(�3�6�.���= Umh�)�0��2`�Ȓ���j��TB�!��,#\�.��=�kY^j�h���	]��]���̣�u��k�ߜ�w�����V���A�[�?R	D��k>U�R�[|�l��~"Z��}|���1mó��C�>}O�8S���׭�ŉ��g���:L�MFv�����ҫ���f1�®�v��D����ڽv���XJ�9�<��u�����P0[��VG�Fٱ��YL�9D����[J�~�6u�C5�u�U{W�j~W��q\�,��+M�!��Le|�зK�ݓb� ��_�p��Z����b��cn� �W���Ŧ��k�iL���1�%L��l/j�!�����l_�saqw�CMs��x�.F���H6rP�E*H��6�^��/�IU"�b D�f�(S��\�O��X5�<�#�RRf���zz������얡ǈ�q0Q�mٯ/�G�}`0��;�~�0����N��*sv1�Y6_����U\�Q�U�A�$o�7��[��+��<D�&�C�9��� 5ho�ABۑ�n�}��-Z���K�K���-��s��R�_*	��GcP��0~~�Mjрxv��K��u ��j91 oE	�\���������yߍT�'gݛ����F���'?����u6�����f����M���i�`��`���ƶ�)X�EU\G��:m�@Dݲ�Z�7o���s�#޺�s(,ũ��%�ŉ�tpu�s�҇k�$|"�t�\hH5�$P���#�������R�q�rҊ.�;iD>@�	J5L0��z�K��_v�v��{o5}l����0M�b�����m|úa���A��ʛ�m:v	G�%4���ibof�	5���W귅f�?�ό��n��*�$�/P>��b]�����+B��D�퇽��t%�ҷ^]��bI�ak5���U���
B+7�;�Φ'4��o5�0��c#�4���7�"<It�����v1���ya(�  h $Y)��h�x]d���*V����G��m"t<��3��
%��^Q�0Q���܋G%}[,#��#�Y�Vԉ��l�-��V�����f"��Z�������]'��������+Z��a�㵋?��DAxH	��W�"�V���(!��$	_ʨ��۫�Ɯf���[�)��8Ua��}fME�?ՕRZy�i�uo�w��D�Hh��P�Z�A�ֽ=�q�+V�!\�$���O:�!��wcmDX._ՅV`qTŃI�^��%-$�,]|<3gV`TW��T7�C{��쫤����A�?=���D���&qPA#q�� F����d'�Z��OR-P4���������������$O��zV4��wo�x/2��A���K��7�f��՗����HH�a�����^�}+3V�^<�ܨ�1	b���;�Dr��0e�kݛ�@��Ϲi��/���8�Ԑ�g���ܼ��F��b�P3��+_�#Uw�K��*ԛ���y7�9g��	����HI���a��7�b��S��z�Jֳtl��q]f�č�vǱ�W���~Ƿ\Q�Y��~���w�֨y�{�V\��i%�>WcO�$,= L���aa�ڟ��i3��jIq�[���q8��ԗN����	�ۡ�^�!�μ4t"N�H>�Q�#����j��G�1�w\�����p2��v.8~t�:����W�Fq�)��vW��H��9�қ��^�n�h��ۜ{L{M�M2����BIy�=�*⣿��Y�c�����A�~�ܴ������� �þM�d�%d�X���cǮ�e��H����Z�j�r�C�����{�Q�������Ű�R_�w(��v�s��YMZ!±����Z������G��Z����I�}�^���M������:��tot[�һm�Alvۣ��F%T��U��g���gB����|��T����Z�����Cr�B�y��c�!�AB�<-��Yd!��EF1�-MR�E7�U�����8P��@-x�d5�|M=�y�N�@��=�Ž�؋*�D���'�4&��?<XGɁ�i�W[E�n����{=�N��W�Z��l��I�A�;$3Y���%k//��OP���X5��i4Fy�Jkk�/���rHlZQB]�C����>��%O�ym�Oz@�B��tt�yo�O�}���Q4-<,[ЀWbr�<�J����<�Zv}�$�i�_�n����+�!���T�mE�@�'9L_O��#)���z�|�8N�X�N�غ������!;3���'��2u� �Z��Y�[�r
��cG^��?Ї�NƷR�C�'�H�|HĿ�(3�%��:�K��^4���������������s|�P��;9Xױ2Ŝ�]��T�����r����(zFky�9{�s�5��r{���Ckp�1UoΤa�4��m̞�#�x�,���B���7�+��߇�F��tWC���	6^z��¯���P�����6֮|�]V-HD��5�Yo��Ƒ��]r@�����M��g�j�ݨM�����.�]����V�i˶濕�p���D�LWXp�|drF
��©S0X���b�:�|�ړY�
Wם�w����/��kx�?����Q�	�M���W}ZÅZ��E�qI�vRͥ���%�'EKÀ��� ��b����O�!;�'�FD�>�5��<�B�7w�p	:c�)1`ja�Ku���9Še���4^�C6B�$Y\�WX����ֶ��C%�
Ku�۝�PXs�������2��.�][0�Q��^=�&������
���������Ӑ��pŮsE(�gcX�ɬ+�����?�}O*Sj�	�ʯ��H�d�V�&]����#�S��hr�T8�6H��~���h�������2a��Z6��w'�EE F�u^d����R,������=h=�� �h���������y͋cO�40H�-��5
G·���!�g���Ø"�����,O8s�U����{v�ֵ�:�|G����t�f��ƌ;��@&��G�
T��5K��U(�����f����UA@�����f���B��&����?�����m�AfJ+�R��X��������H7��up`��	*>��s
k)��k��jK1�T*��y0+*]�Eg�-��]���.X�`�h�W���_��� �a�n*��hS�}T)ȍ	kW8� �as��w��K����Nc�ZS.��OTI����u�Z-��KZ��e��� ������}�'lpQ\����Dd�
�a��,vC�d� s�d>$���=�]O�Žz-�d$�lΩ���{��߃��a��7�I�=�H���fiov9]�.�.)�(���D
_+e�Ax���Х��MGӾ���?��׽�.y>�r�$kq-��"��m� �H�oR���1QO1"�r%���Ktݟ!��9�@�\q���x�R��"`�V�c�.���$<��er�0Y+1r��I!�&V�i�|]kiԉ�����P�Nv}�J�BQ/i�yD���!�-`�+G�s
�g`y�a������7��z�?��������Uu�d���E<���T3{w:L�A�*]�3�I�͒iI7�")�
%���{d�Ӥ�����]�C�A�D�a�3�$�J�m�B���i
��T�c�hM_�9�Q��]i4S��?�o�&��q�|Sṙ���0�%��3p��-�Je�B� ;���a$�3�J��C��NY��P�K��H��]�?�#З��.>g{0*.��?4���&%ǍCl\0���Қ*��G>E��&�.Z��u�����TL�9�ڭ\��z���֥����C�t?��DZx��>{ a'kv{@��e[���O����u[BxF�x4��ywV�!] <5� �
'����{,]V�具L��\xZ�N���� 1����~N��VJ�|�-Ik`��Ũ���Q]�f�5x��xcJ6E��i�U�r8d��uMK]�g��Ȑ*N��C�T��WE�.ZD&F���eY޿��&�?����2+�9�dD�ĬTUI�Bo�������/����p���g�pr��I��V��P�֥� P{��J�l
������Q-�(��Yٿ�|�=o�8��и����tj"����,�V[�Ç��C��#��g/�boE��L�h�'m{髯,@��2 ��< �{W"�Y�F�JUt|���) ݁m���Z�"�@�L��Ҵ�=�\+1�׼�*���ݱS.lyv����|����O)�#�]0�r�~��C@�Д8�"�<v�,�ȴr��ꂚ��x֤rm<SeEB��!��/�X).�S�I���YQ�%��XZ^'��\C��>��QIa|o�*���'N��ض������YW��o;�bz��@�����������H�sf�rH�co�_��똔й�W�$g���/��o���������� `�ö	Z���ú4xa��3��$�� ]������I@��� =�K-�K[N��oG��8r�4}�����f��`�v��L*E�X�����ul%�'sA>WL��$�I���a&�H��,��J�h	;�ʳ=�O�b���r��ݒ�cdA�9>�4�Pxhcz׋�M��,c�Z#�nM�����&�=�ݾ��(���4��c1��u���Ay�Z��>�8cy_��r���-r�+r�A ���j��|�m�ԏZ�P5��S<�K��vx�͘_Őtp��IiG�	cB���3���`E���4~j�̛�n��x�<�7�(n�@Î�ZSu%�`�#�Ը���MR�e�~)}NQ$H�{���������3�O)�GrOIU|.(3�b�|�9j,;�;���P��Oݷs6�U���!��&���'�~�Ǐ���!F_-��T��z��Q�FP���v�/��z�]�X�FAJ�������5�p���34�R���bS&��5l��'!�j��#��&-�0cɊ�@>Î�m��2`O�)��Q�<Ř�����B�q�3uFp3^"�a/��m��M�|�c��� ��k��}���:	�)'���!^�����u��bJ���{���r<Ѧ�;�<08���Yv��P�o�G��=��n�j�y�b��\Z_]K� �ٮM��<O��a�/��đW��� eE��H >���iH�MH�m *�� �l)Y�`��)�D_W�-2��i��dkRD����7�͚�?r�pt:Q�y�Y�8����	J]�3��f�`�?��J�
3��#��Q�����>�J�����GF��3A��������u2��j��br�ܬ�㸮s���T q{�}����X�x>NA�{B"$-/����4��`�J����ڻ.��b�ۙ��jSl����|-yx�<�L!'Z�cMc��uWF���1�������?f�bG8��
,a���
�Ƣs���d�RU�.�1�hy@P��B���b���Ii�ցG��n�9 �����eEIE���Gӂ���3Y��F��^ ��Q"�Go�X�	���,M:�:G4�37.����Ȧ{��(����Դt�ҡͣ��Gq�O��_q}8�*�g!q�z�
9[�P<j���D��G��}'���UkE�|�A���^��� ��!�ԡ�����[$U�����`j���ֶ����M���O^az/�ؗ[�'����#�-5u&:��B[mF/|Ҧ��V�lLKo�hv�Qf��p�Vr�+q��YaA>���Ƭ�]�b��$5H�e#"���:�}s��c���1��=!X��J�����д��s����b���co�x<�v��\���cI�����!�FŊw;����.��g�M,�*�B9�~����U��q!v�o~CE�ml��ske�`[Ѹa�3�����Z�InZ��% 9�>e/l�7�ʣf����%��Ҫ���QAp��w8����5~8?�N��7 �#��x׆E
H��
q�*e���#��N s�̬�y�]�.�w}yt�YਬQ��T3j�H!!%B'8'�cہ�1ۺJ�u!��uy]_��]B� ȇ�э9G#�7Ίks��X�Ya݄sF�Zo��
(���o�n�r���X���E�wD����:C�ӈ*0�pY�z*L@%�k�#nOe.ڷ�H�-�����Կ�'�M��$�`�@���/��r	8,���Tk{9<�N)@��0��hSlO�������+�e�m2���}1?�j
���a)wB%��5t��7:�ҭJ~�V��Rol�w�nN���˟>Ր�cI�&I��c��Yu�r�(�fG��h���%�`���+�(�mҿ���®̊S�|�G{�ʒc�F��"���RJf���ϩK����0��l�+İT
"ɹQ<�Q� T!MX#rK��>��d�A?�����:��D��\ä�)2y�&CY�v,�M�����>[�SK��2���9��1��w��a&u�ॎ�um��m�`����e+7Ӛ���0��^0:F�ձ.�t~�:c3�b]
p�5!,�9�Ƃ��V���� ��#�/��Sܷqc<�n��
V�g�h;�H���7w:�'fB(i�t����\3�.%9��z�ٷF�X�)�`<Y�5��P�k�y���௔�v[��\їi���­�\�%4:pRĥ�_��6u��w]ȽRW�(v��B�M$���d�"��5uy�f��;$�,�p��Կx���C;