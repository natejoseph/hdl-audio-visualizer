��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�v�-Q����n'�)Q��Yo��a5IH7Ul�ޡ�ѤK���Gu�@�b�)�}?Q9.d#�-8N��6e�NKJ'f�,$�-*1!�w$'�ݬ������i����Ջ��2�z�m�#��o�*�S5coD��<���m��`A[�{|����d����#g�k$�C��<���+BI�]Ӫd�t34�&b@�G��{9@����}�MF��u.*Jm����E�2�v��"��-*���j�w�>���I�abM͑�0L���>�Ψ���z����^c}��1�vĥM�d��QIr?�I���["@�e���w'T����������<�Z�|�eh$��@]��	 �9��h�őa&X�F�����+H�¬����p�{�XZ��ǯ���usZD\�_�Rg���_g8�af�Ń'Oz`�]�CXRx��H��t$ߑ�J�����o�M��BX�]��ۏ�ײ߲^�]�����z��y�c ��T��ԦJ;%�(3�A[�R��*=3��q���o�ϽA%��Кr���h�EQ&Nu�w	��B��x��?��:[G{$oe6��n�,P�x�L�,��HW��Xc.:�U�):�K����V�
�q�ѩH��tL��
I�5�LR��E���B,8�ۭ��J��e�n����Fz�`Ց��g��s���eӍ5j��a	@k-����Rf�c[cإ|K��z�d��nD�B��	�c��xy�[� H��n	3;��Sv���Ol���a.��������n��Q�(��Y����?V�=��]���դ!��y��q'I�}�w�8��4��YI�Ĭ�:m#�\ˌ���M��=�r���ѭO�
 J9��2���A&�
����TO0��E�$撰(�JYXA�� 0/W��I�A��Q��F�/���;�J^�=���4����ػ~�RÞ5U#����Qc��[d	A�F{��o~��\���Rڌ��$��nd�+�8�<�$'EWu��d��݄�%)�a���I/�<}���&q���# �J����o���2���t8�cф���g���Al�R`�2�Z�R��[^��9�H�������dŮ���6�TQ�4=���*��g4��!�"���������У����i���8�[�n���@�5h|M*9MHlsؒmϙlaI&�X�I�h586��Q�@'�?������^���N����dk0��S|�#˅6԰�B֚���2�yE/b��?���]V�ߍ`���C��:u�T�0�(U��JG|.� �T8od�5G��e� ;�˅3�=I�sD(5_���8t*|�x�����\��i����΁���	*��C�����B�|8���%�Nh$��[7�Xp���uo3�j�xIƼ���m�<��v8��C���D���N��-�o��n	D.���MĂ7RCx	��P?��vi�j�G�v|��j����h_���@������1��g�a���а'��ď�A��v3R���[�>r�h/8�^�A�t��S���Lr�e�4"���c3�1�j�?��\��jpqoH�]^)����r�Ob�	'H�\�\j���=^H�otF�ő:�.�WV���|1��%���O��]�l��nCH02͏�`��7P���,��u3�s�:�� q�v��Dm��GЯ5	 S��g�i��}�2�9S+V\����*�����ؤ�{[$�D�}Z�e��(�S�T1��ȧ~lS�B��h D�Wٝ�*͞�k��"=�
�ѳWS��cxU�2�6�Vp��9��{XMI`N���E�b�ǒ�	y|ǿ��*��Q7D����e��Y'ö��F����m�y��HQ].5y�`�'��ܦ\����-A��L���B�5�9o��`�oKO�(�N齟�a�I���
9�e��z�_�Th�.ʗbƬ�f�l���v�)JT&����Ç��&^O�0QNɒ�~�5��������^���6O/`����3ypPޖ�i+�oP�(͏�hș���9�k=�n5s����Z?2DG���1Ȭ�&ѷm�%�t�6���GzR�e�N^�ҏG��#�SbiH)���Kf&�}��M�`�;`ϼ�={0�����@$�Xz���p?�`(Z�R��7���؋��`SS�R!�����<R��[C�z(㿬�Ԁ��)�
�R�g_E��F?����8X���Eh_�@�|��^(ua�t��� ���7:pZ9_d�GU*�\9���u����I[�H{!�ҋ��7@����u�(Z���׆�u�c�>c �(�/�8K_��V5򏒥�˾8�7��pҨ*�O
q?�qb	���\��˰��H��f�L��6�ˣ+R���v��һ���|�]��h~Nq����p�ƒ�LZ�NzT/;w�-DAL�C��YF�l�m��%�2�T� QaKCsdt�]�A�#=��uЄ����Ո�+�m��{��B�wzq���I�PZm2���Rd������u)���7�uƝ�q�ƨ���l����H��\	���+���d�Bh)�T���l���v�t	ɮB����gMG��oV��T>w)����K�:�O����zX��*���<���-�Zn�n]U��zt��{�/|y�7�+� ����7�b#�u�e,�?3����mesn"/kҦ�4����r����.��O�8�IL�!�앭WY����$Ϫ����Q[��H�����R[#�,�jVh�޳�#_��0�A�	
E��&P.U���2��p�,K�P�.%��8���1-��nNԶ�Ya�Ս[��h,E�y:h��^l�z����1�n݊�混Ɂs��Y�����{�~χ��F��� �濽v�4��1m���R"�)<s�1��F�,�[�c�(J����Kb�9�]��7�g;��)&2Br&~F�a�W&9�i��M�UZ�e�
 �O�,�j���5����k�z[�5������ֶ�����>*Kb�ܛM�LT��rڡ�w��B�aI���R���9^h�x����g)���x��Ij@�J�;���d�l��J[��4_���yh[�*�CcH���&/�@C��A����k�'f�9&K�}��L�<�t	�����5+"
X�[�#M`3�y~f�� R!��o]a����9:���s�S�g�o켈��7w�
��,гzq����q��P
�ߡ��c?�[{��Ů�it3�4i���&!�����E�gv�6[f�� %��j[EpF�&⬞�N�r�/l�Co�H@ֶ��NTu�M��z>��Y�w 7��8��H>���ˌ�ΰ?'`�k����3�N��X��89�ߔ|U#��Ң��m�"9f��qS�����-�4�>�%Ȃܔ%cE�VYi����[�(�~5~�O1��%Y{�wq��˃�z.l���y�B��`�L5j�/��V)�����b�$7�p�-e.f�v걙�u�-���8�<<pfo���dk٣��'�7o��)Kz`�DeOs߳HT��K�$������7'kT��)�=�L���'i�FK!�Qef������O5s�54w4��1��`gG� �l�pAێ��7�J��%n`}���k�+E��>	AӐ:"��z�IW3�Qkc	�n�t����T��4h(���b:s�R�Ш	�+Ag� ��Rm�Q�A�DC=���,)c{�����(/�RO8Y�Sޭ0��d z^�#����r"���&O�Q�1�L��u(4�/72]�$�'4�D�
���X��rov� ����;Y	iH�<���^���(>��Lm'��FC���>|�f�{h��RON(�\fI\_�>THF��a�c��;>��}���~V|>�y�l�}�#��yJ��41y��5VZ&@һ��x$q�������4�h��;�J�%�v��\��삉���Vb=�E�Q- U�������5���_�Vr�@�F�o���`w���Wa��̟���gt��'e���8wܽ��l�^�'�e8���r�h~�`�9���C
vrFTձ�AH�I���(�A{2ua�#r7��� �ެ\8����E���-�v�1ϵ_��#s�*�[��h&d��A����G�r�Gͱ��&|��d=G��� 0�W���"Dc^��.�7�"���-^a��P=H�H�uݙ�m���h(����TCN�0��^vgi��*�1VSn'���	t��f�I��sð<�EX3s�O�����VEB�y�+�K�E����$.���s���0ۤ[�1-��y`�/V���&�{�;�B��=��S�k}�b����v�Wi�ĨU����sR1E���}&�	fF��J�E���n�T(��:���9$a������V3qi|i�b+�� 싢MD����Rtx1�$w����C|vZ�a�b.�P��zɭ(ɜ����ZA����T�'��E)��{!�<N�0������4���?��UeQ���NW����>��.��J�9$�wN��5���Q�I������,���v�=��4��
�0D't��NX�PK��c��\�