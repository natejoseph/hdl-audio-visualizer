��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C;�t!�𲎊�$��N�ye��B�Ep���ĸ@����I��F��NG��Ӊs���oaxɑ����7pl�^�ǿ_�P�W��98�N�����+s;��:�Q�,fq�E%ҷsM�Y�`1`�էOk2Lo��{+[����Wy��a]{H�)$��ļ]^��+��<�eh���Fȝ�^�M�HX/J�M����E���)m���C8"*R�"GZX���mNz/��=���`��qc�%�1���c�W��D��)�&�G�@v�oC�ddƱ ��:&�)�ԊG�e���/5=`w8��A�#�-2�	���`Fb������ w3�);mXr1�o?��o�j3<�n�m_���E5�q�7I�U �3CY0+�������
�f�|��O�����uFm�k�@Y�A�䃒��	�7��WJ�؇��S�{�/jy�� 6��U�U1V��!����Ŭ��-Va;Qy(�0=$�	ݤ�a���-��	B�z�ᯫ�}O��F�A7�8�.����lU_��B�ʞ|���9� o�:݄��?_o��Ѱ;؎�Vl��qA��>���9v���Eq��;��/ʵW6-��t׽��e~�w�d(��p���$=E����f�����&c
X!j`����w�2����V6N���J�a�ҥz�����:����Է@�nv������ǹS6�41�	�l|e���>�n���,��ܕc��Hz5i��+�yۺ2�iT��#-7�R#)��6uWg��·����dn���˓Z4I�?#aup�_����M$�l����ۺ�-�C↧��`)��_�Ҍ}���1V������9���9�� �'��#���Qd%x5�a�sgD�m$Ո�|��z�?�.ﴯ�FN@u�ڪ���q�:q���D�o�K��[�Z�T�lf���4�g�mQ�rWy9�R-����*���]62�� K�����:�*�<aL^5�8}n�$�vq�+���7ڼ�{�|v&@�)��I������]½fCj�O'�K�^�$��g�p��ፔ����J>m��k�e��O�+b�6۬�ܣ�PU�v��sʗ7����{F;Cfuso�Y���hY��`����N�����m�	��l���oS����������,�g`S#1N�B$�o�'�\���˪��?�%K��EȢ�c�J�5���!�<Bo��|Z:�VyRe��6��a�b���,B��qt~��k��e��&ǲ��m�˲23 x8�@w:&X��a��+'�N�׆��5���"�:Z4��>���@b z`6�Na��,F����C;D|/7:6����y����l�<��0����A�W���VBݜ/�-`�x��!��.�-�=�Om��h2M��j��,	��(CίU &������z��S2�b�B��Jo񻪽�A�N�>>�{�*�R0w��Y�s�{�s�fs�
�ҝǉ�nEz����ϡ����-\�N�zH ����zȎ�й,�<ЋM�W4Pң�k2JN�#{̂�V���Z��
���E<h����Ƚ[����z(94'^+�3���G�?<��#�$��/���;�����Q72ZF������6�,��1�p�JH:���1������Y����C$��H��b��h�|�����w{�O}vMJk��\ME?�榵:c�]�o��J��9K�.�D��Ѣ���_e��{:�d�(��%]����vF�-n%�>�e$L��+���œ��vԆ"}��7�0�|���InL{{�	H��R��oZe�T�D~Y����;�[��v��hteT�Y'�=�o��|!{x�&�s`�Ԍ7A��o��ɩ�v�����ФD�:*`�H�����K߇?\�U�����52M��:���t�����-��l��b�/i~��A�� ��-H��ݧ��ư�=�Y�@���&tM|�@�/|�\��,��eG��|�P�b���\���e�C��E��]-�r���4�'�6�`z��	h��Q��lQ���f��B\ �K�5~��d�/��ԥH�'d����C�{�ׁ=�/���L�͢*�?����R�s��h��c�e�޻++R�6���s�D�FRVP�4~ӷi��jr����9�}�j�U�H9�몯V�����j��6�������3F�3=�&�U8��|U)S�9
���n�`�!$��8q�pXΠy��թ�VA �`����繣���~�~��?�]\C5_𫬲�i��\�td���.u�q(��M��e�B&�!� �,9֒��#K�-Vr�ʱtXq���bo������G�:N�9���1$����{QI>z�H�����߄d�74~�=j"j�]�1u�Q��0����*z`df���1��K+\k��uBnZ�M$��r�;�7փpB.���V�W�X����;a��aq ɇw�>=D.�i���1[�W�ՙw@Ew Icب%����IdI��Fx���#gs)up����M���H��;#%�[ߋ^�}�y��R=�7�#�L㶫�왼��lJh�Ӄ\`�n�p"%��7R�*��ԡ�͍;�OSx0^6A��nb�^�5\�ɗw1�c/@�+��{�ĵ`�����W�լo/6����ϜJ�3�����[���IH��ok�й�m� ��Ag��m`�3|j�^^>-�CʃϜ��u[�4�֪ISS�����ʵ�����,ssM�x������%x�J^�8�z�
�堇��@n��Ne�W��M~B$$�ƭ��nnPn� ،za�#�tl�ez�Ș�i��Ж�~#.��xHXKV>v<�bj�u�e�C+8%�vb5�kv��nĿ��
�}*�bb�F~�%���V']��0J՜y�����5aM���G�p&M#��y��{C'pa�TΥ`��jC[{�Y�ʟ�яJ���2	���k��2�ao�(ġ�z�}�/�������A��U3df1�g.t���V�{)���l0�����!?��tM����n�����?��-J�|�3p�*1��#��
$��i��m	�1��0�I~�}˟���Z�����'�9 �c.m�jE>#D�����bZ�9i5P׽�`)� rD<+\2"�iWu��8Z8�T���ɝ�z�˾���4�S���<W��A��d���Ky߭o����~}q��֢��&��I�7P�M��hi���\a��Q�q�N����2&�ҧ�w�]A?OM�?��ET�մ�:?C��u1 <�

ٶ�69�DXc|�{۶��J@��9�@x5e��>jh~`y����UB�V�&3�y7)�{de89��K=�5�4q�cH��g�����:np�#��h�����Y����(h���M�x�3����!T.-����˙���)�^�Hן�ވ�|�A�G�ӏd��V���G���;h7�v
��h7���?�(nB�lF5Ն���+�,����'���:��{�u������/["���az
�w���_��U��4r�J"�c���t��v��&�(v�\=���M��a��a�\����M�~잏b�$�|�x4�W=c;�)"�v0m�~��2I��b��gIh����<z����aO�`��kW�8�PԘڔ��]��Z�g�J�E�D��r���~�F�y6A]��5E��3v(�Z��cJH�a��p�}5z�����#�`��3�΢{g&`����6�ôJ�s��&��>M�\MӀy���M�ᓽ���L�����yQ�	Q����h,�`4Ƈ�m�c�U���[ oʱ���,/ ?&F�NY2PZ��%�;���&wv�I�v#����T���J�Tm�\�3�g�H��du�^*�T�Ƚ�`��y���i듿��o�':��r�4' ��я�w>������bؐ�^8{��4�y�N=�G�%��e�~U�j}��������N�\��?&���� %W<z~�ڐ��V�F	�ѐ$VBF~����'#�飡M��eF[>?�@�EOFM)֣_W��5�"SH��9����q�5���P�վm�h;�&�R[߀_�<H�e�����bk���?w;Յ (J�M��m�)m$J�5:+Q'�:���B��"pUz�}V�R��-����EL[�D��b�O4�G�`BA*�᪆�w����.5-�g&�"5���M�\'��U�����{��It��&-�̡�˽�Mv�Pܘ����ڽ��qs���f�C�����i�B�e�cˣ?!5�����"�;��Fj�����*�f�Y݈l�X������"!���y�F8Io;�y1n���x�lb�"��F~�Xz����Φ'�GY8E`W��f�NY�5ߜ#d�WԯO���;j������;L�n��1���0Q8���5��	�D�.ƃ2�@�$&���R��:��2��l�d	�Q|O:��d}{A�$5�͜2$�����3���ѷ"�R���3���Jf묨^�ş�L��ղ�t/J�<���xf&pb](�Oߚ��t�XO�t�	���8c�HF��]�����1�����U�o�C�f�ֱ���Qf�g���{����r�l�pw�n���q�����Np���3oW��Z㭇]{�o�ق��Ǫ����>�ղ�z^q˧�?��g�}7�)�֯��ܓE,�<�a�8�� :�N���
��eۑ&�:C_x�-�a�9s۔ٟt;��{���y.H�5:�4�=#i�	��p�Vg�4�?]k�2:�������6O�k[�'�
a�;-)�O��{����B���1�z��In��e &�BX���,o4���µ�p�h&`��`;'��Pw�F"�;yj {.�6���L���3B��S��A�ٵ4ރ�A�a�ķ:m'�][ �����Aq��_��q9^1�ME!Q�����V��&���'T��ڣ�2��������J�,bO�fG~�撏}�������bP���� �4Q>�g��B�E�x�0���3(���H=�Oޜ�>6O`x��z��f��y� �ߘP��vc9�����s5X�c�2 ��D��(/��T�m�9�MM ��ol7�eq�T��*�Z�����Um<Mi���-�s[Yy�DlŒ��e�唊���ћR�e|�Y+=�� ݗ��>֪�e����Gۑr�ʚ���h?��1_�T�y��%#��D��Tr���l}\蘒nС�[�v���τ�iE#d�Y\��k\�����m�,�r�{��]���d3"a��Ϟ?iR���j��� �~���CiV��F'q6�_�_3O�3"��[��d��_��b��pCuF�z��a�B֣ϊ�6Ӳ0��:�z�ARiK��hH�������O"]p*���P�>��zuD��7�\=2:�)���~�^Z>`ʔ�z�#B�2����ا����M�i�G�di���ڧ��mVG"UBp���u�X��l]A\O{�o7Su����<u. ����?�WM�(xM"C��KE(_��nfN���T4(�Z�!���(�0�D/�i���%�4&q=���G2.u��Y��]�"�Tb����!f��ʏ�+�;�>П����t'�?�ק���o_<'�g�K)����4�j��pR�mj��E��C(tp=nK���ۉe��Y߳�MXXݗ�u��4l(Jb(���愸h��_U��j��7~3A*8���;7@c�4<��p
�::`š'�Ub�A��V�$�\ik���Ĺ����m�&�I�S����Udeq/arVjW��
�w~�P�j�μ���5�������&X��p'��`Ag���>��c��ٹ�B��'b����\���'�u�GA�=�X��ۄ��9#\����_���h��eu�=�ǿV��G�%	ɒN(k����d��B������n�K]�\|�����ϫQ�6a�o[vF�k���ok��7*S��ۧ�gyd���}�(���כuf�/X�7�2"�C�X�$I��5(/�b�C�XIv
���׻ϓ������nTN�R!_���@7�uN�������� )�N�
��'=�����x2 8w�8of��y�n��mR�l�@�<K�SI	I���<)L	}[P�C�gn��5�#����a���>�}��c��ά���|#X�nD_0O73�	e�4Q夶�ڟ쫛�by���k��+��RЮ���A8�J�bN��0IDn� ��I�rHr���K5xY�0�Ⱥ��.�a��CR�Z�l�9)ټ�ޚ ��Gc�����ӖgI���ڤ���.A�]J �3 �$)G�q~!k<���AE��tt�κ�bn�#iK���MX�
 )$�������w@=��.��<�� �dE�YCh�O�.1{�4��m�; 4��𰐽�Q;���qTv"��o�����R�E:���wy��Ϲ�U΄�$/~����sC�ݤVTk�� ��k&&�yq�}�+���I
�^5�Ѫ�9�p�3r+�����%������*��8Y��hb��WuS�J[�W�S��#ȥYC�=����Oч�.���I�����&��M�Ch��;�?)�2��.���S?����/k��7�ݘ8^q� 1i���Qq:��\叻(���0�P`8$Q�G��z�A�r(�n
��¾�PW5�7�w�F�P�?8�7xK��S�9���/S\;-�RG���hE�1f��
���uxu��,c��[J
�U7�Q�<(�y.a��t3K���=�����9�
�F|��>2+#¦���ds�H������g�s�?�>��ߤ�b�
��3�Ұ��F=�z*��Ͳ{�/ğ\��[_!��[!�Ԇb�]B�\��?fsu��Tvf���s�n���s����j����s9��ŨrK`L�}���LS���%<��R�j�6q�\���`����&���j9���/�rP=xpY�*ɝ��Y�Yu��S�sn��Y���rn��=M����O%�
{�ꗾ��i�ˑ�8�g��K��7Z[O���X)���t�ذ��}&�&���m]�r�S�򦀘�H�=�u�����.l�s�Z�d*�9k���I�$��$v�0�!���S��;�N�bzm��(�<�����I
+Zs�
:�6�˾*�[�a�KqE��K�ޞrL$��|ˋ��/��]Ѝ�ax�k;�`�u��<�ݖ���w�J��# �_g�~Z'O�\|b MK2�چKMOi���%fzA&�_�נ�:�N
�b��U�V��l��,���ED(r�T�x��{��9���lǊ��R
n%�1�g�j�R4h\\s�K��+��g�yAS?"�6�}`Y�B�_ܱy��]���]�&��ܚ$K~D8_���ю��r�w	�> �"��Js�����9��V�4*#�2���� ��7z:��
@�����ٛ��������H�@��vIg���[t�U>�P1
�&�iŞaG'��lx����4�5�� ���(W��u@'�޿%mm��!������Lո(K5!�LE���U� �\�I̿��`�������|�'�(Y�����ŷ�O�uw͚���*Z�e�z���^*�(ET�*-54�����"�n��n��:���2fҚ�lc�T���ɪ�s �`�8�sl=���B;���qM7S�2�@I��� ƾ8T�R���a�w4�
Q��U���#ˋN��������b	�g�u��
E�
o�F%�A�K���!��j�At��G�=�)��O�ӮCJ�8�z(N�8|N���ĳ��v�z���يCh��`����������Kq!8����^�{��S�e�S��8I�c܊��1���J�e�����sq�f3�.ڟ����kϕ�{II�WoV���~�s��_�4���5]���I��q$K��[�u�)"�I����/#�A��3c����ht��؇U������K�;M	���y\�W�N�㨍�C���wE�J��7����^��7