��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�ɬMn��@\��NΉ�+!��?zIQ�* �G��ϑ9�'��;R�� 0����.�<7���C-,d��P���M�	����y,}��Ϟ�2�L˻h�-*N�)�����xM�ꫣ�,�E]I����C� 2��E7]�^Dd ������y#��ÆK�s�%ڗE�Ż0�{_�-7f׫%i�𶋹M�SJ�d� �lȃ�5 �h}�르�.*���?���?o.�
:���ZD�,0�X�+�Q	o����?���8�ӌ0�S�9��C���(�,��d7^ZwFZ��=�<�"��OL���]��7pX#����:����l���_��g�)����J��s�ex[����h�S�������:�E�K;k��z:J�;���f}LQ(�C6(������R������&��	����8����p`9x���C��"O�
3U(��w�p��2�?n5��q-H�E����[%F5�����C	]�9�6N�qh�I�����;�ؠ�6����X���4�n��*@�F:�#r�hw�m)N��%����FCX��l2�{|��o�����Lx��T��$�}#�\��@a�0��[�-*,��L:���"�n�"`��?ܬ��8�넀u9ލ#c��Rqf�h~� ���~��q�~`o�?���3ݽx16>E`}��׹�F�L��)�TW��q
ҲKE��D�v�$-[���R��(��ćd�1%�@���T;(��7�1sz�;��{M��V8��ݛ �l��t�O���m�����YY�{�Q2�z���3���������p�*Y5P�΋��u���d�gm&oj�8,�I�V,�Kv������;!�J9�#,fɍ]H�3�:ß[�=���x�%y��=�H��f���=����HZ�E}�1֝=[�(܄���|l��<Jw�/�+�$�j��u?/��ٸ��������0uA7	sa�1���&�\�W�<��-��W�<�I)��`�`sx
��#f����4�س-ԪϺ��V����S���AD�|W|�x�yR�,DQ4*�q|'�J��KȺ�_����JRvl��LR�����'�:�N-]e�LWzGx�g����4�@��]%��k�6!T��s�M�w��eY��a�o|�!-�TW]�pG�4��[t�C~�?�ӘJL��������%�P�zr�Z�:͎0�#�����:g����{�?�E�b�X)����F3��<�M�Η¥�X%Z�d�|6�ۓ�@A���]Otmv��j��+��j���|h���dx�T@uB��U� �S��r3~>��I��$a̅���s�:��%��˹�g���A����Q��KMұ���^H�`q���U�.-�?g��~V+�S���������)h��G�賸�9��v���260�^}rI�����\?�x,PGt��q����Ø�88�P\��
�F>r]el��.�ֶO�>�$�$�w�ZS̆�������i0�����RD�O�ޟ��-��]�����>A�w�Ыa|���Z�՗�Ѐ�QEW��5� ����P��]�S1�-��v�J�t
D��	��<8)���$Ջ�h��j*���A�@6K�7�jw�@�l��9���sŨ�-Y(ڈb�)��,J���ݥ~L�k� 4Z�(t����&�r�sE$��qF���y�o��y����a��G�Ĭ>:߸��,_w^�@��)c�6�A!T���c��$w��P�Wl�8��C��<`t �ڣgT�xd�uj���^R9Wơ�#]}��K�mY�B�y�e�8�.���j=��E2�q|_�O�X����E��U�]�*��Z`6otHŶRh�i�� �b�`��>���?�9���$����ů���5��J?~�8��9p�Vۨ&c���1U
��#nx��ӆ0�	2�E"!��II�xp	����~���,�:�H��N$�T���h4�a�W{�X�b^��oC�ȸ]�S�m���寂B��� ���(v�_�4�����	��f�ŝ�:9
�{��D�ʉ)������/)�G���W��y��^Z�P]v�
M��k�������>�m�&����V�-������+B(Ղ����6��20��-��t���Ϙ�I�_��n�"����z��,v2�^��9_&:ʮ�;�e�LI��U ~Jp���f66EŰ1_���̕ϸ��m�t�x]��C+cT�B^i�xPU��|V6���,�>�铹�wTv>]\��!��#��ʾSR0��9��U]#"�����_�+��u����3����a!t�z��� �`�IG\X?�{J!y��K�zl�g�J����r�ij����7��#&�)
ˑ�����X�Q[���b��/�$]���^mo���_=F0V}q
�	��醦l��{co� iӘ�i����$�YW��,�2B�b@S&]3$z�ڜ�"��Iw,_l������2�9��A}s��_���r_��t���c~���H�7^a�6�DQ��L�ș�] �6\F��,��_*�rr��	�6h�?K��jN�L���OzqU���\�@6A��ѹ�[�rw�:��ܹX�eUQch�h�x�;�ِiWW>����k��aK���E��'�~�i�V�n�[��N�7�;5���w_W5E6�(��Y�����,S��)��|OTz4�y��C#t8��	��d+����_.K���0��j�>��/op( CF(N���3"�7���g�dg ����V�b �j�lɒ/���_��*J������ļ����{�P�o�*Uz@���PV�Bi�LRa�I�1ڏ��WS9^mm��޽��&�r����MM*g�����2����Bwβ°�����k�W��Q"��_�"H�L��NV�(�7b��+�
�)�n̴�*���Ŗ�~���<���b�C�N��s�lx��7�5��Dq�2�#�IBM��9��Ɯ��<�=j�m�$u��^5�&yrm�J� !g�頔Eޛ($�TG@lj�-��M!*�y���?��C~����	#h@���e�!H��K;�����K�j�X>zW-A��e �i�W΅��q�>�#(�����WYԯZ�W�2<�:R�ыe��4+FiG #�	�5�i
8<�H�}�zcHui��R��|�\���d��`L\�]��Q��z�=@K�4�>֚�lk��h�����"&����)`j�
�[\�F�{��h�����Cr���H�O�����H�b�1�%=M�ldZ�F�~J�m����;�n?>�MS6c=D���^݌K����J>B���D����|zѯ�����G��2.yŒ0�ʹdס;���~-v��;���R�jW��L_�y&�W�>�#���̧��W�$�{2#ˋm��»�T<*�J��0v��n*�Q-f�ȿ���ڟ3=�R�,�ʁ8ñX�TdIE���u��i���07��5�F|!,�B�O*�%�F�'�~�z2�?�J`''v��݄�����+U�I%�e�u�&�(c�!,��+�N<=K��P~e�Ь:���9J���E��Ank���)��˰I��R�f{Z��|�L\���0}�aP�AL�Ȱ��Y��G��+��U��Y��Eq �<Ȁ|���
�gG��>Y�^�Pź_-Yr"�hW2-�C�	�9`���V5&���|�{�g:r
�Yz�*D����_��JJ��+x���E��>
TR��GR�_�2��9E�a�t*���.��-5�~5�v�R����%��'8��2J�Aw����q\?P^RMH<��-�#�&��t�,�6���B
��:K��Bq�z����(د�^�Nh��
��>�'�{T��}���#ss#����QT�Ѿz�ex5�R��֏��C=&�l�??�v�P搂�������=B�Y���'FL��\�y�K�=���!������k_�<�����a�ů��������M���G�O�ߝ�=���Cl��]g78m�D7�0i�ʄ�/C��:L���EQ$����l����ĭvխ+E����ݷ*�|�
�>�!Z��P�K�ô�ڑUWF\������E�*r�qГ�i�=�P ��`#Qj4X�7�X���O��2ˡ&o�����|����<PU2,Q �2"�P�_�h$���+E�]n9���Ǫ�x�T"�0�k�#�s��,T�"�h��Ie�.���z�4b��s��7�����e��!��=\��]������q%v^�j�%J��d#� y��&MIn�;*�]Lb3�ݧɩqh�j�W��_��J7�m�ͺ�f���Ѻ�h >�~���3��T�ѫn�A�Zj�p��Qtz-j\����iJ�6C;�&A�km/� �x�KM�3,��b�_�^p��q3_�I29�ں�J���gme���ת/[�B���װ�����[_��I�=�#l�
Mi3� �;9�DO����$/�":��e���I��+o~��L75�(d�2?[n?oWQ���.���Ԙ��&`yed9�Ƒ���S������~ԉڹlOM��;+*Q�y�
�끃_ bܚM�ϭ���^�R2��f����ܭ�m�0�i��~�NN}����_Mv_�NF�c��V�3��/J�G2b&ذB�W����D`b��xRP��i��j��3����<Jf�	4���.P�Ն �Y���:�q�#-ԝ��a���QQp����T)��`�S^��"��k\QUh;�'|^����`���6,�G#~�7�eg�V)}��H{���d�x�����VtzSom��tڛadء ʾ/��1i���tL�Y���x�����rٜѳ��1;#�dֳMY	BYwch���D�9�핀s���v�]���Kv�O�&��5A)��P#���oMx�m蘡,=Y)e�r|h�E�J�B�o�K���~��d��90�0R=T��z��1�>;�N�f��DG�*��)�X��]��27�IB�d3��P��gH��Y%�B%C�����n���S�Hc����0���\��׾��D�SUieTr [��&�g&��bs�)�I�~�S�$hj"��־��P����i����6[�j����X°O`Tr�2�WF<����*eO)!���\k/(�kon~$H6�3��/�[M+cqTWXѠ��h���T>U�ddXtw��`
)1-S/4tӢ�(z���qJ4�<Z~�^�B΋Wm)��&�W$����+�S�}�d�z<�0@n٬:XwF ���i
z �D�,�W��	�k����8,2���e��5j���e�H`��׷�S`2^E?Zݵ���r��o4)��FH*��{h��ɱz����c�5�`)!O������!%j��D���J�M��2����@��sܿ�	�f����.�3�ƿ/����q�6:�P��!/C)Qd�Ⱦnx�os@�",���|�*t�"`��ȼ�y63�isHh�"#��+4`H~���`�Xi�F��ď�\�y�e��8�Q�C�w�P�q��R�!�[ D�U>�m;�"*S����pj�9d�y��;Sf��,��&�pv8�d�T�E�q�S,�0㭥VD$r�����ت�ω��3ɀ*JIL�z�,��Wy6�v��a�o�I�Łq�U�۵���I�"���ݼ���h�|@|#<+��2�f#�bͩk�M�^6s^�;����<����	�~�Gm�R�;~G���"jzY�{W����S�0����$����8<[�F�*�`�-(B�͊�;����Vd��g�.|]u�n��Ӟ�������H��a�5 )F�O�w@����,,<!�U l���%�O�p~�0��F7���A�_�y%�n���$��Ur�w2�j�
DW{��"i* �{Xp�#^Z��Y\�H]��{W�����y�S$sӗ��&Gd�l�N�7���Q}�U�p���ܗ��e��C��X��z����ߋ!�z�aǺs�ͭ@��5=rK�N,���-n�!KG������5����â�� j���s�M�o��������W��&Qe���>s��8\fQ(���+p�^pZ3+�N��xW����N�:�������3�v_Dߥ�Fh��V�Z��,��kD���'P�_4��k'��8[�Q����_b�@�/�Q葉��4�s�H�}�訬�5:�km�D�&j�43��M���$ϖ2������p�Gq8B)|������ט?]���Uw�9Do[�3�u��cU����J<w8<��6��ʮ���}��*Ǘym��=k,.��v�������yL�"e9�a7ڱ(�"�=�7�P1���0Η��QPA�.�0$,{BqV6
���=���A8��� ��d�~a�#�V�K�-�Kml�%д��֫�X���cJ�����)��<��}�O�_�&�k�@$���z-���97���H������W �*���32�9��ջcS!�i*��g]i�'�ScF�j��b1G1�S:��]��{^7��:���(� ��:��M�CTg�6JD�����܄��f�����1�y��Cլ��F=I��`��h�b�3�����tդ�`.*|��:�#��"�UV �셱�zso*F��2̹��:�_�}Ƞ�4�Ⱦ���Ӓ��g�����r�za�58��<^�#�hZ}���d��0HQ��ε#]�˭�~��	>�4�_3�'-d���sZ�f���Sh�K���e.+@U��y\`��x���'�������I�c�ɇ��{勚�T/{U@lx~x5Bӊ
_���4H�M�H�,�'��$gq���i&�"���cd����E��bp�W.�e�4竘0;���X�߳�)��u�>0V�=*ʟ*�{�L�&Z)S��(Cbظ�����o��v��G�����cx��U9�t:�4�O��e�aɎT�JP��uKb^+�B�mS�f��	�K���|v��w!��ȢG��e��������N���_D�!]h�A�����n�ؓ�	� TL!7;����0�e����J�{n^O�6�P8�ݛg�����f���_h/�\��͕���|���r����UPg<d�J�����aZ~��p]cD|����݃�~�Q�&Xv�V�n1���93��I���}����V�{?��E�S5��`W���]Y�|���ՙnGEj�Rh+<��tz�6Ŗ5h�Z��r4�3�ָ�ܫ<WZ��	j�"�uȹ�녙�ǞV�h�1&+$�����}<6�_�N��f��'��w8��%����XD9@�fX:��};�H� I�s��z��5TkhY����c`_$I��?�ay�͊ם��1���χҺ/���*Qh �+�˖ߦD�'�N	u�c��MЉ��;���_�+��L��cǡ0ʉ���ˆ�-�''̽v�p�����.ۻs����hIC�e�'���G�&� |�Tq��6{o���[;Ԙ���
��~$T}j��q�ƢC*h�����w���,
e�[	V��ц,�䄸[���xZ����-�A�� ���&�~�Fm���#q��2f'�R�>�p�d��Y1���������ˢV��F�t���e�3�ɫ��1tQFNGt��n�K;l���*9����֬�h����Q��"C΄5�x䪀y:ە��&p��f�`���,N2r��}�־��Y�a�QkY2GB�c�-B~��8�2��c�FyR���%�'`�]1C�T"���	-��2$�/w�a�]܁1C�Ʈ�ܦ�I��-wE�Xw�sX�v��2�(�(>��|o��nnV�7�Y�e?OP�@$���E�$>#��d�b�Q�y�{	>,��$������Rr@S�/r�j�%�p�EGCց^������Ku+��u��W6B��#��W�)'�{�Dt����2v�-<�%5Tiq��A���蔳T�C;qN�*pG�r��0g�O�Rg>��"|���� '��,���)�N-