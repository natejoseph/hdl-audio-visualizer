��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��S3x�K�3�}���%�����8A����r���O<�`���434A�pK�x	�uD!��h&x�N�:¯+mf���V�(����4��Z��[������`�(�!����	(���|�ZW�}I�^p���^|� �0��.���8ޣ�I+�@�6�q�P�۲&�sY�[o�n��XW����"~�@5��L���s�ǀ�=��C���'�x��tP�@Z�+E��*GC�}$H~d��o�3e/lZ<��k�'�嵅�F'�����R�~k[\�b�%1X�a�_����y�:c���T�� [�ъ�#	���Z�x@����*}G�+Cմ��f�����Z�t���b򖟈�5�-��\��b�#�s*�k�Ȧ}%�A�֋�oP���"|�\�Du�#��t;6��:
���������h����7����2*-���A�U��-uzhW�͙�Hs*�� ��&�͞�9�Ǹ��osӢ��������>�㙥_x�/|A���"�~�c˥�r�+�(C�(N��{�:��7n=B��8�r���}{�.�ٕ���3�h�(GbJFr��T��&�Q�/��Է�D���I���#�����}�;��Jl�3��6�B�Ko��g`����;��H
�d2($�z�(2�ķ��U����Z��3D8���7�+Su�������u��-e�]r��ůi��M��������kb����Zq��X����i�d�����f�t��M�g�H��9�9�䥑Y1d�2T��~�Z��l[Qǉ����V|4TL���Bq�����H'�c\.\7,��Ӊ⽇
��pċ�q�$"�]�^�`�Y\�7f�e[o-ҁ�1��m���0�o"L�W2B��"M4�#�y\S�H� ;�:T�Ĺw�Y��-��f@c)�����t4W�Ǭw�V{/%;E`$�H�i����ԥ\3���E�C;1(]k�F,��Mb�|��L�y5��o�`�˰l`}�0r=���y����z�3��P�@D���/df�({;�30.�\w��n�_��#�TxLv^wo��4�u�d@/�tį�It���d���K�^���<W���E�sZi�;�y݁�!�$����Y��yK��'�X��e�vH��嚖��x��d̚ߤ��7AE�eux���@G*�g��_%�I�CQ1�� �ŧ.ą�N����~�pq]�Q�N�|\��;x�����l�����X'�~.g����p\]M�,� 0�����&*��m��z2��O4J8j:~�md��ͭ�#N�w�蕱$�o�Iv�f��h�����\,�������
q���C��
�I2��#��]MK�o�s���R)�{i����0�����7�E��0fb�6���x�qZT|��s01��]����E
k�y�ש�!�Zl�"��E��Wz�S-qA�I�˯�3����Z���E�S�H=I�D��k��-�u�8��udw�\;wA7ş�"��n	���qc������� �MJ�zА�;?�0�
A&�C��ҀM��46�b�j�w*Gw 2���-̙˙1�J��Q��c�wz�g�8�38���>��x��X�C�k&EJBo�o?�H��Y�����qr�i~_��\]��*,G��j
��3�����r����h}(��*������=��/�X�1�ʡ��o�K�4����0�X�C*�u�Ax]K/��+c������n	݁͛��:�Lܵ�)볂Ԉ��=�O<}#��=��q�n�5�,d��#�����J>�9Nťڲ�q����>O��������m��x���K+]�9��