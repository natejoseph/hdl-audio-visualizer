��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���֚/�뤕:>�l��7ϭn����ď,ttB	Z|�}�^��^&��j����)��\)xf�̉��d�F�P}�h��yg!��AK��+^��H��|�N�v�w`}S��"�<Hh���zN���`��I�1�=/��^��O�m���f}�߉�?�	���&ؾa��[��{�r'���f�;"�]�9�#���D���:$m��P�łr3Q�د��Kl�6��ɤO|a�_4N����#|���[�C�����<k����&KH���\��_b�YJ�^��aXK�-���.EB9l�pH�|c4�/Z���x9���>����V�å���m��/1#�G�`^hr���ӯr�0t
qƳaW�A��4�oش~�,Sſ������ z�e&7�Ber���D�̡+ٰ���Ձ��Ȑ���j��OMq ���c�9]���K��gwG+NR�S�mHZ��	��b��~�BTIC��_�Hp�G�Q9�f5!��GR&���ܛ½��X%�'	�*��D�����������۾H��3���m���o�I�T2�������'�J��N��]�~A�����O�� ���o� ������_���{����������sbIcߎ�s�`��N݊u���I�̏Z��:RJ�����~&cZ���PR�U��=Q��
�(�o��A�v��;y���ڷ�躠�iG�N"�>~}�8�jmL�4��˺V8;����
�e�vt��\����-���ų��)�3�.Jޭb��J�������',�wߩq[��EU�
�]m8�����e�� ����x_"a΃���V[֊ɓ<C���<L�6Yā��Ռ��Yv>�g�Bh��0���Q�,��������)2\i��'�VM�	�?�'orh?Wۆ�m�����ěH�,��:�]�X�����۾3�1�Z��/��� ����;��Y�����G�X��F���MUv,ɷ�o�Z��3A�ȅ+�"�6�g�`97<W����q?�dݪ��C��x�׵�dDq�JO����l�h�\b� m�
B��n������Y���%��9n�m�"���K�t�:
@�/9&F�|GQ	VMM����K�����xR��M�cnnV����G<�V�p��t����*�꣼�N�?���A�x��~7���n�CU˴޼M�i�j3й�zn��q�ż��aߍ�I�39}�khA�"�\j[Z�"�5,5I��;e�����n�}M����z�t�NH_�dt��a:�i�f>�=Z?���g��*���Z�x�o�-Ȫ7-�7�1����K캉|��2��d���_K"� G�u�?:�kP�I����	��"��ł|�Q/4��de+}�z�'�� �xy ?h���]����Y;�:Y8C�,�7s��������Խ�~�0�
�2�9/IŸˇ=��[ ��AG��M�s]�t�`XPz|Vfe\l����c+���W'@�ǡ��FB����/���o8���v�*���DL��� %�/-H%AO.Mh5��!^�U�6\��s:v>��DX4�@8F�\���+�'n�I�����%/u��1����xG"��BX�r|�M���������� ��J�dL���
$�md�V���]GG��T�����K]��Dt��ڎ)�
���7}	�9m,S,h��B��y�!d�C#�������v���1�c��EVG��F�(��~��;],���w��P�s�Z著��χ��|�b���`���s�)����)u�Q�1G Ҹ
��?9Nj)�Sn��(tn�E�c�t�{����|�%��[��颙��a\K�$���|P�K�!:?�%#=P�>^�N꣚�}NY�����IԙԺ��Dqq�Q�ڐ�1���^}���Zt��T�25	�}�M��'���Nup� �|<�I���M��nh̥�n�?��N�L�+0����+_�d!rs�\$&��^�X�:a����t ���y�����jt,%��X*|[�O�Dɡd��u[���s���n� �i��)M�~�+�����iP��e{�P��:K��À��j@S�����Nla`W;����`��7���"���ǥ��!���00�u3v����"~�$�l�R>2��9Z<I���ʷ�^pY�1��3Ǿ;��<���M�ɩ}p�Q�P}}�2|�c�0�a>f�=�d����,��?ɸ�8�en=�kd�<�y���UvY��x~
7M	��[?���T7�
��oh~�� ��Ѽ�q[��t89<�.M��K�q�4;�LS�qܖI
a�#�B��*iǃ0�ƵZ�����l��>��Gv��ٺ�N;���?B��g��)�M�^Ap�����M�� ���n𵥮�H*�O��-&)&i��^F%���p�"���}+���{�,�#ߋSj�90f�&�@������Ԕf�Ԛw:����L6}\���GHӡ���f[  )<hG�)��B~�o7���ֽa3 
�z��]ݭ*@�ߢr��',�?�W����&Ahp�	~���Lb��;�;����Ȧ�D#����,�Wa�zh6CLW�lF����:�I~�)�8a�Fp� �Ij������
�i\qK�f!,�`6�,���S,�v���Z������I��j]��̎���^e�i9U�U�����8�!�Q�Pg�`e_���_@�>e~2�~�
��\)�g�ѯ�l�rcD��0���/z\��['�����M��(�~{(��D��&���T(�$��3}$s��c�(�����An��Ʋa�G �x��\�f18=�C��&�
��i�'���rʹE�MpdI,��	���1��LS@��n�mR����A}-Z/�u'���Mz���/���ĥ
#����+ã�6��	U��>��>.�J`#��
f�Q0�\!�1�	"0�N
���+ƞ0�⢉�Bl7U�QL���g#v_��u��:qyK\B4i�@�I�y�X൞�?^Cԥ�A�A�K������ ^���J@��62.y��t�}1S�w�F��jÿ��<h����B�IH\�߸OD����>�tk�L�,�ʼ;���&���0͑Ơ�tL�7��-Ke��$$�er.�6�e�fX���FֿAJ��8������m��!k�n�u k�M��kYƞx�vWW�QH�IBP;��+# �7��1gU��9���̓�������ds�`�9��u>�y�K7��%���v0^�������+����c��$�eA$��3s�a�ȉ�^k׈W$�4䚘>*nY��;Uf)Ў�"�C��*��]��5��3,��-�_�{Z�r!�)�eC�PW���ON�S�[���D�8�u������&�;�Ic"�GN8|,��Wk��Pэ���'���D��U�7�
���$�壙;X�y����Un`�dL��np�=��N"�G2�����?1�Nl<��wm�Q�ci�4$��^,����y/�i���-�����w�ͮ��Nҽ��u�9�k�+�.�*7���b������T����yB�G�jĤ,�Y:Z���c4u���vn7��y$#Y(<�g�>�a�������2�ɾ2�(�������s7�uM/�O�)���� Zf��1?��V^� ����k�<?�ڡ(�@Uۅ��]�J��Gp��j����N6y�s #U��e�tn�+�缢�j���t�������@�u�#/2�\��E+kg�0Ӛ�����,�T�UYd��L�����ݗu�� oq=�Ϊ.�1��MS�$H�� >?�`��cƙ�|�|��/��\Q��?U(��j���� ʖ���^�i�Ҿ�}�"��]�����K�_(�*�$I�X�pu]�
%��8j(z;��#�\^�0��c�0��E5��+_k�fؽD"�MW���}������c��;���[�[�_V��#}aE�1X�V\u!#�eLD�Ĵ����><�Ĩ>�I���~y��q�_9�w�D�)v�mTNc?���=:Ộ�	�i�t��
�8d�,k.�S�g�I�mFj��P�T�ϖ�+��P|Ɯq����/ %���1�Cr�g�»*�'�&fV٠m*�th*2	nnY�� Rei����y:�f��<���n.T�Uf)��h֍�ۭX}Z4�
�[��>(*�-��SqU}�_9n0؍-��_���B�E�:/	]6����S.ӿ���Y�<@Mb{0NŘ��/��l�'��l���-��&.��YV�u����˵V*���H���t�m���C���hx��V1�:��j��4�2 �y�N4��q��y[��lZ�9ؾ�����&S++�P8����7`$QΗۓ慴n�� �L�e��`���{��Ċ���R�{��_�d�[��wR��J0t�D*�^�4!!mIG����!J�]��Y�J������j�eJL2��j7s#���њ��٥�ւ�v���(�p�T!�䭋c����F�I��颠��#A��2���޸Ռ�P��F�5�&�+���@�@�j_Ⱦ�Ku'�;)���=�Tm1j���� �)`���쩓e�XT��mJ��Uc+t~�v6�@)慅܏&V������4�M����姅�^/�^���L��&��k�g�[��	Mw6�*m��|yK��t*��b�b��-�cы����1�\�]9�[��R~�c���̏��D��bRk����"=@U6<׸����GC�跽M�>��5��:7�����)-���e�@�K�ݨ1;�nnׂ�}�D-������X�����&���������oOB�lΒs��o�u�[{z������G���.��*��ܷ���CX�2$*"�p��ԒNo_��7ߔ-	 ��kLH��qt��p�z�W�$��S�j��&���{��0Vz��&Y%�����ߙr�������;�J�9�[��CX�c=�KK��lSQ ;�l�P�F]���)7�Oa�h8,��}' �� ���?�#�I�,�8A��RuW��x��B��Xj	�ȗq~+�ނhEk6٫B��з}4E�:~��F~����,�;���
`�G&ʘ7F�%2�%��
��l�$b;%\jv$��UW��IM���Es��Hl���]�l����:`�P����4�	0�,��a�D�@��N󲓹\�zd(-^YD+���R��uD{>�[zЁ�ʿ-������*1oI�
�R��N^����#��C��i��{R8�(��1�񪻡A0TDÖ��2�DO*��h��..G�jÞa��c���ql&�����>"���Z�O��|��q���2�^f]�d�v���߻�Z����I�jNw�-[��hEסA4���J����^�*K�IoJt��(�|ը������@�����]o:x�:�.�0��o�3f����+���W�@LT�i�~Z.S�B"f��))���9����T��5V��[pǮ��)p�S��j�V�)�4X��PM�m?��'����J����3�3�lʲyl�>��	a�d<�efy	���J���̪r�<k�-��TZ��q�.q�:�U���y����.>��b�n�z���4�$�h�%���8�>&Kt���D�,�nρ�!; zχ�5��0���!>�d�1�6��1S1P�n���w~B6fn/���&� G7c�8�ӣ����zK��t���KIʅ���j�����Q2�����s^8��^�0c��0�A�x�&�k���'o8)��M¢,��Wq�H{�z�/@G-����Up��~3�*���۸��o/W�`]�Mkܭbd���5L�1�m���Q�ig6K؛l��D̎�k�0�7���X�%#QW�ȅ7�6�I�Κ�� J+�E�c�tuZ�޳�9�<�������i롈���R�˺X>uqW
F�Ŝ�ՠ�Nؼ𞒡�mF��&�Yɐ��=z̲��pHuXq�Lx@�}��`a���b�i=g������N�և�Ɵx����cwF����$�e�Y��&���`��jW�Nsd��4}D��ʪG�	����h(�P���;�D�P0~~�T�4��'z��,St��e+7�2�0-F�]�|�WR�������Lu{W��" ��2�y�sӈ1��X'��65ap�Dӥ���r��e*��o-�˻>·����7�uL
k�;?%^�0L������s�[�*C~��k8F==?u��e�K�S1=`2"a ͏Y�� �K|v��@{�q����Ӂj|�e;�&����NҺ�a�i���_���� e�[�p��>��5M��V��s�� w��V��4����ӑ��B8\R�������j�.N�>�$����F��]j�u9[{vL�7|�H"d���<GY�fV��E�Y�q��$���E͞jo��:gS�3�^�@��K�O)D�?5�|�R�j��w#20�҈'R�8n;,P���H�Aˬ
@���>S�j�	�B�%x�V�&D���fY��-�X�֥KL+���I���ϡ�U��f͜J&��wi����`&,�hн�#�ܦ9�7�` �#��s�&�D�~�MTy���u��qT�Kľi��\�Ds���Q&-�w�� ���.�t^���wo���Z.Zt$�������9V�qa@��ѝ��)(,�@х7���#5Q�w@�����7ֵ�c�U��l��leT���./`*����N�����ԧ�۹U� ,��%WEݖ�#~N�@��G��
���UO�ʧC_!���ak+iD��,(�wx��[j�ãw��$��[T��D��dy��Ħ�̌�e�"h�o�:YJ�c�IrB��1��m+@�=v��s�q
?మ}_o*v7��z����Td��z���j	�`�!�1nX��Au��16�?-�Q��F��1�?�|9�]>�{�}f�B�г	��૵vFx1M�S�4�V���t�?K�qm���"#x�Q�1�p�2E�@=̕���M��ǰBE����a��ͥ��q���H�s��PC>�-R���2��� ��G �oເ�X���2�;Q�}��R���r��EI<X���w�<��b:S����Y,��a�$-z��"fo]ҧڔ��P�3��r};�:«Cp��r�O����!��n�\'���ͲUGtGȚtq�4�n;����l�;�Y�Q&���
2q����

��Io