��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CG�ʜ�S��m����un#�::d�y�a[���d�������9��1�oJo��9�����,�F�m�هE�EB��0�ZD�[z?����0`M��|z[��;��Vw��\���Z���92�}�Ů��@y���u�
�*T��xP��b��(�b��'�wP�X�|�(���3ӷa׵��������us���Vw�:W��c�>F�?F��[���:��y�g)+q 	@H ����^ ��Y..*r��~dGә��-<+-���Ϝk
y�Y��J�Բ�(u��f�?�����6'�u/�}m� ��ګ�"��K��-XݘR��Hzj�moM�!{+8��W�:6���sp�0:�N��W(��!�+P@d�4s�um_�w���6d榄�Q3t�p�*�����E���e�lKr�)�rlaY�n@/4��i���.U蚎H�/����6e�?�74ۜ��+�Ж���W�D�����ݗ�Z�2�������!I�YYp�_�Ϲ���/JvOq��'Ul�o�ўV|C�HE?��3&3���4�'������׳�tV"W�f���F�J0R�_�"����a�u���E�p^�|�lҡ�R��3�����~vlT��|u����J`�!^�Z���_�h �z�aI�Ӯ$R�'D88lL(�����:�P��̼�?��"�*����� /#`$�X,��s�|	������喙4d�|�Qdd�@#
�\����@��cʔ����F˩���}AL����'sJb�>�L�`�#�9a�uS���7��A��m�̀���(H֏~9l��	���9���p�Fjc�;���l��_�ߝqx_~h��g�%ɤU(�b��xa��~z���k��=t��"��G� "ХsԺ衦5�C@<#!U��Mp� VGR�Nơ��<��'�5�Ѫ��ƌ]˽�Q�H��{���n�ؖ�G�6=�,��)5I� t�F��Lx.�͈xƖ̙w ]w�:�ښ�D��每�axU�����t�F�	r����-�	��`�x�w\5[+S��)PqcjT��G��&��V 	��0��Ry��	�a+R/^j/�+�%;'����{��}n�Z>��p����o�'5�����Qe �>�;.[Eߩo!�;{;R�q@���뤨b�|�؃�1�yaS�g�������"��:g���K��J�5Lw'�o7x�߬��3��w�"k�ۛ�0�e �6E\	e4�鵌ű���2�en�,����.�1:�	x�) Y�c���i���B8�on�/�@�j殅-6
 ʚ~��{rhՌ0�.��U�B^��qx � u{^�{Ъ~�Ƴ۽>��X�r����hp��?F�eHy���@��!�TIܬd���V����_��R��p폯�V*9p�j���>�L�?^D�.� U*
�����G�<T��2��른��V��n��O�!���ÙA\���+̣I歕y�)�z���t����ڴ�T\V���
�C�,�W�3�6I��\�v�⽉-�!�FV�P�P���=<|Y���S|�\Q9x�F�Z�c��k��'��k*��Xe.O��������eP�5����2���|`筯�w�3Lz���}#�_a %S(�;;����z��������ay���\���$+�=�S���M۬,��e@��E��,^�P��?U�l����Zo��m��B�`7`[{�D���`l�&����˘#R�b�9m���S1Q�w~���%�*�z�?�J�T����g��Q&���bÍ���x�謐�P�#g�N~�Q����f�u��??}il���8.�8R�1��xb�S�$�/�9T�~[+<{khn��ۅ��wV��L$qLmj��ٌo�]]�Eۥ3I��#����M�<2(n^�5���5�ar5��H~ ���%�-����-�z<P?�c�N���fL�q/�����L�� ~�zX��Q����[��"Ɔ��S�~��<H@����[.����4c�#�`a!��
A��Å�|].��sէH�tJZ��ܕ���VM�i���Tš�|���D��ޭ���%����M��w�i�Hc��쿧y��?im��OQF+��Y�� Q8C�˛�w��p��
��.��c�K��sg$4��J�?��ֈĉ���g��!پ��1��!����H(ta(�
�� T�O&$KXK/��x{�w/�<\����N��r $+��ƢY(瓴vW����I�T�)	�jghN�<��p?�2��ʝR�{f�y^�$u�ʞ�{{�I�Q���$�!��ܵґpAo�
<�^�(�3��/�ٚ�B�Lx2TV�m�r5125^gܖ���!��o�쐝	��͈i��omS�M�Btֈ'g���>��\.]H�4{G�Y|	���A����0?I�b���f5�tX�p>+�Iw�/=�����A�l��99������U��Ƌ��n�\vFg
��'_R�B�%rI� CC8ެq@�x�9N~I=�E2z��T�>[��:��4e����f��ۋn���p}ĵ����`���dͯ�����Xu������	���Qn�o�1c
�������[�x��]�#a-Fc��nD�|w�fR���K�� �[���o���Q�?� �d�+�Kj\ ��$aw��8o��0lM�͇kc��	+t����0�M�v.�k�pb�R
����?qrjד)�&�wsA��A5��
b�'�w���]���&�-��ކ�e�Q,���vD�	ƆU�l7�p)].�u0�����;�ەa�?$�)l:A�m��#$���X"m��i���eez�4|YV\z?�H��rIL�o����ݒ ky����p5zTZJ��^�iz��N^���DF҃sG�ѻ�ٜص.v��}�o��_ �0@�uh̡D�vo��y��:�b�3���A���Ά��~z��B���U�m�B��T�,7��v�������-�X͂�5I��L-L�&-����\,�#RD(�#_[}MH����^���l���/*SQ�K�$�8DK�^��#��5e��"Ro3����>aG1|��*��1��k$�]Z���}4�%&�S�X���$� @����ጴ�$�����{^�}_%Ã��쌄jt�C��Y�~1	��,nD���ѻf���p�~�X�fy��V�M�MU�Y���2��Y-1+����V����y�RA�UzF��ۛv��Q6�KX�x��ё�ʾLh��Q��
Q}��v���� ��>Ҳku�t<�Dj�]�}���@�!��mFeub��;�<?��OO�Ji�)B<�v49T=��N���,�MBA�4Mu�97M:���$�ޥ�j拆�Rlex��='�!���!O�_wLz�T��Ҡϕ)oD�-�~3@2�����h�馪͢^�&�����rB��.<zCG���Xbc��7dO'���Mwr��P	�����I��zQ�}q`eۢ�<2�hxQ,E�_�8�z�#��M�z"?}杹
:p�B���Mke, ���JN5`�>�	ղ
�>t�P���k-I�"���#���]z��'=d���{:GЎ��$}
����Q�H���r����{�]{�"�B���`]�+F&�Bo=��}S0�(�������Z٠.�7��8h��E��7�g@d��1a��̙&X+���(It�Ф|��η�kS��r�ӄ;i��r��XZ�]��m�ѐD�7�X��,z����y���f`aM�_U=%��I�DH�sg�Y�����f�A݂����4 ~�K��%ǯ7H� ��Mq]�F��.�)�ׂ������{*�]��D�R�������_|�:ʉ>�ev��n8�`	HZ�Ȑ��LJu���1���d��p�
W,M�#%�Պ@��A\��/�C��L�)>��d;N����`�~�/&Pjd�kv���W$��7�𑲬� �灾�Ԧյ� �f��;ghΓ����Cu���9��"n�w���۪0�Z���Nl?/����C�TJ�͛#B�e��u��cvX���0������>�Im�4�#t)��Ӷ��\D�>�$��N/+�:?�woC��r��g��O��!����zE��Lf-���'Bh�
;���^�.�6���dK���V*��O��?�� A�ا���+*�!d����)Fk���/ �h���ل�vڔ�*��O�\ڮb�3��V]�ʹoh�(��L�Q�P�*~3�u��T_��G,�^C^���>,2��h�*��@:Dc�e���	�̂������W�*f�A97�p��RKY�t��,�)[v{j���T�ߒnk5]����q&���xf�(��fC�6#z�
�>��~��|�w����q�&)��%i3��<�����
����"��^�QÚ����K�BU�����mƃ�^�-�-Q�^�_�\n��jHv�&�;�F��Ⱥ����Ԏ�A<*�c���4��Q�̱�ɪ�:�#ӭ�o��;�pP2���\�k�-_x�hB`�Q��wL���e���6a$�t������:�Sz��~�_S��������2�@�`�����0ҫ[��I�n,z�Vc���S�N�G��%�o��+(xppr��@H+'wk�%.	Ћ�G�ݥ��R��y��!�-�nb�����G��?����^Y6��K�7�Ѽ�
�O�R� o.;���h�k+h��b��0N���Y08$z�/� �y����"~���R`X���weC{f �Ǭ��S�1U���2��y��,���'^,&*�O{�Y�� ��
�a� 5B�:�Y�c��X�ȸ�^� {��NJ ���(��Xr���'�.֟�p���G���=ڄ�6�_;��l]�g �-�h|�y,��f��
��D~ǌөw{#�u����"��^#��)D�6��P�N� QL�F;���cǅ�9Ѷ�n���������FVM0D}}��3�{? �&��]�M$����cJ��Gr��]�`�r�.����)�y6�Շp���(U-�-�:+f�/�K\��jK9�ۻW#�(��ǝ��a�����*����(���\V }�hfD����G��3˶���A���D.����M �r3nu�-�.�ZU��8��#e�wߤ'=$��WS���4'�Q_��X��5'����;O�O��a�N����#\�˱w1tv���`�൪4|�9�� t��.�Ag�eЪͷ9� �e^��LԴ�?O�e�u��JG׻.�MR��*#�	ay����iBG���Y����)o�h�����)o�]oe�(7��55/'��(χ1�O�Z\S_����l��P�Ұ�D�FkL��Y�Hk�I�=X�������bT�8���<�QnSI�`G[��LG�IT�(Ka��7ڎH�_G��׾�q:m�N�*N�����W�2Ϟ���ў��!�VnKU�Gx�G�<��s�3�k�IZ���)��p��M���uo~,fo���ǃ�2��>��J+i�>)��vj�9���dg��/&���ƌK��i�s��[G�6��B`�� $��:�ϒ��+�r���#Uk��$�!�}>�\Wt�v,8���"L!Pl��H2����x�>��^=9g�'_��4P�w�	����a�^�U�|V���[櫍��D!��7��JoW��^be�C���.6��{�E+YN��(�g$F��n�
k������%S��,�*��G�֘$y8��~��,�_ȃjEF���y�i���n(v�#
(��f����bil��)0�:&u�a\�EL�LA�E�w��ꇻ\�/�I�Y��^���И<[&��������2�*��������c3[�k�B�����o4B^_�a02��� ;��T��׾������t.��0���c�v@����M�Ő�B�D��੕w���G��=��H4#k�L� z�G�Lņ_��oRݞ��Xٯ��n{Q���RD;@���(��gfZB��{%j%F����%礘��:HT
e�W����B��P�.ާ��y��ep��/�/f7������-��t���z�P?��K�(�@�)�%�^=�T@������ )��4�/X��L���%��`>�?�x�������˪_4D��s���B�;
;;�}�%-�[[|.�Pu5�eAn�V���Q����e.���s���`�/(tTyY��ʊ��/�EPAN�|2�Y�J�&�y���u�Z�����Cy�U�_w,��a���3:l��W瘵p��!P��E7@t@�1�?��u�	6ۡW��{UC��Ƴ�ME����GЅ��\�	B���5.U��>���vX���{aw�=�g�θ�����n�U�9�bL�b�
[69b�C�]�ob&J�?V�G2�3O���H˰(�h��H GmB�ղl� ��@֭�`}�W�%�$x'� ��噷�-��#g�+kS@�Ia�-��U�>��x���
C�&I<�����,c�f�*���SX���1(������V���z�8Ќ��{���Lܩc����c0T����/��t9���}(�R���+�:���Y&/��#������/���МQU<\ԕ�j��:��>b
!c�����;��^�i�ˊ) :�N���.��c�Wu08����'���l��(�ݢ@BF�=<Ilw�6�%��9�H���SgS9���T���T*��x#�wD�9x_�\o_�~����7��}�HR-���Y�������g��T�Y:T��co�T9 ���ݫ��i�M΃���bx;���,n��<CaUY�+~���mQ�e0K���e�WJR�}:��TP1�g$��Z�/���9X�j���Z�X��A��9���1� %@1�(Bs<�|�����贲ڃx-�'��I�O��ֿ�a�R��AR��4I�F�.ïo���W@�D8WWkc�j�/��U[��1��E����s.�W��V���B`/����:��y�#�H ��T�����G(I�?���&s*1�+8�5%ݒ^������b�7i|�[" PT�N@�W��kM�w�Fs�R�&�����H��%o>]� ��k&M-P9��Hc$|��@s��wQ@t�D�$�� �+�\{~��T}qZ�]㾭M�ْ���PtO� wgW����e�z<�3,��'��A��]��Cf�����=�J����C{l�BIk�-�2=����
�
~d´W1�.��\G��ș�:?@'�+��0��)��
OpQ�xv����/�9D&�Rpsy��
(�g�)���aG�f�`e|sr�LC�Ԡ(kRR�u0��ODf�}�Ш/k0dGG ��S��oV?.��E�rpQ�KJ[K
�.����J�㱘O�{� v�Y�7H�c�}�U!O?�/��l���Z��"t�Fy���`��Ԥ��f��זS��z�+�.H�R�s��(�ONu��^��q*3j=�T&��+�R��f׾����Ӣ��"zVB��e���x��g�R%�k�NJ}�k�����~t�n�s�_� ������&��;�2"v�fv�J�ǻS=D�wf1T���D��*Dfc�?���E�-=��2�{,o�sx"��^���W$n����pzdK��)���⠎"��=�������z�nP)��h��	�"Zm�v�U3�V�Va��h���T=�"�V��	����'����4��ւ���S���z��6��=���HK ,A���"�"��Z
�E�����W�Ѥ��5r�vsﺴ��AkH)miD%7�ۢz��9Qɭ��8��y�p�����E#�'�>{��>t@d�Jfy���K=�s\�)#I9�I�'�末�89QQ#�ӆQ���2�B�����~�~��F�d��U2�Ż�$@{�D�;,�&@��_���/�R���!�]��:�*� �Az	��c# R��u�������� oMF|_�\��2�<oy��x`�f�d~��%���p^�?�	���>F�+ct�|&v>Eɀ0��7q� �������sz�5�����qx�	aV e�ゥ�\:��+g���e�ߋ}D�TAI���CnȖD�F�,��s�Ǔ�HB����v������sa��lL3q��k]*�����1��Z��WI�si�(/mpX1q�[��$��q��x��BJ����Rʉ2s�w?�M�4��$
��p��
j�縬��P��)	��n"2��+�����z��^9~��:��
�L��i�����+J����o�gď�NBI�Qq�bL1�G�D� �G"^�0(0�gq[� '�z�m�Ja��~D�v'A�����E6�Q�7�z	5Ŧe�����KJ��#��8۸�1��Xv1�ԋ�{.���b�K�lmќ5�}��Q�_
��j�^ۍ�^m�{2���$��!r��\�&��'b������i4��*K�r�/n�([�D�Jg�\<��x6�G�\�O�q��8>.KY[�	��{v�m�&�8�J�v^�d���DA+c�W���brz�I9IX� �ЦwD7����Y��}\�t��-Q���g��@�!���
��]v<v��I�L���D���"�۠Z�>9� _��a�!�vA�K\AQ����P�[K.�����Pڲs�?0W�{U0�5GpH�e�<�ͯg�7���ac~sN� *����S�'Y}J)+���(��ϕ����
�j�=���^;����n�`(�q�|&�^���Z���B�Ï���Kh#ȞK�*��v��c�Q0��^�@̄t����-�e�V�^�\���C
B�Q�B����D�E"2Y�7�G�,4Z�v�g����jV�T�;8[ـ�. Á!?/�]"�t��}����@<��
�����\�GehR�g�.lU����КS�E~:�'�B�q�p�J�
=��B�KX��}�ո$Y�Ԋ,)*�o��S�OHn~W��P� �k�@H^�W��X�E��V��`\��Z��y��[��� \���<���{њ���""��7;E)I~MLf�"k�BHҧ���׿+��ᖎ��D��6W��F��ky����/�Y��Ϲ��b?�|�ZYIċ9�Ir�vH��B���۵��*�<���n�P�(��oU]��р��R���~|"Du�S�^�/�Ѻ��z��il?���F��X�%ev�6�����ޜ�t��R"Y��O�ꏊ@�uD�z����J��q�HR�wϟ�b> j%I8��ʢ����:���1X���3|)q�u��nN� ,ff�~6�ٔ���/V|�:�&	�s��-�/&�l��y?y8e�Vk�|���{��Vw�_dŇ����MGMm��?
G;L�E���v�@�c�N,��/�(�P���������h��{����m�ѳ�DݺΎ_ɡ�,u#3H{rf���R�J����#3��AHA��ӶV�(	�C�q�zk"�S�1��)=�2S��41�>�ʵ��j� r�v����Ϩ�kbY�?���K'wAI&��Np��b�$U�+8�����s��Ճ�'���/1 /�Ք�������j!ʕ�_'�����}�����p�/UyeC/+i��I�]�ݨ%'29�R��-��9x��B�:}9�W�w�Qߩq.�r�����j��uS��fQ�� ^Uj�M�����L�#b&S�*�
��H���/�.���^��TX�ˇ�[�������W��J�s akU/Q� ��1�ct��'�S씴 aH���\���,�2�C�ם���i�k�.e � {��4-yX���/���2�g5:���f�e��`c:��L�9�]�r%�/�8�VLgȖ
����:iJA������\�ΫX{]��2d����5roJ5�M?�=Κ7d�zqwG�eyE>pIv��2����D/k?�s�8p���3lk�2BuC�����m��:����kY�k�}=F��`�O<��Q-����̍]���X��{�"#C$M���+Jy��[ڭ�Y����x�?f���ӷ����k���
"�6aH��,~9�us�-k9�q5Y���.,�?��Nb�Q��f�&-l&� gFXtY�a�ԑ�kٷq���@�m�9��	��yKl�21K�𩗐i#�;�;�tPb5�3_M$
X�Ί�&U'������G�Q	.9M������R�M���������A#��Ņ΂l%%*Hj�}y�%���j,^�#�=m[��@M�h���,����RC�y�?g'��{82Z?�c�1ۈ�MVܐη�'M$����pl�+�j�k�p�ݻ��=nK�ȕ!Yq��b�|�ɍ���o��N�||P����`Z�6NÄUc#��(�H�1|���<��%�����YʬB��(�#��j^v�v�n��+b� �(���֑��ef�~�=��Pґ�.�lъ��C!�{��tq���8�/,T	\�򣼠*MR�dI����#QРX��rE���/���˸:o��r�qޗ�����?r	Ō?/��c�ـT�����D���l��(?E8��ׯ�+V����'țĨ�@pQrh-��}͸�M��C�["Ɩ�������PG/���� ������q�k܇�ȭ���� S���nΪ��#Cz3�N�wc��I+����1I�^�%�*���Ff�/�<�u�
�^����w�]d=v�^D�i�Huu�
�Yq�x��\j1�^�W�^�+j4�(�h�J89�/l�2QPa��O��(Y֯3���cft��,�@�9G���j?��+�~7%�Ç����~�0���U�K�`ӼEzީ�4ޯO-|���>^Q�ܢ߿~_�%%-�W+H�"Z��+Z1����gNy��hĕ7�@����̳��3cL��wc�k�%S�
�#
��V�e$~�X&Z�;: �d�-;�?U��^׬�Uy�~��1Gu�����$�sU�� ꠑg����fL���Y�$�1��QJ7���A	Rs�I7|�K<!�ʢ�K��?X�ZdL3s�(�ޙ�4�g܆li��(�WtϬ�:T��ר��e�������@sm�1n��h"y�'�ә��ܥPT*�s\&'n�ܜ�HR���@�x^�^�ݟ���K���0�}����j(����I�U1�v��f�Xi*v"65[��[}
����_�%]բ�RZ���� 	C�?�ӗ�u>/]$�6e鰴n;�^ܜ1�h�V&v����C�y"	-+'����p���6�	;>DA�,~���yܬ�l(]����~�]���>�f�>`��Xv0���+����6[>>S���ф�l���ϛ��������)����Ue�Y������#�^OS�!���c,��H�	e��oAêeYV`T8� b'�.grK�a�+��G�RӲ�̤I�.o�הh�=[?��5�;��~D�KW�Z�x��AY�����:�ѐ�\��\lQ�b�����ʙ�o���0��ӯ~ �΋d��qfp�n�q�����l��LB�s2�7��O�����b,���/-�{A� �rR@y}�]l�S��Ӎ|z�V/���(���a�ݮu�q�e��6E�e�s?B��{[���(�6��~�h[��w��G�U���4��8Y,V�WR=mQ�?;݆���c�|�;����w�qy����<�v�O� s\w�P]���T��NA��b�I�N��4�oL&�v��ǥI�Fr<X_W!���b�m�di��H0?c	.Ӗ�r7�H
�I�zW��nܛ�,�����䔡֖��0���S4��¤{sk��t�aKc2��<H��#�Og��8��N���/4�3��a�Ʒ�c�������LV5v�t�O����0;���I������:�����4~5&-����� �Ao�頩/��Q�2{��0ǚ����l��'X�ƝE�'��]�[}�v�$�� yˏ��!��[�����z1v����N�f�zƱ\(����I���Y��W7���E>/qQF]Ƹ� 3�$�4�I�5[��eg�Sz4
��prC`H>( Ӡ1�V\l�����<�]��r��ɸݝ�����Q/a����'I8�6ǜmmgg+���o��}8]�T��mu�?K]&qჴ36�����,{�J��8��o�f?��wr���J�
�n�X����q���n|-�׵��(,q,�`8'���I,�2&��9xM�e�b�Kr��S�p�]}(S ������j�er��da�P]"c������x\��K/�\)ɒ^�xM�MeƔ_��϶0���ؾ�Ϳ�/"�L�o��ON�J��
Q��R���M�Tk�1U��B�wE��������6�Y7����x��|}��� 6=�!V���Ǘ������Y1�����%Yz,ȟ��^ ��=%ŧBnS�����d?�>+̷V֡!ބ_�x�ǐ��Y����\�f�p���ʂ{7�B`�-i4�+}K�_����z M�#��UN���3}Ǥ��]j��+B�R�T���5R�����
�n�Ԅ��H ��~2�H�N�1ΆR����x�	�};}#��"8��}��8�]9�-�� ��Q~hǂ��+��H�:
?;��3�M�T��Z0p�WJ�͝	ψ�a���A]oxh�S�8�IR�'�up�&C�	�ɡ���~;�cn�{����rX�Z�h����K�q6��s�kl��@L�刲0�1v`�kd09��5