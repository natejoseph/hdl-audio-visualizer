��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CB��na��v��4_u��ש}6L#t����b���_�`������Dc���rf�p�Y͇�O�@TK��}�,jp5��Ub6}�e��������HY�q� �mg	��G�c����RLL���=jϙ��禺dX�!7�%��Xv�A묇~<�5r�V�V��|����:��lC�����T������E���z|���p�2��+/���HP�3�ra
r Ex$}�4@ǐX^�_9���9#f���`%}�!Ԇ�	pd)c�+�R�%~(+x끱�!�p�ñ�|<�������F��.��i� L��"�\���c�l�����]��5ҥM�i��rk͊ep�in�CQ�)���僎�6}�F#"�~���D���I����g�/��@�q����M{�9C��ybW�yT�)e)[��XSz� ��U�%kg1��� 1K7��J���94n~��� ���%N��[{1q&�gA�S�v�va�xIkl0����)�^-���Iĉ���>����՛�Y�y�2Q����J��I���[�r�ڣͅx�W�<�j��u���?g�K�*Ѝ{�i���A���^�04P0VW�益2�y�y�m�߳�|#�q��^���[&�ɁAwe+�����\[�6������>�����H6���h��&cJ��~ 5��<���熥n_��QX��1��9HІ�T��_�����HB���2\��_O�Ӊ�J�
��V[�l.7�m�����n�]�|U����4�a��f9��zU"��1�k%�ڭ��s����c�7�0��[A>;B�����t�_��r�:!�U��Q��{n���-3>u�9@��pf	�����۴Q�X�ݔ� Q����Y�;~0/��5�W7�Y��0NXܭ����	m���4����Ͼa���X'=O�e(���MQd�Z����9E�+��wjuWp`ʡ8�{��8�Y�1����Ea�O�Uٙ�L'tW�{�����O|���dam���fs��5:��{J�icj�螁r�O�i�.�h�O#�r�������Q�dv����U$i�h�_u���T.Y���'�(G&���g���*�u�ٺ�n�ܻ�p$�{���s���N�x�������Z�9�zv�8���d��۽�A:��3�u#��&#����',�r����~��J�L���"��hB�0,�g�����R�QX��[%6bzP��b��"ڝgٷ$[�a	"u$�����>c������婗�!�[ Ӭ�C��;�^�Sc��iʌ��a����;�F��eZ��]�m[%)�����N�qݰ��3t̍��8�2��N��7��K�5�F�q��~��9JDx��+�E�Ր�n����?�>��,���;�>�˯>��l��-��#S�ȠNb�{󈁐9ƥ��k� 
2�͸^�V��!��ȅ��3rD��b�Qs�b��y�?9*��:�3�G �Xn+���?jXe��0��y�:#�ϨM�]��k�w=���jo��:�8U�Ȅ�!$^/W@�T�J�SN���*���ġ+�m�E��J� �s� 2�~=m�0��8�=}ۅ$�3aq�x�7l�SYXj��M`���^��.�蜢JC!qЙ���`�#�/�����%m�5�c��켫gc�׎�|(�|uN�>B�Ge_���k��'{-iad�p����
ƌ�'|h��� �*Z�>�ɍ�R�e���}��l��Z;&�S����L�n�<�n���l�� �vZ��&�r��ciǤGa�CbH�;	�̲2�/%��#��_@�j˟�	��ڧU�{~�Ξp�t\���BW5��K���p2��-�L�y���L]�$�|"u����Q﹗ ���{�h���`ҏPkL!���y�r���^�5S&�������LJQ�S��*�5-[\l��J]�@8�D=H���
F��M��Xy�0A����wc5��G�
�wɼ[Iͣ �����o�z\[�S��3�4�%AH\k=���$��'k��Mf�OJ�`w��#���ku�v�s�c|G�Fh��,�@�M_�?�~�����FD�
ޛ�=��HE�����g?����PҕsC�E���+�&-bHxH�s_�-��>�"Έ�� @��X��u:�#?�iJ��ᕣ�&�8���j-tl�*��_Fyq��\)\��ZׂbX)(�'jI�f����`�W�ZV�U(#Bn���^Y!���~+.|=��[�!}�)������֊�ǆWw��IrC+�?vRr{CޠM���N�Y&'�fLN�!d����*�/:ԅ�^ğU�Sf6[��t�Z��y�>�D��A�U��fpͩ��1۞�GOU2��l��'��!���M~�]Es�DK����7B��*�ag����K�~�E'�_�x�}2�M��8���Z�j�'�k���M�;�O50*h�[�XfP�Rb��Uc9�i?��Wf����l�@L�
��嬴*�^J������� ���f�x�9��I���f1ixͻ)��G@�r��Jщ!�hyH!�� �T)���rQ��|fsk���R �b�xQ�;�HA��zޚ�W��82��p$jc��%�1���Ə�4I�6�^�AH3���:��N�X����6r�SL�.�!LK� �㌑�R�|��i���)�2¨aѩ.�y+a����5ϵx�xX��*�=!��ū~�(O�/p�t}��
�Eg`�hGJ��9+-)�X��V���(����(Fx&^!�P͋az�N��0�[�ԦJ4ػd.k��yr'k[@q$��P5��c�o��,�X�ז�m����a��I�I�d���"()$��!�.'J'5����\nM)����ۉ���2ꍦX^�)m5���>��ME�.灞9�s-��O\Zr7g���;;q��@d�B�/�,��� D^#��{{�v.�J3�u]��p}�mQ�`s� X�/�Z�P����P�����=q�
d�q��(���}��Hu�7�Ť��K�'���Q�HY���&͟�p�xd��ApkN|�͢G���w0��8�˾b�0���Z:ԩ��P�����Iȏ�R���e9π1���z�E�{��0������L\�C�/G��i%R�˚P��h�y��X�<�*>t.,�<�o��n{^{�9�7<.��|n���`	%����Pr���%�Y5�4Q��0Ҏm�O�aׄ0c\>���U�U��D��3�������5��ί�� �(����G���tB�'���O㘑�c6R;�Y�|��@]S|yqH�����PNp����p���!k~%m�������E�r�B)i��-xUu%��BJf��I�x�����Țs��
�No����YϷ]���w�1�Էݼ5pRT�rj���Ou�Cig��A�Z=d)E��H���;�
�kT��
x�i��5�b�;[��Y����2٢]��!s��(�r���%��ћc,�Z�n����O���������� �D����Q�fк.o�4�\YϘؒ+[b�@*ժZl�.Sj�`��
�	IR���^v�D�Bcl�:G:K��M�KD3�0|f�����S���Y7�1�) E����q����`�$g�/���Ë�0�|��v������^�'�>EU��`�/b���Q�n`{u�mL���d����.���P#J���0����]K+@Y�(d�}��u�_�*���l�A+��~ۉ�s�
�t~�{2�_s?�gǲ����L���=��腡��i�0�$O����;��2���M�� Y������&�¯-�c��3�q�9�eZ�;�R�W���.�S��w��$��Eɋe^c�d�j�l�53�R߆HQ�x�E,d�k�J:�e��4K5�6c�Lλ���!���m�-����mi�,E�	 ��
�[bm��*�����������j߈�
�3[�e@۵����#7Jޭ���� n'F�f�&��F��F���[��4�V����2%���Y� Q4l��� �s����3+l4栤,�����#d?6*��BoF����g�e�C��.�p���7��,`-Jڦ!Yj�\V�c ��1�.�~ O~�1��v� �y�]ǈjZ0kM��j[8[��
r�Ft�%�I��jP�;*� }����X��M��b�(� �+PZ�݉wDM����'~�|��}噫�Ͽhv��P�Vg�^����G�ƪlY���]�^_m:��K^��
��m����>QŉN�8�G�s������|�0B!x��a�'��1�Y���G��S7n4�X��nc���3�"H������LM<Jʶ�4L��faѓ/vW�������N��iLph������(�~��q�r��9.[�d��~u����⌮����zK.�D
�u>l�~lU����j��7���f�>��@�{η"ə�?�cT��#�o���&2����،x�^XQj�!�`�(�H��\[s���ao�٧�tk�:V��@�R_OI�Wv3�Ev�!k5}�.��Y�e�xmϕ�c��;P���;���5K5��؆��B\�3-���fbV��[69�bi��r���#f�~��FI��n���č������V����W-��\���7�4��x��YOÓ�L�T����5K/
�pY����L\�Y +ԣ�b�yar��:�\uL]�<��
D&�̯��Q��d���*V���]�x#��U�QS.R�Ҭ�T�!����/����gS��Y-h���c�'�\����sJ����|���c�]��k��kj�W��&��¤u�ե��)n�X��v�(�~��s�[���:�����_��V�~)�/������	���(�7��x?�S��>���|�����I�8�n���4�:l�%�Sm��[�}�7��R[^�}������m��AT��,��1���okw�-҇�++o\)�id ��_r|\��n�9g�z�h�������IN�Y�7ct�3�(S����`��N>6p��;��R��Ь���� �F�ו%��'W�d����tS�C�ĝg�.մ�[|>��j��s�f���^��G�Oǭ!�F�E�a� =�m�����I��Ѽ�BT"��_~�H��E�A�~���3^����I�pn�[�Ơδ���ތEY���7�z+��skDԈV�0�\;;�@�+�+��T������<����MD��e���vk��X���n�v��t�,��+J�e���r1��5�p���J���t����:?��b���� }&ؓ��
JX�x��6��La`�R>?�MA/���~�j�}��Y;��?�T�e��i�$����b�ϔg�(��&x� �ⳔC; ,Y0N�H�Q�V�G����������'H���!�"��kJ)z��6[�3T��F ����ۢ�^8>��꾪�F��fRQ�T����b��$��;���n��tJc]��b7,�L?���Ŕ� w�<�)�:�M��ڶtAM���`�H�P�w!���l:_vB�G�-	��i��QK<���hi��tT�����3��Z	���O�F����
`LBi(gI# ���Eƺ�I�#O�-ތ���\�Y�4o͞ZkfB�nLR����bZ����p��9N^�+@k�"":�$'��k
}���1�<�>��[9l4N{�����P	m��2�E^]@̝X�F�N��²�ty�,c�m[�"Ϳ	�d�N�B�-v����|�K�j����|��1��^�f��I��rɃa��\�V_:�i	��H��! H�Ps�Wv�fәճtG-n��ү�8����D��4���o?}���v�I�Y��g�!������Q��=���@q[}�0��B�vwZ Z�;1�ka>���^�}j�r_�����9Qw�v�`Jaң=I�2���H��C�e>�v�ĕ����u��.�ʱ�xJ�gd^z�V�i�ZY�Lw�$��_��ʘ�SZ�#m���y	n�ɀQNr=��1�*~k?<���8,�~����9������&�u	��^���W��w�<#Qw��,^^�T���Ɏ9��d���zX��f�柌�Y(�sYf0��0UG��P/�w%�1��z�$M&�A�Vh������`�%yL����N1���o�|Π2YeA��*Y����X�b��Me)�.�^����&丏�
<�~k/Xf�4~�aȼl�Q�1׃�mD�j���x4���c@;���Ës�j��^���'T����O�ET�����d`b6�r�aŰ<��JNl��S*�(Sp#��ӬL�t��|=�4 !�r��V����΀��B}����z��֠���ڦ��rP>8��WG�����17�B1RC��th8^���0��ܓ �i¦��T�FZ��S~v'g�� ٲ��W�W
�l�iH�ew=�¯�$���Lg'� Ί�4pQY�Q
6�BmS�����xDSz�w𳢖��Nc��	Mq�[c$����)�x�*�N,Z+�����v[\��4���%���_��-�g�M碛�/��!��_`iX@x��E�5�����$ᱭn����yL�=ţ�/���h���0�ek#<����L��Ar���b�0��h,�\��^s�Z�J�@B�jW���M���\�����=[�0�B&-	�f��pR��J���N�7���i���"j/B�RV�5�9Ճ���c�P�|ޔ�-ܳK�Hm
�G,�V����T���}�b-h��]�W�L��dl��ɏ��x�ǜ+z�E��d���@;�����N��b��RK�!R����Ԟ[�O�:�����Xu�4�N�����������>������I�/��
�XT����8��Y������A�'�Ob6:�f;-�t�8f���>o4�r��'��
c(O| �)hM�NuK�C��U����ӰŲ��9@�5>k����3�>������:«{o�7�@��6}����iM�����t��
���ĳ�M�Z���@@G�o�N$;�6��.��t�P�o!����N������9�7��X�هY/�-���t����t|W�!*w��%�:�m��gG�=Y�`F�}4�邸��Wm?���EƐ0gx1���h�QF�E�#Bu���6S=��x�"X�M6����$�ߜ�<z���G��Jć�����(�V��+��#,�T��o�w�5=�np"���w�@&�@Sx��T��Ӷ.>��MG�"���%{a=�"-)�����.?�K� q�Z^.��vßS©�w�h tF2���"�8��PT� ��= ���Nef'r�'��Xy'2��t�Q��s�Y`��n��S1AqJ��6�C�_��㨄��	9��tX����-eB���R�d�u��(��?�#�h#�]�K��1֐)�Q�F����Υ{F��iRR�O���=9��y$�%Ţ������k�H��e���S�l-�L*��:���L�$�Y�4��4��!�A���Dh�D*�(�����>cy�˽��X\�Pثޑ�qЯ�R�>�W��˒!SP4� L��s��ku���rﭣt�Ypt�I�鲛���>�Xw&�+iQ���cO� ְT�����ө��8#Pw��2Fc*�h�9�X�� �',�!���X���?��%s>�����͜��wl5��<X�7!p>��Զ����E�|�6X�q�5uļ���D5�as���U���o���N��y@wR���YuF�-wj�P�O[�}���K֔~^��eJ`�D�T�`��E�k�����R�X�U���?+lf�#�E�4�믡�8��76ǚN�T{��k:�b��