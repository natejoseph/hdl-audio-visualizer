��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C:�>K['Q(LW�,W��:+c|l�@N/ٯ<:R�*C�Js-)
�-pȎ�e����Wau���#�U8z�'�5�FH8=U�jIJ��6�5�I�ϻo�Cldy5��1�y��?�cΥ��Gǅ}��zv�~�y���	X"~��t��V "j��oL�F��lL�,����VH6���0gA�;0!qX{�Ο��z����f6��^���<>?��3�ш�������Հ�C�>Q�@���;���;ZE	ۘhE0�:a�/�D�W���b��.�ڡ)�#%��:D�ud��@��=on���|�C����,�Li���Y������4�(��W�Y�+�Z��J�5-*�	+(C�}tt�T-�j����3`����x� O?n�5ʩ.��"���P�kYy�lŁ����p ���B3 ������j�y0D�)�9y��+�`�;�o�a���+8oU%z�b'=����d�x8T�m O�ٺΚ�c	�TJ���%4\"0�������YSf���$�N�*&�R*�3�p�{/��<�����H���;�����YVO#��!G��'!��YJH��)z��~߁&�|R�hUfsk0#�����vI��\n�o��Ի�S��zN���*�d01�Uո�2)��u1�n�������J���u�Q���g'o��ɱ>��q��:�6�	���R��א,�o�5v�c�xr���c\o�8�r"�agR{�c>ݼ|ΙQZ�i@�J�!�	��r���x����_�M�3�	� ,�	3�0���4�_r'|#���|[�)P�I���ӡ�����Yh�\N���A���5��QS�#�Q��|¦�}O��co�YD^�����8�@�%;������'�gJ15ʗg؈�h��"�	-d�mB�h:��gi����?�h�;���3��:_�0���Kx�a��X7�Y6�n��cI��[��p�
R���jj�J��C?����V���qs5�-���'x@I/�������.#1�#15��N}��[����&\�j��%��T�XJ��wkmV��a��z��$~�}R	�$�P��[���?�g\Lu����yFCf�ɿ26 a�3��*��`Xڂ
-L��63J�b��l�]�W ���ǧ����h�X:	^fk�zryy��e��M(���n��؊��F�j/П�3s+�k<�&��[��Y�	v�)+Y@u�Dtp��l���
���?f��� �X����F� uj� �g����ڦ���vr��Z� 3<�]	�&���_#������C�5_��ָ��8O�`�4?sR*����|��RUo�G �8<�6�9c2�$&�P���Ĝ����d��p�r���d��"ǈ��
b)�����E�U벯��S����<��1���<&�5e�/S��
�4r��:�J��D��"'R[���r-௃+VB7U��l?��2��\�l�f��1,�`>��M2cewE�Q�d���d��}P������d�L�8�|M
��0{ruGۘ3ԉa�O
�Y(%����W$c��9��?x\�8��7���h$߅(���C�b�_@w��N��W�O�U�]�3��Avݪd���0�9�]�:�/;���m���}ݯ_��D8�!檁�^1�����XG:���cQۄ2m���!f#�ʦ�&��+!���L�㼫��QDu�0�u[�8�\W��t�����n�(��<Z��Ȑފ�]�������J$�V�?��#0{�}3b�� ���x��Ye��4)�Ѹ�@��7��?��5Y�_/�+|O�a�H�
�K� -DR%I%���A�F�R��g5 	�nMQ��.���v��G.����� �W<"#�����I;c��&y|��s{���A~hxp�W�V�r��bt�x���W0ʣ_Ĕ�ԣ��7ٟ�V]�g�w%Ϩ&s)|p���p����Ђӭ�F���5����r{\;��C?�,\����r5�G��Je��� U6���D���U,� �5���<z��|@Oʳ��D����~�� ���^-�},:��򺭬�ֳ�=��Z ��ǥ�"?s�G'�{�y}�Q'"~��u:-�(�gL \�"Ѳ���\1��V��?�}n);Ed���P��(���@S�?�-������X��y5*�+ؓ^"��x.��٥(�}��om��ѽu_���&ޮ�?�f���P�L��X�K,��>{%���� ��sP�/�2}�Y�l�hy���&d��e���L��R�O�<�H��X؇�wZ����@3R�Ջ��<|6�9�a�|��5 .�������,?��m<�02zw������_g�C\������f&��UU�e���j%SW���������A����a;T��+�a��_�f��R�� ���ވ\3�ٞ��)��j�X?�B/9(6��Z����+���8�	i��a���W�o���9r�SbzBh�ߺ'vx�$C���|��(-'�Pk	�)��s���p`=��M_��XA$���Ҹg/�7�Fv�����0�`K�Ί�8���B�`�n�BQ4� V��&��Q��"E��p?]�:��Z�~�@�h	��_yR
� ��e5ݨHqh/A�
BKGp�Z�'����i��[*I�iʫц��؊���rͬ�ZKl:��d��	s���j~���E�l�?˲�\�5t��/�n����I�W���l?�	�Q��-�iՄ1NWH��=�2��#>�JO���4��m�L�!P;,0]:��B/�t��6^��4����bR����&m�5�:cH�h�,Kr�l)L� �s2ӼZ�:�HB|3�'��T�we�ջuwa��;�6�Yl'���h�j�y�'����#7q-��J�C��	��tHa���u��ɞ@�W��P5,;�,����Z~�5�o�E�%;�q�Ӝ�+��[{`=�_�h�#YR<!S�Q��k��a·�� tO��������l- QS�X�ES"�Je���~�����Fۨf�q�)�0�ck{�8{%�
�$�FH J���cx�lQ̐eY�G"�\3ōJ<Ɨih\S�ܢP;s@gNC(�����[e֦(u�ZxH��|�T�`��!tR �wxt^te ,}�U"�/���A{�.�1������.�<�w�]v?�f�=����,�V3M�b࠽*��e3�)��]��FI��\�ۘor(y&^i-���7J5��dF%���
���JMCvٷy�뱅TG�4�����\�N�ۦZT��I�(��ũ��H��H/�%m9e�$����Jy|���Ž/*�N��Z豥��Q���$FǋRU�<��t��&�R��6�b��{��[��3�_w����Zf�����!P�"�xFH�&ak��cΘ}�F���({�����?%�&9�9��W��	�������!�Vw���ٌ
���1<�d��W0��A{%����XL����I���wQN �\��$�${
3�Z�m���b˴��oڶ�_�Ų;^rEd�'��(%�5>3'dꝯ<�]蒻vq���׍%��uQ ������<�[����"z<�	Nr~1�œf�D%��^����0p��x��!�v;x1պ��|��: F,Ȇ�u8;�XSګWc�\Vf���e�AL����;�ѱ���Di�{�wx���P�U�Ά���k2h�*�����W�s������.�7j�_�b1��nەH��w7�C��:�����7��U�ס�p:������ϓ��R�oL�2yw>X�m�A��cWGe+��.Uf�}��G�:�T��{���.dl)�'����`��NV���1�%��G�y�ٶaN�Lޅ��@��*�2��FS�C����=r�L&0�I�1~b����e��e��9�F���D6�
Իl�ۧ+f����K��O����w�i1ߏ(Og%��V��)�<�. 쿢)6C����ʮ�u�
.�P�RWjiKS�(�N�Jk���Ņm��D���׃�φ5sq��ֆ5���M�wh���r�T���K�ȏa����,�%�ّ�����BV�����.4;,,ه�F� l��8]�@�!߯����y�IR�y8�������6H�'����Y��G-�ù(����MÄ��7�N�g[�{B�a�Vuv`�p��LŸd;��&A�?�Ls�B���y�t̐8�A�H{>�͍�|-Q�-r{��R�{
g��.���-�NQ`͢��=/�W�����
�$FD
��B�+��_e�  ����t=�<3t>9SuB��mU�3}A�-Q��LwZ�c��~�H3�}�mΟ��9Ŧ�[�T�|��xI^=t���ޣ_e���r y"jT��bB)�1dģ��4]w��e6F���I��Aɶ�y?F�0��U�:Fb�/�jLA��-���]��a�c���-�JeT����d}�>Uq[�����\�۱�\3"*�	��)�`U#h�LO�Il�_IU5.\�A?D�a�}L��%�q@T,��6|�V2����ݚ̛N���Lg���vw�0p[{tz<�Z�tN��D�P��J=���8�@���^�����}�c+�| ��z���xK��Q.�ix��Ү��2}�W�� ˨��U擴��%d}z����#@dd�Q��npn�D�����Sj����؇� n�u�R��8�gR���_0�ըnq�P)�q`�&����E���+�i�#R������ip1���0F@���td�Mt�\;�������}��WX1߮������L�8"~l]R_l��v�U����C1G��&�+Y�E����@.6͊gbc���2?��ob��� #�8�I톳�D��!�f�纞��)�����>8k��N3�e�U�ٶH&�� SI��rNY�$������z����A#��'XM��)E��ۙ��`��f�ϳKX N������l������T�JWP�
R>n�Q)�)J��-!	'W�|�(�5�C�6���?�K����O�/2�e���D���EJƳ���v1]�AM���L'��H,ζ8O��,MC����11�Ćz�IT�!����fRt�,'⡎
���(0�LZ�}�!p������iA|{Ks�~�RL��ͥ,9ؘ�]Mu�%Ϙ�dg���"��3,f�N&J���+U����$�[�W�k6τFm6�C;����{Q �?�>�`
51B���9�H��yzҕ��,DN�X���)e��S�~a��p	#��E�ƃ�-�v���]��W�x@5�}դ����p	�-��y4%<m�9e֙��؂��Ю|�ګz��Sû��D�q�\�_�[|���q�_�Q�8�5�9��C��?V��ѓ�$�T�a���z�.Ӭr]�W]@�S��ڰ�\:�k�=��)��]����{�h��o-Hzi:�����f4���0�t��$�l3�����S��>t�A�|;�?������g+�|�kJ�����0Ξ�U��[}e�=F�X��/\�=�V�:���ay��BN	����ma��+߁^�{�&�����H�=�=v����L-޹_T/Ս��;e҂����<[���<1���),F��w����5M�R+��&W�XtT�y�7�|J#���x��~��	��"y�� �Ud�|�]s���9E{�.�a.Wk�(�i8�v��7��
�SV�G=��]��Lڃ���qAQਁ����T�&c�0��Y���_��d��Q�`��Z��BՐl� �\fo*7�Ȓ��ϊɦ����_�2��bn��	�S�*}�sԣ���jk�ع�߳v}j�s��inĕ��"�
*�CTH}��+
�k�DFi_�,h��M��[��[^
��cF4H0�p�E�RT��Iȥ���].��1�)7q���@��P���\� e粳]H�'
ċjث�&U*>�;��Y8(?���C#�*
mqȐPu�κ~W�Q��a|K�H�=�
��s���Sv��B$Iu�P��0�J�~6�!ܞy��u&Ta�>���~�;�>l�f��,��e�I*��{U!���e-�&9\�q��yO��)+��Z�����y全^�-+�+_��4l5�o��~�D^Y_��g
�_2�5Y�~I!q?�m%�$��1����|:$r�Hn��ML���%�S�J�lQ;�6[q�.�˼�Lk\Ҝ�3��	�z�GVe�=�`I��=���������x���3m���A���ѧA�B��5�r�@�,����l�,y|L��NMz竍j7V}g��d��bo��ރ��!6��K��巟�A�OK�E�l:���I� ��h�|�Mv�g�B�w���8�+�����uSǲ�ݷ�2Q�D�Bl��#j����,�����G��"���u�-��@��@�6"���W ��r�n�_+F���@P����B�Y-6>w�"�ҳ�'$�Ůlqh�������u􇧜�+�x��r��	GN��TJ�_v��<m\�Dκ�G���) P&m*=�d���nn~� e��X��[P�*2t*�μ�ke�{�\�S,}Jڃ55G� �b��ѷ+
���B��xwuj+�a«�H3+�3W��=�\x5���w�������-[�*��FѶ�ȘIUɉ]�8�O�9[~��<!�Lt)��]k�2���Z��l�9e���ퟃWwi��:�,���xR��!�V���z���?�M�Q-�b�\zK���\�i���_��B�U_=�s�zj�;�Ɲ@�(�O��i;[��e�'�vg���������y�t��,���p`�6��3k���|zt����>u�I-�P�[�K���ov�!w�*Ƒ,��P��&z�����b�䂕G�� �a����@,� Q+��� ��j�}�[Rm_R6ݩT����uǰ���C��c�o������jZld�N�zZ),��Gj�yN�ݠ�*�ݔX������&�
�N��Ut��%��(�<�Rߛ�@$�t�S�0S}�T��ݺ@y�V��>s2ŝZ:
�J��ؗ�U�,�j���@zuV��f�{�~�A�I[��튟�NGLB��k���[��xx�1�G�V�H��q{j���QZk�1��Eh��AMG��;=t���EJ��B*)�㓁�#�I���N�k�Ɔ�ÿCS�&��{��S�ᖧ���z����b��1�����7Q�.w�T�p ^���$A�y1�ԗ��j���>�;�l�T32g�����!�p��X�{z����[:�(��yY(`s�_و��` +��h�,
�"���������*d�|���ԕ�>��'�5�X�:�_��+�7��Cq�J�{b�}��Ո�`��cI��;�L8L������_�!?l�B	��AjTfbk�i-�t~dT͛j�I7�s8�`!K���|º�}�$Z�{���|O��3ԗ��oS �#���@O�H���5��{��M)��N�=
��#>��WL��	��#�C���.ξ��l�`�[LĀ�mch��;�~��w�Q؇������7c�:�wu��@����lS�ݧ��ZE�Bg9��:���f���@��'G�WԷ���2<��p����.K�[+��i�o�3x��3pA��g_��$9:>#y��ǻ��;�"CÏwοe&�$��s6���:�dߖSc�B�)b���� �nSgU�n&b�H$��7���>h�^REp=r����[��I���q���)�j�qb��ҝ���D�t�Sn9��Rmm���P^&vf��X��H`��z<x�֦��Tk�A�N�@���Eȍy�v������kǨs"P�wYO�����Y��_�y������u���w�"������G]��əx�DN��*͠P�3��
XF����~��^t/s7�'�	�/7q6S�����ͼ��G��Q�-�@�K6���w("!<�7�E��p�O�.Iq�iY���)VR��H*��g3��ǁ3V���]�G��B��jp�Ayiܫ�#oq	k����`�<�*G�o�1鈲���q��P��k bd���Q��b@����e�|� ���_��T��k���/=XDDY��3���KGxg*�&<�ʢw����Z	�!��Ԕ�#�)��A�P��Lgg�����������Z�+�	Pz8��t�����I����O�Ru���#m�����+� ���p��׼�n����1p��J��é��K���T�����'o����w�Ĵ]-��d񗳭]���������>��Xc��^��m��e�'��F�Gx�Hڕ�ݪ0Y�V5jS�"5U 2e1Y��[[�����6ܮ����F���B��5cqcE�B��ZG���o��2��u{޸;䮗�,�÷x���� E�\��b���N��3l��0)Ry	jJ|݃�aM�0���jdѥ�M��`��9ľb/%=9�Lpzb')��p�0"��'D�EA�L��0�P3ƕ�4�;痪�4�}��څ�� �p���5�"m�����D��aU`���5 �-�������3Q��9�dE��)$W[K"ۑT����Bƌ#����q4�	�c��Ŝ��X3�^��$P�:Xe�$}��|�"��� Gj�s�)�
��F�C�h�H#�&�����q�W�y�T���auӺF;y��|��>��������8 Q^�� ��u;�)�+�V���� �)2\v�w��D��#¹4Y�8�g�y��)T�<�$d���>�-�'%��Sw׻)4|퓹Y�Y�ȸ��;�����>�Lb��֣wZ���y��-9.}@����T�1�K@�xz�-ڀR�=ƚ�c��89�m܌u�s\���m����Y�PfEKpZE�x��Sy	FdM�c������ĩC<�kRH�����:�-���D����0v,j5����$����Z��q�҃Ǹ�� N\�?��G'�̠����GU��y�n�6�膙�$��X�\�^xK�5���٦�T�fp���魻�� �U%�e&=ғ���2k����  ��3wZp#Vo/m��n��|��yox�˯�Y*��:�)�ҕ�V�@EA�5XK?�v_? ������|/[&Y��2�
}�����Z�T�0�N��D�����k�Q�� ��XV����t'<��\[z����X�
�M��ǳ�f9�|8�����.��0����7e���#����� �y�-B�n`�$J�RbF�O��%��W�x��� W"�����L���h����9f��_zI��I���Zե�Ż�y�q�㯼��lxT�sVg.v��|a6�R#�u����wT*V5�5!��`�	�{9T�T�����0���ab!3��7��օ_����h�	�B׳gq%�)�'8�I�'ʖ�7��o�&ϓtM�7�I�N]�Ԓ=:�>�� Ű���k��ƑF
��+nt �7זD� �{�f�!n���e��:�˖p��`#�&`o�w.��a[NEH���~r�֌l�Hs�C!l�;��oc�hc�����������$Оd�-��3�pC�[��v����//==�8"mn�&W)|�YN14H��t� 4��O�wt���[V-U�:O�o]	H��3F)���\��~��k�`ke���[<�0�s��ɓ�.}��Jt�v�����G�;��걀Lr�s/c�$�z��W�2[F_�z8�����sΓi�kSeG�C�Br�[�v�/g'����U$�CLY:�`_zH��)�Q�O5�@=�eq\l�<�LqA���i�Jd� nO^�z�C��/N����򆶿�KL�z��Xa|�.�ϟ[�!A���^���.g��z BI@D�2S*����If���vmC�g�G�y �X�I�ئ��9c� �&�v.��J��F��fp���H����9�w�u��^%;�����ΒA1������Zq���jp�KAt{�����ߜ)�˴�#tɏ�T���i 8��gX���&(c0��Y��0��KV���Y����H����Ʋ��M+>��h�V�V���'�,�W�C=0Ɩ3�� R�u�rMX�˝��U@f�\m�o�{��k�~��R	n�5[Sk�u��%�D�4�4پ�a�8H���=WYf��T讀���^O���wb��sO�%n�H�u��|�	Vjۊ͖�5'�K|�S�,��5Tz>l�|W�ݻ�zA�d>i�a�~=`W�`�R�:�n;/K�^��'���I"(�83�I��"b0�k�v-�ӝ�����	�oL�Gڈg�����(x�6�_���x���3g{�}�`�[�:4t�{/x��M��}hȑ�d�����Q���T�$�p�})F��;���&��K�(��k�/�"� �$F���;v���#$��+�`"ap���϶ z��H\m�����W���d�Eoi����O�q$�����V�E�^7�K#��'��ٞTV�`���V��@�Ϯ��ƭ�Gk!����a�t�ٯ4���lM��
v�p>����x%#t`#Y����l�t��EZ'��G������7�CN)���؀XL���J��%{�pI�;�^}a⭠�罪2�=�KaN����MR[VȂ���Şʍ�af�l�%pZ쒲��"�7�"O	b�a`4�iC$Y�s%x��օ<EI��61�Q./�����4��y���7}/�$�ל��]z��S�n�y�?]5����m�2�e���e)"#k��[=���^���BX.�w��@��4�dQ���ॐ���a��c��"� m�ZQ�I
�ׂI��+hܸ�o�|ǅ�ͬus�䨰�iԇ����DD�J�S�7��_�M�6��c�� ���s(S�jF���ZFO�
�[�����1d���j�6��5 �\Ʉ�Y ���}�&]�^�&��:8b,�% SF��*�jC�V�9��@hʕ�b�3:l���p�Vis�e �1T�'RI<��rz.B���>Y
f�j.�
'a��Z�4Z��q�Z�;�a�m=����'-U�k*q*�QfH���
��FU�5�����<
D�:�KB`���>�Ņ� 	���v)��P��SI�c�MƝ�C	U`�׊�)�٨���bֺfdV�_��8���f�x�L�U�O���T��(�[`���Ap�I��8eg\amQJr���x�Y��F�6�p����0<3��Ó���L<����q�]�x_@E�9���$�{�8m�(�=�Z�W�ABɥˇ�vv秐Խ��YK�De#��4+GZFv;({�`b��Y�c�%�/>å�P4��'o3q����y6��oEyL��]?����>�&��ǀr�N>���Hr�S���)$�M���V�L+�t�S����A@�Ȓ�ɸ�1�
�"k���\�Ok�c���*��_?�GE��Ѿ.�U���m��fFK�!Xf4Z�-�=���L]�D6�����9_�m���.���Zp�̅�}�{��"���r�X��Z�6.(�EʞA�lV.`�� 
��o=s&��y��hk���_��s� SI�p��g�a1@`����9B���|� �w𗑩&�ʎ�v؈D�ʋo���!�j�Pi�ބ'-���b�]ɔQ��X!D�$FY���֖M
S�����%�]E#6�mwCP�/�>�9"L�R9M9�P6�W6;Gp��\/J�\�m9'#�(d�h����6H<�zP��i+d��i-n//�u��A��R��a��Ú��K��x(� {��E�<S�2(��n�"��!hx���ϲ1ߦ�̅�L�@��s�9�4\ ����VVF�RZ�׊"�8�v�#`r�g�ܲ7��PWR.�o �1 Lx%� vWU�1IB��ʁ�%��0Q �H [�?����F��8(y��U�<�����N� l+f��,��b=���;L.T6&it�.1�[�,��Ɉ"|u/�p�����4W��?5�fM>��3�����$�k�)�.% 4t6�YA�_"%*)�v(zy�N� Zq�qs2��ٝ�O栕�D�#���h�_꼤+�hS��A¡��_���ʃA. �st�۫�{~�$#��!�֡��Fc�	�\��K��ŧ5WQ��ع{̹N4�$xr�'���?���������.���AƮH�n�z���.VO�ǔ�a��t��ˡ����杻�(
	��G�]pI��VФo��
B�
���/��&)d�q�,XX�Y	1`I<X���# ��%� o�0�땉h W���$�FJ
���5'��h�q���j��O�#����1���q�d
��>H��Y�-uڒdS�6�W9M8��W>�����ТM{� c�|R�G�!�`�����MV�
O��~t�����V���0�s�6g��%����Q�P0�c�{8�/�⃜-���<���k��FJ^��������/H34.2"i���[長.����a��-� s��`[9T0y�n^�猑4��;� 9������:�Y��th_�&zf:���i����"*�r?��y�ڶ�o.~����Q�Vߕ��d$����Mml���{��Oq���T��`�dʗ�j���l�J���s�R����V;Y'6�;��{��
D�����S<C��<��y�~�tD�#Hr�ݑ04n�u�$����MoN��-�0(��PJ�氽I�-4�v1Y :�C�i�Nֆ�T�lM�����&>|ds"�X�bI�7�34��?{����e���y���ϝ��8k���I�/�'�gG!�7W�JNg��A{C�2��S+�Є�)�qq��cz�������r^�Z���o��&�ȸ��?7�wH��;��!��Ik�|���&7j��J;�NZN���=�r-���C3}�ߑ��,WK��ǿV<4eD�z���ݶz�5�ǌ���b�Z�H	�4XH	���g��r4�ݗU�z�m�x8��ơ��5��/!@$&��A�w��u��J�����cP��������g��`2 {���t��\������n����i�8#(&���Ӹ �o�|���Pe�{j�n�<:L���rU�w*��ɚIqQ��7V
�'2�M��O]^!�=��'_�9-�Pi
t���o��wLO~CH�؉�D��-ha;�$�^�WzSЛ{OD���D!�u�wNgAx�_$�s
�i{�0�s��;/+
1~�g�{�z�$�-��]W�����7
�l�	O3ᚒU�۽T^y�}2�R��]`�A�Ldf|��Y�O陦{�Ak�K"���<�{.:+ql�%-s�z�vtq��u��D�(�4t'wVW�䈈{^��7�_5}�·7�ɖ/����]�m̛�oq2H�p��,�HY)��^����4���E6/�*�\��1|Cr�分z
@�.6bl2p������i��#���-��}�|&!�{������N��s@����prR%$������2;��r�Jg�*l]���,��ȥZ�7�9��ؙzT���,=U�ЇO��&gr���<�`~?��<(��$٬���i��S��ֆ���}a�����&x�BIsV�����)���AA���Tވ��W�����BЍ�b�J��=�V�V�;��tD�c��WQ���y8o-oi��C��|�����ޠŗ|)�4H>c6cf	��Pĺ)�7��KƱC�<��:��}b[�^P�О��$C��g��\C��b���ʂDȳ�Q�a�h����=������c7�H4� װ�
P9 .�U���;&݁`�c�|��u\$��_���rM5tn�,�E~��f�~1'e��W�_d�`@w�j~MYN�܈��f�>:0j���@?S��	��w����+�`�2�шG��nW�LF4� ʚo�] ���b_I�g�x�DSı��Q�Ć�_�dX.��_�I �1�k{1�D���k���"��p0 �@!Z��uQO��ݜܚ2U��6uݱR#V�PX5#��g��҂'Gn�s���?�A4�.(�����ƨN�5�N��e&���8����B#�����s���~tP"�ϒ�]�0��m9p�l}�r�>� 3�D�'MV=�d
��D�#y!�k�^���#o˫C�������M\���[��C�M�R���DU��NS|Y/E"���xa��h�7�
|�!����J�y�c�ш�zv��ޒ����(����\ßd�:<?�$(��(Qs-��4V> ��)�_���,/O{��'��×o� x��[��}�vwHkb`>��d��uz]�4V�u��qd�]/]�4�NS�`U�� .Jٔ��6D��<`����0ւ���$l������a�S'���?��s#K�~i.\>�W_���hx�G�M6�/�v�0ْ\���Ņc�ȡP�joo��٩ڿ�^�wi0�>_�IoY�,S�+'�Ƭ�9�������B�<��3��0^�>����Wk�������壁��1��Q/�zS��6�滞��3qɞny��~�f(�L�sƨ�^2㼕��\��6�����6������e_��})�>%���@�� ���S� ؝��*߬��<ŏ.-���)�w��Z�c{u��5�����n=��EO/N4}����ZO���13�v�2����'�N��7���x��K 15�>���).��M��S��=&H�=`f?g)����]�U^�s�e$A:Y�������.��Ԝ$�}�6��D�.��Ys�	��\VHۮ��9�D���%-6��ZĬ�BLb7ȣ>�2�g╏�v��
��Ϊ(G��c�C0�[,~5���q|�L�{��]/���<��)�n������^��	([�~�9\��NX3۸�e�ƅ�~@"pf�I��F��=�����(�; ����~�u ���w6���s�ށ6ɒRK�踰��}����^�`��צ�1M��M��#&�wz�*�g�v��go��{�E%lqл�9�BHb
��衝�Ɏ7|���܇�#�+5I��6z�~(~�J�4w����9�N3��eҐ��� R��l;c�dn�`�Փ¯h�����YB�(7��vJ2���]ֶEo}hu
6�}M���o���K�X*�>Q��{J�Pda���1Q^Ezߛ;��5���^hc�Y�$��4 -&�	=Y�/�S'��ho܋�CI˾���\f����#:�|)�G��ť��ᰘ�jf�|�)n���֛AP굳���V֙A`GM�P�.�����Υ֢��?�%�+@d�Nni-�tE���ƹZd�>l(/�~��r��>%0���T��[���}�< �m�Kʑj��E�.q��'*������'m����
����[�@���9�(�0���(a���ɇ� c�n�O�m�.�\jt����b���,�7��3���$��L@�S3���E��̜���nl��l�W�p��&Kb�u��o��T�3*�IJ�^W�
C�t��Ӑ���aޚ%zw"o�'�G�2J�W5Pqos"��o��L�DT�qCn�X^`'9�����v�~`����ӫIG��R�Z�h��1��� �?\{��"�le��C#���n��W�zu��ǟJȑ��sgGLd)%�Ű����K�uYE�ˋ�)8���Q���yrb�W�^v.ؼa	�I%�,��)�Q�P�Ӟ,]�*Q��B�,j*�)6��Ѝ��M�$S�Hs(f�>x%��
��G�K\�ЁP^���T��tMLe�Ph�1]��c@�m��M޾���w�d%4j<�t���O?�y.G�(J)^���m�j��W��t4�ϝ�H�>�
U*z��	��E H"������5�Z*h$S�S��X�CEJ�;�x2��"���o"m��,J��m�G0xUb�4F��ӾC��aY#'��b���ZJ�DM3�50@FT�
�^Oz�ܑ��ɺ,��sB���
�8r��A�L�a�{F\6	[B��������%+��4�Ɨ����;,��}W��$/���ұ�4D囔������7x�!�&��|�)d��.�Mb(�Y���"����2�`����7Y��8����o�5;ZT����X[�x�ʜ�H���_�լ�dlo=��Tx͸h�c�5M��G��1Ùl�e�!<b�-R�#��Z}�vR߫m�Y!�:���FY���e����%eT����<)��k�;o�F/0�yJ��,I��+�Vʆ����vB!���lY~�2�ю]ɝ7zQXc�������H�h�yTN���1�Z�i�&'��s^o��md!�@{�o��Il���*���}y���}��O��G�IȚ��(�_�S������Ns��3gJJtJk���2�j�Ϻ�����?��9��Mǧa@94�m��nw���i�ZWG"����5aL���}�:��oE�b����֣ֶU�C�ު�[U��	���d�I�Ĝė��4K�$�a��V�LH�iF���Rq1a'+�t�8����7�d�B��d1�At���̂	���̣\�t���]P�l�'��ã�%D֍���!YfחS��}-q��� \�^�H�y����VĻB�:,x�?�EC	1�,����F��a����,���'\P�{��:Rh4a*6�`"��.��Dߡ�y=�8z�}]�sWP��H�W*~0=���P��#ɡ���������B�����ALψ�rͬ�ǵ��h��g8� ��BqW��Dh�"`�a'^�g)'-�-Bq=w�oT�I&�E<�0K�qO����Oy�11+�_�(M0�4��vB,M��d��J
.l��p��ʢ�PJ�}�,0O�'
e����9�UF]<�DT�G.��n^���Ֆ<8���$���t�
ŀ�j�]�.��/��Y�$l%�­{��(D$�DvI�����Y6C�vʩx�2��k�y�̏Th0u)dҒ@�#���*VrW�L�Hɍ�� ��X���E,�g4Y�����#���^6���p���8?Y�R]��H��s����Y�h���.~н�B����ĺ�ӗ֖Ņ�x^m�{��w���%�l�����F�h�W9%Ps]�	h�_���x>O�'�\9�Ĵ�|�d�Xn足a�9�<��������7m�Yi�r�:�}�}�jц�.��;���3[�-�@l���:J�Us��k�� ��4�s�t�DǟΠ�ʪ�*��)[c�Ė�
�@{�V�h�$�y��L-�wh��&v	����Lep�z���aT98>�*'-���蜬��m��⥓A|�g �l!��i��nf�-�Sm��"<9�K�J�$�v�Uo3�S^w��͢}K�ب�z	D���2-_��:tՖ,�j.���[��,5���]��\��f<:�<�?˸�C��� tk��uo���?�����I�t�%"�=b�""@ �_�m+���1�
<U	��_�F�*0%x��
�%`���E���̇VM�8��~6��uBC�3�� h�z���R	U��QT�M�-%�u�FF�sj�kN�.��]OG~���V�g��dne����$��=���h��<'w�,8֛{]�y��;�.�����w�"�@�Y�Lx�0U�_�v�Oa�Y.�/p���i�M�X�ёD:�6�C�4=8"������IƥR)^ �D��$-4c~���J�����g��y�Ḓ�+���7��Ą�7<.h=Z�G�4{�̩K�t}I� �b�Uڢ��|��������8��-��*걭�$�E-ߎ��j�n�Y�~G�%��C��b}���ey���y÷����0����5��ִ�y�q���d�>�t>��܌;���<G�m�P�3���9b��A�a����,�2�
�n�:��^)c��k�pdᅅ���N�����M/2��w �״���"6#%]s��x�|�.�@�e5���� �:}m�9�����(IAm�7x�/k���t(�sv&S"��<óNhM�T.��%&ة�����G��;�%x�������'�����u����+I1׌g��o.U��$O��8Й��>��d����f��<ڪjHn��(���r��p�����v
��!HC�!ȶ%�2K�%��u�<��8F_�����Oql���4�j7KM9�P+p�I�IMSMiE�g���T����/��O��]rn=�~#����� �Dg�7#8:�[�ݵ*�GG�B���y��7^4�9~�PF@�RF��]@������(.7�.SqD���nJ']��#~�t��������� �44O�#�_�$�oh��F��5�6�Wt6��t�C�� ��Q���E�V�����"���D׹�p��c�iX���O��ɍ�;P\8�+�Xv�TI"~hG�8@("���Ǎ�dV�RՖ{.䍄-+N�Ԏx�_�T�7������U�_�KO�4zCx�<�Y!i> �&���j:Ys����Se�F9拳���QWn�����J]�3ФG�-��#�o*5�~5|�Z��V���"�*���tL�t+�?*v!��ܬ!�g6�6����}���Bfɰz�����V�Ԍ�q��� �g���AFrkb}��w5]]5&;�f��pROkAz����w�~qN��z��v�X���6�T��o%�,!	�+
'~U��@Ftg���@F�n�d2��j��K��nNY�6����P��H1/
=�6�qdv�[��Hpd�{����_A����莤^�����u���Oz&��-�\`��)���)�s1i�|����yN2�#z�l��Krj%d@��%�=�u�X����$�)W��h��Hd ��̞�dA���]�i%�ׯ�n�|�Ք�����������'�?%N�������KRvd�S�$.	+oO�< lL��RE)���7֕�!\W:P
�aV���e�8������(E�~qpf�zh�n����vC�z.�tA�����L  s>�Bf�t�y�س�b���4��sv��x�=~���(^�މ����E|乸c�#❍����n��3���y�~C��S����?XXj�_-RLz��FS�`�2���`3�y���]��M+-�2I<QS	���e����t�PKg(ȩ1���1��Of��zԳ���n$��O^���T~H�U��� �*^���D�}�Bޜi��(wl�|A� �-8�dE��Ô<�����T�U
(���W��L9������T�Ǖ�&R��������^o4����'�N�赊�Z�^ȍ�cX���U�������;�.���΄>S��(�l�}h=IHASdg�Y�� ��`��R���J�ɬ�'g���I۰͛g�\i�7��j�nO�����tvF���Mf��ʱQ��H���@�m��S��I��Cx��9;P>a֦t��1L���5�Jg,:h�zB]1
�iB?�L.d���;zG�����`��\���@��g�5�c\��@ڷ	3J���cg���~��	�i� �����G���"a
����,��6���@���S}u�����FJbh���������8fe���Z��f�����d26�F��-n�s�[Ñ<[� �~^A��5fK���e��/T����W��|\Dm��͜�v���1f�ز�0Ï�����l����n���|��o�$��������[��2:�mVL�YH[#��LR��2��	�f��.)�(X�\�Eh��2<4�D�b>=V&�I��CG?
s;����A�
@P[H:|�e�U�OAB�LQd�`P����#̩!=a�s輡�M0}�E���`�� �(�QoXp�2Q��}1���|B�[Xz�>���ʂ^��q��a�AWw�c����FO�7^�c������30�Sd(P���fu�6���3!~h�qj�l�>��Ӈ+�P�����lC�{%f�?���b�N-.��YЏ	�E�}s+&!D�Y,�ڦ$\lc�3꙽TY\ӂK�;$+������S����h��a�/A���Q�Z{FS��ܘ�6��5��~C�s'�|3��l�=
)�����)�"�%�$C��4I܋N���L�t_^�h�TS晕��얟�� C�_���x��!,����q�M����d6�O�
�a��'g���0���o�uzv� �aik�,�h%��f�\'�U��wa�k_����}
�SS�W�56���"	��Q��s����f�J�"wn%p�����`$�-x�Z��c>z���(�l�%<�G㾨��hP#�&����� rU��gVg<���7@��%g5YA�B0���*�-c�d�S��VXe��e��F~^}-+��mB c������\�Յ�n6X ���ow�7� �
.'kzx2��ߙ��\=/#�GcP3��O���j Dq{� uQ?�ЉdXS�mq���i������N6�(�b�[�������e]+��.�����+��7R�.'9�%{6ޤ�����9@�9n��T�J�/��J��t��1��s��{��f�X�U,�S�x#V�DX^�`�C��n�leq�S�'���ʂ�4vn��E]�L	�������[ה���iRe��?:�d�o>mL�i�� ���z�^y�l̟��:��xj��0�j���n�۴��W�7}Ń��my�ń���8��z��=�'X��y�����G�2:�V�2�O��FM�ʭg��B��oō��|
���*=؊}	v����H�nX����e��̠��}͑�+�d,�L�ǤU$kl⾷Px�����o,"y�]6�5�q�'fe������wK�\r_s>Z�=��0�V+
�q�#�t�V���=F4���9ˁ-�����P��:�^2R��b$b���Z��L E�2R^4��K����h{�0��H�N�t�a^�X��T8�'z�g`$�>�T?�=@P?���\KP/(A-��lh�2��T�!��}�Vċg1��.��f��믳T�����*�7�U�
v���0�o���؟̗�����W�ySAG�ߔ���oޓx��x@���@%!n=��I�(gv{h��r7�Pi���S{�;ʘtA���̬�|��rw���fΤ*>�
�$��0�3M!׭mƈ��0���J3�˪�m#�4�M��'ʶ�W�(1���UD4����YuՔDW��#ʫ=�Pv��Oߙ�)���%��3� Jk`9<\�Sf{�鵓����6-�<��P� �+��	8��.Z���q� �Es�G���ǲ1��$cv�Mb���|�$I ek{t�S/�ةC���᱁�2m���D�_�MU�#�h��K���u?)�-�V����C�M�ӈy����!�ғ�@�l��N�<.t��q�#�y~5 $�3EO����}S�ok�Ml���}�Qٞ�T:��of�y7�#� ���C�N�s�*M1Yf�x��O_�j���o �2	�3�R!�>�&m�K
0Vz���w|t���np��l�,�O��d�S�%Q��׬��a��Mo���u���ٮp���/���X.¨�$+�*���&�!�,p�3&Hd��j=U>6��!~�O�&�4`̏����_�����������m�R%��L������W����n%�̝H1�7X
�Bi���F�+mнg5:y���rz�a�=��*��jG����Ɉ�9O�P��f���P�� Y��#�y�BGr��2B�8}ɴ{,<���H_���~5����FY�A��d+�neCZ��8+TzC�f`��]̛�{*e��'�K�W����*L�!�v�e��{壘MUs�b���G|�]�q�@�X�F�C���ܙ�e���e��B�
h�B�������焒�P��f�&�7����$�aQ;�?v#��dѪ��?����"d�rJ���}5s��,��e��*�_���R�8L�)��&v)������
���ia~��U��@et}o2uP�v�����j����p��OH5��|/��׿H�Ւ\:5|p;�A���܇�XW�c��L��_��e1���mQzWPC���VE>���wxh���uxbіzGV�OT(v��{�bb���u�#�߅M�jLȻfs?!�&��X����D���	K�P��������s��43,(dR�)M���u8��x��u���
m�_!����;B9!TX�vy5i���nŤk��� �@l���h���TT�*Z����ZF�'�Sd��)*Z�9�@n��8�=��j�͎�}N ���k�v���բ�q�0��xɟ]z���8*��M�{��ŀ�DFj�t��2�O]�:���%����k��b���憶'D��YXm�s�)��2s���w� ��ԭk_�N,���?UL"�	��>=�<NՄ�m�6������I6����I���6�9F��؈W�&�F���F	��}����/-���F̔�Sۆ�|��
<��S�b0�A����9��[Kn*��M<I�D�TC&��4�»�R���d����%7�Tpc���Ɍ���0e�E�MoX�-��7<��+���{�{������O6����P
��=�����]h����AY�`v��/�|o5�9��{�`�H�)d0�b4oՎ<��b��Yk-�<��W��D/'P�y����<VBH���L@�,���Ê?��~���MI��z;`�����_~򺜓Ӑ�n�pNk�	�'�L�j�T®�@� �U|�̫]��W�'!�e�ī�A*�ְ	@��.�_�ۥ�b���k�A�{,�X��֡	�4ۜ�tެ,֒>����ɹ��F>䋃=�=O���*�]7���4r�De-�q&!ũ�95-g����~�/�e��C�+Jv�x&3��R�)^_j M�3mA�_w�Q�v,��S��	�#&��|�<�		CA�7W�(b	�]J�a�36�3P}�y�x�?���_��z� �;���?p�ٌ�3�s��5�o(i�[��{%�A>8͋�B��S��"���!����^����A ��Ӝ_��=*f���1�c\)���\��	���B�2��e��v�`nI:�F�z��@��<b*4�CJFD	&O��;�~6<���8�{^Q���<���~��#0_ld����{j�I��0o�N���/f��J2H5�z�_����'Z�K��f�||�=��8]��'ר!H�^�Q�0��[h
�)�k@)4���0(=��,���l��ґ�w�F}�g=�V�&�1Lw�S�xӈF�[c���)�P7�8���;����s��Sd�	q7ߌ�	�M�d��"Ơn����V��i�3+J��C���TG������W�0n!CA��2>�uԦx�<2�;<l����.�ts���;4Hp_��.ю�ܸ�
F������s��=�����7U��B
8y<x�I� {]�-������sP��>��[�����&I�>���hֹ�M2�7�7	[����i։�W���q:�XX��R3@�~���8G!0��-�eP���OX�ky�gm����%�>����졥�9&�En�_�D�x�R���b����=1�)��^�.R�H�J}��[�Be\5�H��g��),n6V�zd>Sf��I@�1�ﴟ����K\��dqh���0�Ǡ�<Gf���9�@1wS�M�vS��vM�Z;E��籱�F�X�� ZF��>#�J�S'�!z�Y��k�L$ɐ9�2���mm�%�`;�j@Nj�C籩A*ZM[h�G2��>@��R��x7Na4ƙ;�;�.���J�Ԙc,��ktg]�s�@S�:���
��(r��S��aD�#s�!��_��l;n�W�-H��N�f��SFs����p�ŞD�(+*��m����恑m8J$8�J�����
T5�ĘY�!�ty��Z3�+��D��Z�A�'�zơ=ac��"	u�<��0�O*%u��=�Eݿ�h?�5����ڒ8F��:�L0i0{���d�pHa�?�����q8l?���F���#��9�e�8�>b�H-�5�ʡ�f	��=��<+0*����S�>�@'Q�4R���\q<�qV�:��B�|A��զ)�g�!9K�C�������3N 547�G���kȿ�셣�7�y�j�#�"N�M�ѨD�sN��`iy7���V_t;���V��� .L�I�0م��^�3,���Ķ��%w���M/yl�m���.H�gac0��Ǒ]+HKX��*#PR��&m��	�gq�IÍ�. "��E7�����x��l��5rXP�u�l��2U���_]�r^TӁS`�;�,�@Z~��d<&�oj�4��K�[�k����NU��jtd��F׵u~�o��,���I`:uo87ж	t��K�lO��D���,x%4�f�X� �;qxi������G�Dc~�>(��L%Մ)6��~�,��3b����TDF����=�F�w��7�AάPF���h^��:�|�d�Q��*׹q;#�<q�f=٪���
�cr��+�	Ƹ�AQ�	�l]�w���5�2a��pp�mLQ��U�kE��h��jkmo��HI:�|�f�.�_��_��L�l���a��^f��� ���r}T�n�C/�,�skt�.��N_$�e�A
�SQ"��g�S�*����|����̦���.N!r����;j�=����3��R�b���xzP{f3��o���<��Usj�����T�F0QM�;�����L�8��l)��?fs�sJ�ʾ]���y'�����+&u�K����IS0X=�\ꭠ�G��l��J�yl��
o��7���'$�{׼q2e	�|N��(�0G�a5�7��X��dRc��Y�q�Ãhɂ�1](�s��+^	ak2g�-=ݣ��r���
��?��Dn-�ڧ��VW�P%����\G����z�����)��W�ǁ��vY�ӇR��y����
�!�`a1&<&nM%���k���(9
j���k�����U�K]���[���'m�?�@����JAY]�s�?�5���fF�C�X.g�������G
A��%�X�0aG�����z<^���c����{����(����Ur�C��AN@!�F�w�5O:EkL�W��z�5S�)sx���R���C��4)�e�D^���9K)��c�����Cq�Kce�e'P΢�>�	�G�^��( `�V =�0|��@ӁTS�%]u��ӡ�)'+=�T-[��P�\c�؛�%�9��"�8��"$��Φ�h�'e�����]��?+�Ü귱�1�S�;�˒I�=�$�f!��&����{��h@��i��̎�:)�݅U���I��S"��^9S�;s!�*H���(>o�p�g;5$�Jz��V]��{	]¦�t4����+
��b�Clzw4Sx[Zupi���i!Ͼ����г�����o���gmjV�;0=_�*�7�\�H��QXH&�	�_- ���'=���R�)/ʺN豈�-���Y�}P�/���w�K�+��.{�E�9"��Mo_�1�A�A� Xr/��d�~M�ύyۚÇp��Ȑ飂W���^�iC��Z���2�`�k����o7Q�U	֟��)���`����&_=R�(sr^67�h�����)���H���xz��ӓ�1�j���S��;>�"���k��Y��g�4=���i-�^�m�Z�l��>j��g��:f��K�3����� ,]��]����(5S��m�L�~׬�O�ik��sz�+�,U����3�}U��"�����΍�'���L^E��:�'���reO�(��m����H�і�lsV��S�7^w�����.F��Cz��1���	���F=;0�"�L��[=���"��%Z����X�p� �
��t����!v�}vS
�^�2z�.>�5�V"���s����Q��rQ;�_��x;ڹ�G�)���=�8��`a!L󿔡��O��v�X���C� ��B(dLT��Dk�F+�o���W=��M�Hq�j\^����&�(Q$�[�W����o��3(�۵˕�H���D��Eu����F��Έa�aM�ݣH�ypM�ݼ
��p:��s;�3+ 믢W���f���y���R�Y�=�FT��ei]��~G}�����
���L���������`���/�2!�+�Y��KmT�7��ў6��b�fX�,�>7�A,�����L�����ZS./��2��D���u'&e��l4�hz��KY������EqxE�.�W�uE!�=��Wq�n�'j����슱E�QO�"��p%�̎2+��X'��	u
�뵊Qa0���S��gx��<ϑ"+=y�H
J�F��;ޜX�ۜ౬���؋g@Ģ�}�ж�.M��-
�$���y�ځw����z)&	)�MG�~?����PA�h5�!r��`����\$b���I �YD	j�|�K�?5CC�,�N2�ލN ���6��/b<+�'bu�-��H��)�����v�{�DH#���dkqH���,T.ϖ�Oo�8C�|�v�,�V�ĳ��)�Z��{D��+o�5#<NC��-C�A�@ߒ]�ϐ2Ѧ�n6&\/D(e�/���3��@��?7�h����KD�Vo��5%0��%�i��x�
G�ɻ'��]PB$-�Y���2���C����_�Z�#��ǧ\����xpX@��3e��$zP�	�W�L�� B�T�?��\v������^�>-�����m�d)�+(@��f��-��hß��7l�ғ�c;Ayo;�����ꀅ�ތQ|l�~F�
��b}ɱ����U�{(�-�D�<YN�K���LI���Vժ��.�F�T��A?�*#�X��Y�0�I
�yi7�p�?��~Ȕ4Dd��=9b�;��F% 9��2�>�+N��C��>%�5�H��}��ch|��a�P����S���	��~�N3_k)⎨�������)d�l6m�I���)�n��l��s���iܿ]6'�t $Xxn9����ܝ)��x�ēl2��&��Tm���4�kS?ЏC��l���*9�p�,A��؁�[�l���:��Jh3d}9�eI�4~�u�������!��&[��7.v�Ã���L����I<c�ɵe��#�S�xtAh��V��,ב��o������'ӭw� �}��=a�E��;:��l2�E8��j��j�w�s�c˰��ӜX@���E TQ�n"�^�T] �l<,5����P�N�0"mC�{l1�#&�[fumQ�;�\�0�̠b� Q�qy�z7T�9z���8�R��G����{��LO��,PE���Jc2E�R4"cH>�kȀ��ɠ��к�{3¢��@x�2~��`bs|�,v(k�O�Κ���zLa!�H@�=�H^9�O<�О�u��$���yf��Y��4�y^-�G�:_��2�2ŷؾ!�Y&�����#4�V;VP�:Z|�i�G��S#	ɾ#�{�xaL67$��{���8u�y$� �$/\�Vʔ��k`D���F����'���P#��l�#/���E�r�ǒ�$�_���0ڶ��w����&���p�zd��FΠu���԰�]c���m��~nށm��j��E!tQQ{��
ጟ��Q� L��L�@�9��v������Z����E��5{���e��Q��ZEv��I��r2����X VhCF�����ּj^���	�z�i1�b/W�^�sEρ7�SM�<��6jg��XM� t�;Y_���h���\/Ň���0i��"b!�b'B�Js��Dl$mߧ��l���d󛅜~,z�@WV"ѝ��7O$e��Ѐ�]�M�DOūŪ�#<�@.���1	��ͮ6ycƵ[��H��q�G6�=P�� ���KT&�%oH�C�l����OLY�����b�`��B$�ƫ+�'��1�Z7�ŏ�Y���Ox��Վ/�M�>��$�Sal���R��:�b��R�*~�B7W�w'.'��ޔ��o�ƛ���03N�ư%���=1���wVd��z{��-�O4�_j֭����*�s�S;�"w1�Z�԰���Ɍ�����U�1�`�b�̖��C':��tL�4���vv5g�m��å|�sKÔza�N�#h&��3#��\���E�jL���{+�&���W�I'��3��A̷�}�/i�P@�"��q䂰����*7�����8���B��!���x� �I���^�Xԁ��[`�g����$�i�M�
�J��K��`\IEm��ϝ���e-�r"��y� �
�ɛ�!�Md��A��煺*�GmY�A3��9���+U�K��CxP�����&���-Qak6�%(��>�����A?3��ks�j�:�x�2 Fs
�DL/!*�^��7�H]?�$1���{Y"[��1��;v-�	�����h��`�N�ɱ"�������=�c}�7Q�7=:�hc���ڇ�6���[�~�8	<� �?��2��s[�J����71:J�}���
��
~Db�x�9j�A���=�"�����~^��e��54�|�[���w/�c�^N�����.�����63��!ݙ���
&(q`�[��SG��k�^<�q1Qϯc\���j������̠̖�ʗ�d#U��������!6a�������<�W[c��������E����̋F�KT�Ć6D�+/Ӧ�9m���/С�&���a/O}A���8�\�H�8�L��x)q7�Mw���1�`�+�0ׁ����4���,��H�q�W� T�̇2v��1w"3\��v�8�,�����&�g�4�glm�(���
y�"4�%�m�T�W�z�=Um�m�XK9"�?i�fmA=uSFӁ潴�/$��˲A�P�N @7�_�$f�֩:��ȹ�ɥRlWڝr�z=,uj�wj|��:.�t^w��(�>,ޑ/�����Rg͟~)s�A�3^'	vy�yꍀ9mZ�X�iz�Z�9���!�)��S���r�n��no�}Sv�����w<�ǲg���a���r�S�	�񁁫]�j�7�p85wr^����
��"�KJȭ�|a BԐ�j���1)$�"Ĭ��Rv9,�}�{+�K�u���� d<&���1'ӟ���Ox�؁�ä�FPI|�iBb/҃+��&w����=
IfX �%���]��&���wA��)��i��w�Cj�Ρ솬m����e�� gO0�|�Ĉ8cX�i�ld�Cp�L��Oѹg��K|�K}�^�ZY~�!�
�ʏt�a�#��.���ڑ�W�q������'�/G6Ō�g>`�}tx�	��&pl��[�q]�#�\D�D�����rꉘ�7�����1!/��0#h���Gѩ��H�EJl>�|7��!\I^%���܌�eg���{����h^~�T��Q^44��(�h.	��X�������=�ԣ�/f$�m�/!u�ɇ���Y�s�΂��C�Y<.<�jcN%��u�Ht��7k�x����7�g�řE�Y�6
�"�I���-��̜w���5�Sq�gM*r��m�AI�mN���"_�v%Dz�ed::����t��+4��TG�\���p���1�_+�a���%�Zp�5s�H$���4q�n/�+��#E�C�X͓�����$�Ok�|c>L��M�0��W�1ٻ�Y�����d}X�hb�I�����Z��&�<;�������U��5,�t����E�"瑗�΢�:�C1 �� ���ӗӧb��	p�ϖ	tq � ��أ5ÑJ�ٷ���c8�W+y��O�&��!js|�د��G�๔��HL����cLKsQ}N�Ja��vq�C2D�6��(hy4 �99%��+�ckm#�5S
H����Om�;��7�Þ��tg=ZL?ه�ې�����dj����[��.�Bx9Nn4�P�N6�#�~N��c��F��G�G�Z�V7��<�"����c9��^E u�Q�ݝ"NT�����3�8,��K Jh�;jy0���ѥ�>�K�����3Un�	�LP�Á̞�P3&�7�L�n`?:Ӆo.�������v3��ĳ�Vv�#���H�e=�%{O�@�_N���� H�6c�S�X���?|�]A4�[�
XE����r��������*{��Y�g	����A�ro�s������\�k�iq�9�UӜ)�"�Y�O����Ķ��Ʈ�pc)_�x8{�H2�t��K R$=03a)8r�x�6���9ML�ɹ$���q�Q�y���f*;���a��]Y���s�*�]�NH.~:��or���L%�����~�j�]ɼ�����ߒ7{�E�Tb�q���
�*���(jƪ���EiI|)���)�d�2ҷ����/��F)f����T����Z�[���5X�+�E�EQ�w���I���ӲrM&%NYIz�[��Tg$�ǉVHMe��eJr�74������|B���#�vI�/D����� ���F�Ct�
FB�-qr���N0�b�3.�Ώ���t+���땫��ؐ��u���fK��,�@Nm����@�г-��	���;�]b%��j�6��C�ss&�<z��ي=A�f�R�9S�CHIO+�	5S�`I��:>"��"��F�����Lפ��W�Mh?kq
A�U�	A�:�(�`��	����ۖ�8"��@i5��f�b�0��mh�kԛ�Ũt|�nĄ�sqD�W��Ij_�HtY����;2`��4̅��I��@�^�0��ɦgP�!�YK��P}�����d������;�rr�n���;���#�c:5�nH|��1�^C8<v��bev�l�{#�lܨ���:�n��s�D��n�N��}�� ���1�/��@�{�l�/��>�Y'��R3�m%����X3Nd@wL,"�xm' ?���nͭy��3���x$��"��s�' �����X��g�����ҚO�W7A]5�Z(`��nP��l�Z�7��v������{��)�m܂�[b�;A��;l��FZBzԆ�L�6WL.�X#�pnT}��y1p��r*�� ��\�IV�4f��W+���+~��A$�ja�9���1es�~��)a�EP2y��恮H(ǮFq,�`����N�����7z��'����(�����cs(q���oh�s W�T;��2��5��k��{��N���'|qK�m���	!����|�^X*��T��z�уu\wƲ~_�b��W�x����Q�%A��z�_[��f{׵�݀Xc(�p����:�R�/)��ؗ>��3�=?̵���.�"M�#���ľ������㉗��s��Gb��{����� ��o��ʡ ǅ�+H����L��o� ��n��ndb���2�����ƿxD�zvV��Z�9�M�����$\��NX��ߏm���q����\wV�����K��eC�ʒ�Z��HK�A%0�x��{R�����,����m�I�i�	F3>�J
(������w~�I�G�l}4n���z�1�	�G�AƘ������x4:7̑[4���	��|��|��!��dO���� �
`��:F�`�Ԝ#��7��t`�y�˙�Ǵju"�;x��dWV/b�yN5�����u���ML:�[`6�����4������/������7�g�=�?�/�J�?�T��	H���s�6S�$����b��R�����j� K�[�ٯ��*8|2u��7�'Z�hw]��U�l5^$fSBQ��u3����)I�+���E�}7pw��@�}+}\\y�Y��I*��5lLԳ�TǸ�r�� 5{�۫�|�Q����E`�_�}��o�a\y���`�e�ր@!};�;yS�����Dr�����0��W� aq�zQ*^�7�rh�����S\�L�Rt��G��DŮ����j�~ǆ�0�$O���2�g�0�6��P<+���K�)���b>�@���<4D�G>�P�>�I��W7B�q���g&$�>
Kǃ_��lv<ͫ��>�PhTh�Ѱ���݃�7�����8�#maV;ch,bRG˭2����k�}o}_Ֆ�FDg��-]3Ja4Q:6��E�S8e��'�� �����X/9�wϠ:J�I�Uz,��r��cۭy��,څ링L�g0` �q)���}$�*3���~�,��Z8�[dc�b��ʨ�{y��#<)��U.�,�(ҥ}W�"�Z�Q�}�|V�'z.u�%�O�XϺ��)�I��!�*ɲ��K5��� �I��X���� }��ה�a��s��0�,�IO5��ddڧ%7���pB5
����gH9J;}5��?zΖb=��� K��ݨ ���y���/���GQ��;����1�!Y�UP���F�2��@d2i��}��@��I��-E�,�S�	�qXL4�_f~jv��$^2njQZ��|��nQ����괎�{�u�ro�������!XR>�GP��Q��vZן�[,Y#����:~��QT���k�m������f|��\�f��o� J}��j��T��i���5��k��U��}���^d���
��q���[k�|)�g�-pLq������
���ضss�n:0ny�ᘻ����[�������?*[(G85��ח�c��Z>H�m�84��Q5ϟ`�um��E��ێ�Y�����O�4�1�j�.��' ɠE�����Y�]�7G:���^)��E�]�Rsi����3[YȩҘ���$*�[������7��a׹���+P�d��!�y�Xa�V���1��I��cI	%0K��e�{�JSf5��
즫 C
n�PZ�;{�@4r,p���s��1BT��:aݭ�SM�Y��I3C��6|a�\��u7���zk��l��=ă���3���.P�����,cc�0���6�����H��k�i|.���uFx(l&1�ߟ(��GWf��
���ndeS�Ҟ�QUL��guSD+� _��,h A���H��8;�K�7����P��lT0��#ĩy���9�
U���Tgs`�L�|B�u9[���(4'�!��Ӌ�ۮ{)��k�lJ�#����w݃7o�؎KW����*�Xɖ�9���{��^5ޞ��(󖓗��x�[7N��dؙ�@\�Y����N�n�Z�WLjn@'�V��6v���T'B�2����ܫ��/L�� �@aP�e��W�3e�(���4�+��Rj�>��6�'�@�~ #+|H�SgE�#�ɥK�i�@�8{,%��H$��@i�悋����Ty1u#�ߎ4Q ���c�'�d�gϫ��q�L�[+/�/�ɵ.tF��)�D������^��Gz���&�S1!������҇q؆��P�ݪ�U0�1�~k��LR�<Lu.�ҹ5�ʶ��~\3��jΟ� �Q_t��{�� p�{)��� �x�B�T������M�[}��p�E�B��@[|����EW�ཏ8W苖?�\��7?�)��I���7`�OA.*(ez����N?�@|Nbu>���x�>�me/��,/յ�6g��0Z���LJ͕�LA��n�1f�X�u� �̊ʊ�`��������PS*�#j(���E]�� X%������~�x[�C�w[^1��jy�$�SiE� �NV�Ȧ��rQ����sF���3��(�+�9[�:��M�����ꅍ���jV�Sp��SK9N/Q��bn��Yh2V�3oO�o��j����Gp�ChuTB�[�X�W���0���Y݇���)CJ3yK]�˖0=�����@ٍ����J�~W�pEsS}�N�|ht�-��P��Ei=&������;���.e�K8L�	@����,2� ����	=B��=>�wS��V?o�x�gkZ�?�m�,�'�ZAT��P�'�hѫ�C������<P��e
|.�n���Va�I1��l��W�x%�<ŕ����(f��u�P�h�{�'�yՕ*1�rY�z �=�-J�
|�K��gd���7��z�c��%a;� ���:�����₈�����@���e[������˦�` �R۱$������ܳ	,�� ����&it���#
]5��V��Ԑ��C�p����(_k��hM�.VO/�� ND[��%������kS�2A�w�_u��e����Ë��7��$���G�9�0��<g0U$�<��{�q	���D�����
`/?������>�4`s�Z�����[��VE���9g>8����B��g8���|�>Oh��k��]t��Jq��X�+.��FO��8&��m\3c�¹�s���%��R��W8Y�'z�w�Mov/Og��ӏ������i����K\��4tS{�~y��ʡG�<Qr{a,�П�x�v�f���d�R�>���Y�"��_J�� b{�3 ���O� "[�����=EQR*�Μ�%��k��E�B+�o�i}�P@�)��Z�ߢ��Bͫ\Vs��a��%t ���k�7w|.���u'?�k��ߚ��KI
��lR�Ǖ��c���,!�F&s��b�F$�㑬�L���F��;�ۺ�$e�^ɼ,�w;�1pB� ��*ym�,�1�_�����w��A��I|jx�ON/A�����Q,z��ɫo��3�Jp^wvL� Bj�{@s�ݮwlQ5��<�x���~n�!�I-#� Yb���?-~�����dj����2	�0q�VF�����Q�e{4< v�p5蠕}K*F9�d��`(��:�� ���Rd���3�C�0?_+p'����_3���N]al	�?��NV�-������+��ZA��CQ&������:&JĔ���
A��:z� �#���ӡw<������H�d��i1=���8�O"		�l�'ā� ],R,3<�r'�I^����+pQJ`i��sXdq:Pz�^�?Da�
�.��7�F>#�n���!t�<�ٸ(�[�2Ք�w�� �X�B>=�T*T{{���LU)_��
�5n�S���;�vD���΍}6�e^'8�@D`^�yG��A�?Q�|�k�� H*RA�-�#V̊	@T��Q7g����U�̇����*�(}6����@׮��
��2/��fcX�)Gv%֨(���r�6�VJ��y7EI���QV�������Z4���W�*��k/�N/�d�|5�L-'~w C����̇8�WE��~(��^��	����_�x��]C�O!������yJ��-��҅��\m���x!����]���ݘ�(�4<�����d�jLŖۡ��X��s\|��clF&�4;�7EK���@����e\�^��$�+��6�P�����S4yOԞ�	?Zw��� 2�����a��1�"��=<��&A˵����wR�-�L�� P=����8��a�7J���+��n� "F2z��;o��S�ό@W�E?�(��k$Y�t��]ɥ	�wP-�a]%�6B�����yq'}�A�����Xm�O����dxq�����w���w��\S�}6�Ռsn�Ww����fދzQ�(�1d;+UH�+��D-��Qr�Okde����M�t%��/,���ƶ@8�4�����ES�ԝe�x@�F��st���R\��=v�KZc*T~��W!|+��t��yYf���	=i�ňu�o#�*D7�PJ,�HVNwR�^�����A��K9���c7��OJ����/OTs��r7�	��%F�T*zVLhIS�ޢ_1N��n�{OE#,���2l��|��d�R5��8h��� +Jz��*�^��e��e	���c�i�i���}�4^V���4�@��%7��S�t�B�L�P����BWYA�+[�����D�_ӫ�sQ?k���J�MT�����Z��A�d�Y3u�3�\��͈/��T#YR"߅_T�^��Yd.~���7)�ݥE�9��m�y�
�E��ҋ
.�o�R�-aVzt�di�m�֩���hѢ���Dl��KJ�7B�ߑ���o}u�����w��5�=B�	e�������|�>���O�1^ޱ�UD7p �d�?�Ya�/���s���8:ڈѼ{w	ª��6�m�x�>6X�fF�Y	D��l��	[=W��7�u;�'	7�'E�`�
�?�e���V�J�~Ap+<�D����п��l/�G̷��m���XCi���C�P���&��	�ӄ��a�#��O��>�}Ȧ7���v[rU��EŃ0�<gW�IV���M����D�s�w�4�0i�J�ǅT��Yq�Ð,��&�$�`�;A��;��j�*f�M�i�{���b������v"ȋ,��;���5������Zl0���Jk�W����W����o�&7oZ �f唸�y2AS�'����GaV}�NMI>Ɏ�>��I�|��<���
^����<N��
�~�"��J�<���e�2����L̬PB��PV��j��䌭�7L#9�L��`xw�d,��}lbdW?ݤ������iH�����fh�udUL(G=�wo�h�l2�l������?�H或��Uk��	c���6��0u1/���G��E�g���������t�a��U���3��C�����2Ŏ@p}t����Dؤ�9��c^z���S��i�f��C��r�(�0[�w<�ya+�	��,�� �$�'�[��ds�ďl���/�{��`BݦKU�ֽz?���U8��y���[�g��^����B���@��#R��D� 1���T<�<�VZ�ߚi*É��\*0D�=&;��B9
<\1�,[�ûq�g���n��n<9��^�YR�V��{o��z��W���tс������k
uL`|�2��V��&�:KSc�M$0?�B�$�u&!p-cn�U�|ȠZGN��sҢ�,xa�}��[�0�Ԁ��3��vk0t��oѢ�y��=��R�����"�G���?�S�yh���A�|Z/z9�$�3�Ь��)N[��=͓�*����z"t��q:6CI����s� [�����()N}�!�؄�Zg������O
u�x���*�tF�WLS�y�����97���:R��P��,�M'sL�
_ gzx0>r����x���]W��X�e����QN�jn���9��Nm��mD:�N�C����3-���7�Wq����r_[V�C���l8�Yx��Y��x���Gǡ�f�BD�_~�"��ʐ�'w;���BD$�C<Z��?���8ɯ�po�w=(#J g�`��� %�q����^�� 'IZ�ZZa吤���wn�����������ھ2Jf��Yy�*�|ȣjK�S"���Oiv��ǜI��R!yuD>�\��o��C���|5��%�����mk9�t�����.������|G����'�|6�6]/ݣ�AG�I�6?N!{��������."+�o.�f��DX�J/���6��y�����3�[5y��k�3�s�%o�u �����7�!5}d�(�IM��F�5=�m{pU�"IE Tl�[b� df��N�V[V�z	�� ܒ�#3g�ΰjuw���R���&����6IsF�Q%���l�mJ�)��5UO����y�Ld�C�����5�` �>ڥ��B�JH�v�na�e�S#�X	/!� 	�[�p�{f�fk d�� ���\���7�>ސ�2*�% hYw�4���ǫD��Zp�gHw��2�϶MLW�q�,�8~[�������yg�+b�]%� Z.CG�3����ͳ��A�Xz��9/�E�ub��d>�(~�Ѹ�ѹ~0Y:�@��7��f��d<7�6��MB�I���7���Qu���k�qr�$pXi4��u���~L�[���C���ޭ��DW�-P!	��SB�ࢲA��&����3�=�i�3�E����6�O�,����(	$A�VP�}��������[�.*�x��L���|��T�yb��t��$�0�=Y#S�Z��WӔu��p�n�0���x�y��J���0{Tw�Y��1c��^<����V��B��+�#Ƹ����D��K9��y�#��Ѣ���5����0���l�P�@��	s�]/coJj�|���4vDCMI�+ʳ�{�<e�jB:�/�&g�eEo�X22��c�<=V!�ߛ5���R�����S�z�>~�ڴ���څl�Nė�_�#"7.p�Iy�꧹"��z�6BT�a��L&�ɉ`�?�ZZ�d7&�(������ׯ���iKأ�346�&�b��YUGlrg�����ͧ-luM����Op�L�_�����#�r���N������������`uqnY�h]��\i�V��a9��/S���{04jMN)��	�j	���`6����E��+,�H��gh�?e�64t[�-Ǟ#��"������´<�β���^�n���͍�)�L��Q�Ν��"�QX;���4�O� @Q��1`�0b��g 4�������t|���3���(D�>�(mp����k\�.#�q|C<�{����;)Hb7��/�K����5T�l`U�9�������1�I��
��O�$#M��MKn�YT:|z��[�(��iy^!|*�C����;բ�XZo�����i�粠.!�uN�w�S��+�I^W
\WQD�oW��F)Is�m�A�[if;=����e��)+eߊ���z��績��+;M���g�Ϣ�[��7�c�_/��A�v#[h�;���!�(ʁ �V��R���Q���!V���`���(�d���v.G0�ǪY%gd���� ���ĭ�e ��#k�j�p�ߕK^}r�IG�]�"Ę/o����=X��{�MPH���q��XzSS)�t/�]�|ꃱ�ec������#79�V�I�;���5@8<ʾ���c���t�9������Bx�r�X�E�a�|���Qb%�}�J�3��By)?�H��=D�w��&(�v*b��wv��i;W #�m ��qbZ��/I�+�\���^X�xV�?G�.ΥN�*qŝ�����D�/|��GD)E�a�!�P��u�C��b�y��DX��f�'�mڢ�Ϩ���os��qw�b�Krp��EW!VC��
�k
�5S�P"KmPۑ�����Ɏ)y�Z��dD'cr���9_��l�h��y���8��f���}`�]d�jo**+5���*���Y<Tw�Il�������3��sT��yUV��c���t�I���x�o��dKf��Ҧ�w>��ǣ���[VX��c�jf#�5�A���"�k��:��;%ź�5>���zq�-��t�`�/��`��
}�4�ETk�sb&�C��T��U�㤴�7n]������I����e�&��w=������7�8��-�b��E;�%����v�A�TI�0���F��\d[�H�߳������Rp����0.���[S���]�Aa��E-���N�x�V�7���R܉c;[��y~�>�㳧�>6�M����'��(@F��
�lP�J�\�)�QJr�B�' �-�)���z�(�	���,�z�C����ae D>�K��4hm�V��v�Fpr�R�4����*�f��W���Y��V���)��u/���Y�~2��z�B�L
GɸVr�Ν!��IeQ���"݉I>�¬k
���C��T�.t���ۇ�z���V�4��{uh��P1�J0tm9�q��//xm�g'%�� 7'ln�V����F�~+6��]pwgS��QZ"�~}�d�H&�i��@�shL;�\a:q�Bk��f�\̻�RB�/�o�&�wx:f�2	�s�!:���r����ZQ��!�����"�K�E���-��%��QA�A�i��j�N���~�H�}KIڜ,K��@]8s�"���%�w�>'ȿ�H�+bJ�b�'�c2,�#6
 Fe2��x�d �`#�Mq�H�]{.��p���l4fO���I?��EΨI�M�
��1! ��ѧJ>�|m$y�v8�B�E�r�>"�µ6��Լd���5^t�����{�,��W�NvϿ���Zg���5��s�r�ic+S+n�Rc_ �����5T1�x���Ѓ�2�����Jv��э��G�cO�RHS�1�N�OTŭ�-Q�5�gQ��P�k�:B��K�xp*gtz�$� t�,Q�S���m��E73
���7��BIH�ߎ6�*�eE�� ������G4�A��c~���nߡQ�է^;��a���|[	���z�9r*C:�o��q�i�Q|q$7����>��ǜ(�.q���] ��N���FƩ��mf�n���1�����aa�/��^z���,Y�U��%=+��ѣ�	�Z�P��3(�ǂա� @� }���j�h��T����O�Y�ݪxB�������'V�ؔU/�D�̺��w��hԗ$��"�$𾌽��=�  +2_O���`=���@���p��+�ˊ�[T.N�{	�3s;3�e���'�`���A�ؙ�}���p��o8�IY!�Ƒ��,���=?�rM����;=�����%�8���(]�8EX���A �9AկƉ�tę[k
��y���w�U�D�:������5$�w'�	b�ѧ�NG�O{�h'�H:9��#%����yD�`|�pe�������/4?��Ҁ�����:�7"�W�Q�W�{����Pڪ�
��5vT�=j��|G����hU������[��Η��k������z՚�7��՝��2�R�WqA���f���@�'�/�.��T�jO�֮�-+�A�|����B3dQ>��_~��0�G߲`��9޴�^������_N[r��l1W*6����_6.� �C7{p�^�p� 	�L�# f`�5�4���Lp9��a�0z��m�0�l!.�}��ꕣ���ШD��JT:j��⼓��	�V�Xe�Bv����Xi ����D�m�3�Ү��U��~�ꛔy������(eM-��2Q��7N?kJ�l�&i��IT�4��_o��|vU��;c��鞞>uy�?����'k{�]���~d�\6�-6�	V˵�̿�L�.�y��E/�8C'겜}�Q�ޟ8���GX�ՔJ����%`�iz��tiY�>xX��3L2Uռ �����zEr&�o���E��m�H+|��'����K2�ɝ�J�t.�sQ#�NH����v4�X���&����d2���v�������\%��F!R3V{�H���W/
cB�&C�W	M�Q�P Xi��5�r���X+_7eЏ0���O�CI�.����"�ܗ���o��ѻ ^pL��!IBbe�<8`�rz���W&UTz����ef�Yl�̧S����F�:�~/rI����W�Lk-�ʻ��0�?SV�m7!� L��ɡ��)���)��4��`�"�fj���"+,]~�X����� PļY�z����q	��9����߃F��lT��[��A^?�Q1�Xz/��M����IsV£�C���[O+M\
B�n���n���(f�j���v,�aro��q����r��A���'Y�d_E�8����Э{��ݲ���Ĳ��0�p�������|f �>d�[	�����i�;���5k2�!�5l�`H(�J����ؓ9E#�L��6��r���F���\4�p�.Z^ދ($��@Z@�	��<�a��e��,@ϩ��*�@��F�f��I�OM{?�`�ݙA�y��Ó܍�&֢�΅�-f;��6��7��1m�o�v�pV�2��Va�,.��<y��P%[����j��,EFEfP�(֒���;#����|�Q݉ςݘk�+�*ytm�^7�͍�:���ץ�nk��f��s�ںZ�n{_c8Q��d��ɯZQ�"��<�v>a��O�<��p��^���1�lt?X�s�r��Ro�R�R��>g%M�W���R����m�
��
��D�b������2��&%#��x7�n�Á�0u�I�;��O�^%4��g�r�W����f��u��׵���\%�>䑞Ρ�-��qe�"ӐyL:7�C����]�Su?z��՟M������N֝o�V�b�0l-Z�<YE���p#��������-QW:|��D�E��֣�Ox�T�^��y^Չu�ϖ4l����i
.��w�4��y���P���Y��%�ke���v3t����I�_0<9�6����W�G���YP���%9�T��x��5�Oж$�p�w�r��d��Q{�ƙʄ�^L�]kA���Vx��3���/{�:�Ɋ����c �z�Y#0��{;X�l��Iwd�Iȇy���������#���)�s(��e)%�[�<�}��׆�KH���;�2���؇X�X���!�Srn�IxXVy��B|�t�;�x<
��Mrܥ��-M��sZ@�t$�NY�pWj�*����oa���o�<H�≃h�7b\	�N���omp�����8�!vJ'��ɱnbͺ@Nf�zf�1	6���/%�YN�*��z�<���e�H��Ik,����@��0�ɋ5ş�//ѷ�7m�a�ؚ�B5v�OS9� h��j�d< �t��be�W�ږh�48�K�A;�q��
B(j��{�b��9���q�}/d�����AĒ��;r��mN	�刲��7�}l��~;0׸��'0��5�~i�H<U- p������$��K�`�a�0!YBS����:�J_��C��V���ޘA�
y1�Dh�#�M�bَ�I��u��������|�� ��*幠����KR�Z�:>E:�~��9�n����2�8N,�=��qd�6 J��:�Y{ְ���ou%�Vκ�t�Z���R�]
=l��s��%�o�%���,�-�l��1a��es�e�Bᇆt6S�Ss`_������?+η=K��<��7�U�Baw�Yg��-���C�6�\�cy~W`�`�$��t�R�|Y�i8Z5N*��`�,{Bΐ�#T��Q���a��(�!s�_i��ةK���ac�CI!H!x[$<�6��*�?q`��@ZK���㢺hiG%h�k=��89d���1�Gg ���x8d��ɝ���G�?E	�ۍ�@dU�U���7���a\�n�t��\�O�:k�H.�;Y8xL�$:S�w}{�X��E�~� �����xQ@6��bNԄx�C�Q�m	ۉ����?���ߗ@5*��-s�dU�,݉y���`d1��&M׍wu�ӈ �[���@qߏ�t<>b. �[D��i��P�x�х*�L��	�Dl�����c}Ei�&�]��_M�DҒb �����Z�+�/o� E�ͮ��@0�W�>9�h��'C���a�V��&0I���P��'���΍_��;��,��-��*K���2�?��������+�ϼe�uɔ��$Wɓ�����;�������$���l�D��#�b ��oՓ�l~CG
��txW�N�b�r�7.����l���="C�ZD��^L���2�����]ɏ�a�AO�b�rQ�U�,����@F���Y#�}���C�K�m�T[�5�. �
���ODY灡YF�:�0�=�D��_���TVY)���E(�W,�Wt1�t�9>�^]4�\Q���*ρ�b�(VK���k9�w�@�	�%/Y��AՈ���ȭ��{	����U9�Y7�8/š��VNG���d'ά���� nl����w�mii,RE7�pR~�v�	�H�����Eȅ�x7����+<��9ׂ$�n������&�_�$�C��'���Mq��H����s4�A���˄���>���M�	��j������������/[mL�A�սԪ��r�vK"ij)�Xƌv_�5�$o [�צu��\I.���h�,F�u?ڤ��	5���'��NIm7?#�ưe�u؄��k��Ǿ-:��fN%[Q�u�j��u!�@d��/R��ZL����_Y���ӊ��5*����uv_��&/	['�8�?�lߡ�	S� ������C��������"b��;��Ȏ�ɫ!�=���Z��C���$�^�$=�E�Pr¹�q�)��	��Gt��N�ݯqd�=@;%R�N���rR�A`�p��T�p,�7Q:�~]GT�:���Qq��l��Ďs��$<�<z�Sa:����`��a�0�F�}E���	�x������ىv6�W��rBƄ���O�@s���>}��t��7�S{^F�� �{k���t�syaI�|�μM�A"�g�����,Xxa�;��$�WL��dᛛ�3�l.}�G�����J��i=�7���/MK�*��x�ꀚ%F����bB5π��B&���6���S[��D��QvU�Zv�J�RU�s-�M�(�������z+��:�}?��ҧ�E���W�G�Fr	5w:t�o��[8�?��B��""Jl��A��"N���Ƃh^��U������9�!�g����f���a����#9���.���:��3}JK�{3o��=�U!?�T	���4���f�(:�L������h���헒�Ѩ���p�X;�����P�3(^��Xd
1�&G8�B��m��	m�G�
���	?� Q����7�c��P]��+��~���)R����;	/�Ah�I�$��|��w�� }~�ǭ�e�&��'�U�-���U�>K��s�(n���+�Mˈ�IuH�����|��]��V�g*"�3��0�r>j�7�p��3E�@�C�����i�+�A<��Tx���YVԜ_��~~(�
�����D��;�>�(�2]'��e��*3;G�S}<;[��Yz�nX�"�_���V��cf�ҥ�6����t��$"Ą����`���Ztb>�zl�+36O
K�4���E?��2]��EG5����e^�$ǅ��9����Yi�*���v'�+$Q �ƻ��Y�YaC��^V�K��r���-S��2��Mvq�f�V~�5��]����K��(��6�P[>�6O�������e�Q��aSOē�V�;�gg�7.����UDz~u�}�+Dou�P��m��;���|sCj�F�Bj2�b����%��g|���F݋�~������Pv��f���O;j�(4�=8��N�q���I�b���x��;T�WG����T�n/��PC��U|���׺����_y"�F��5��o?�foە~X�>Շ���l���gc1«���!\�b�mSlv�j��q4!-}��͋�⺳�t�����Ȣ�|q�O���:��M�jv����%Ҵ�.Yx S���l�'T�nb}d�����wӻ�8).O_�`�1����ِ��O�׶Z��hN9
������s�9�T��`�= �Nyf���un��L���1���D�Dt�n3pq���Y�`0�y=��<I���yp���g�j�C�XEb
]e{�.;Y���Z�ñ}a����E+�[ U��ࡹa&��D6�)p�M�eU�2�������>zփ� a�'W���!��֬h�!��x���ۚ0�	��BAT�@��#jogGaҹ���g���`�z`Q�Mv��]];�?�;f������U3W_ 6�"lCw8�hm��똂Cǡ"���. �����Y5��h��G|��_��O,�>wM�2L��V?��i��PA�K/}���i�׈_F6�z��Z�P��r=���^�z��R��A�Yt������fa������WH��Ekה�0Dp�7����/���HQ�W���⤷�Dɼ�f�¡���b�cfX�-<��,>�s3������X��Lyп��\��&�t�$�q@��<�Z*�O�eh�j²�[5���ڂ��a�Y�z�S���t���5�����R�g���,�Y-X� �6!<z5��,��J�����P���� t�&�Jp���lG 
��A3�J���}�-������!i <Fd�� �=J��/���#̧^�V�B���4��&��"$��F��o& ];��*�t�tB��*���<i�6�;�M� ���?z�/��tN	ޙ�M�Aѐ����W���ia�}'��ő@��2*nvwf�n(9侂3r��W���f�B�	�sv	��Ur�s����?c�rЙm���@;�uT��t�:_�A���e�R�B�5:"� C�VǊ[����U1�D���
��;j����I��xo�I쵺��ܫ>�U3+|;"�9��Y߫�3¸,t���.�tj}9њ��t0��P�/oR��43��s�
���ʩn�����.u���ɱ6����ƅ���p����j���Ǉ�}͟8Q5���Lu���U,��C�硅�g�3�Ο5�NRI���?xk�ϳҢdH����G��7����-U-�m��l�y�3]�V��Z�K��//��x������&�ï����՞+��n*���H��+��W�/D�V��!�y'k W�|R5X���]C���}X���6z�`@8N�B��c�<��P��n��ŋW���I����3��|tdId��������ص�4�'�`��H���'�'��$���k��Y�PV�{<�^��Mi�l�Z�2B]�)\�%������UE��5Y;�C��-[��x=&�z~�x4�������zx�����>ޡ�m�E�i�\x\p�`�JM0��3Z	$O�`�����T'��+��z���>�#��V8���졋����H}\T���D���L��h��}?���+�B��>�UК���>8�V��U�A�k�0���u�:sb� �$��rU��o�4
^"2u���5ө�#hF�@61��T���wꎑ$^�N�!�	5��#���|��M�h+�Ε�c�f���y
����o�;m�&��c"6�!�'�۲��T�N�,� G�=<�=ki�<��9�����G#wo�~O��O~Gm�H,��
����ޤ�/ZwR����Yf<�9�QvWQ)�����o^!�c����&B�뫱4��Xf���O�^ϥ�����*	έ�+M��po�	�[AX�m��J]
�A��
y|8�����LQ_K�g�����ߡ��U��F��_P6�b�<��ML��t�,�㔼f�wg�fGZ�# �ji�/���t�/����B��	"EHT�J��b�2�ƇƑ�=~�8D�;ŜZk�Z�����R��e�*X��A⺊�L6�'d�@�E��9���
��&cg?��Т�#��Qb�+|�5�o�쇸�N{O�@���_,�x��<�!�zF���1�M�k��L�@�jB�(��h��b�J h�����D����v�#y��T @�ԉսA�@�����T�Sv�+=�^�ۨa�Ӊ�\芢�&V�$J!���D�,nj�j������%�J�	0i��/'t�mF��h�i�N/!�o{!s�d��TNP=J�7Qo�l��֫BU�V�!��N����_���ދt�����$�<l��f�[����I��V�>��ڛ�(.;Z?�!0A����#6�#�r2i@�R-J6LeC5-�I+1L��W{��E	�YT2�{Q�|q�-_�#1�U�:&]�==Jcp?^�c\@�ͷ������_؍:���	��!M���g��0Whi��"�����b�e�*r�����mmv��4���~�7W��,���<)�L��8i�M�8A���\��,�s��鉃�W�$݄7[|[�C�W�S4Gѯ_�g�OΫ�
�Ss \�Ŭa�����z=�(ۚO�6ǖ��Gn�TG���1W��1���;�곾�`m�
x�z��]�c9�v`�τ7U��38zK�A�C=Hi���{��1���
�VKU;wd�Q�[��i�-�L�H�痓1������.�5u��F�ِ3;�Lx%��A�Z�Kk�� �M&��l](z��~��˗�:[�Z��B��~.`ǋ`w��q������z��<W��ؘ�*))�<�J�0Y,��������Z����Q!(g�]�ql��x��W?���Q?a`�+���nՃw��&C�@��v��߁�鿤e=C*���|�w�ȢG��S6�s��;�+�,�Ze�ح&,�t�в[K�bg���&:C���}��H.I������֒�J okȐ�&�0���CJ����hQI��H-_�,�O5*�[����O)G		x3��3���>Q�% ���<���3�`��<� GB�8��F�r����{��y@���VxFԨ֠��m~��
a/���U�ψg�]�m�߹��+�fK��}e��G7����av�����T����v;q6�E\F�-a"V����ZJn)v2œ���'�u�����U�3����[w�T��wr�ŧ���24��X)���z䣘j.��{����|u��yAÁ�U��mkλ�`���Ś���y�%9�ַp�*&W0��k\V�9`��q�r��� ���/ƯSl��I1��ľ��r������s��F��T&S��.��x�@xb��=�:C#K�lϸ	`{qb(�i�[r�*`F��Ge��3�����|�I��Y3��1E�R������C�x0��y>Pj�qb �Ub�B�'}d������z�A�[}�R꧟�1��Y+�����/:utdP��� �!{5�"����=Y{&s�s�BY��[u��Y�c����t�}O �� ��K��'���f��ý*�� ?Gx������C.��w�Жw�ະ�<P�o�Y���R	#}4�\���k��#F�1�x�E�S 4ճ��R#w [Ci�`���xߤ�퐷(��|�$@9������zA�y7�J}�NF, u��jq�r�7���Ld�m����f���x{��g�_2��l����/zq,i���P_o3�?�p�.~ump*�k��7[�e���ܙx���~���@�S�/�Yp��Y���!�����]uh�S~ ����OH�ؽ�Tx�R�w����p]�K/G���s�7��B.UVc���z5?dxOz[�}�0%ZykYI���[-��*P����V��C�������Պ��V���UX������� �*��k+�'ha� �X�u3h@L3����P"��_���)�2��{�i��5�l��x	�q��da��5��L}���8i+_VǬl�}$�Wh�8Mn����t�W���Xɚ����c pkv����c����9�UK�?�$�_C:N���H�Z�ׄ����$�&�ۀ�n���	�mֳ�㲐�ۂҹ�eVV,Q�;Ia��T�)۰��rَ<�/ hD�ǵ�6r̜����Rrkވ�����[,.���a>5A�HM{c�(�Z�X�q���T���,���j_� K��};���(8��4�s�������k�n>�I��9*,�#F�Z���������! vl	+���m)W��HY�O������i<���W��w=���Y�͕�2�����U,��Z��l18��N���7�F�m��>3���T�[��`��GZLZY'�4�E�у���:�����9��v������Oq�a7���zӪM��}b� ��E0	���I��R(����#�Ӗ�|����7��ڱY��9?�pB�b��7�m9��!�)iD���T�-�Ȯ)�������&8D�Qi�u�ЦTv�J��YCZL"�dCT�Ox-�@�n0����cVy���X�V�In����?<yKYbUW�\h���8i���|��a�\�/� k��V���Ԡ�[����|�s	j� �8��CjVmU'u�&��OG���I4����C�}-�Q��ވm�j��!�$�[+�����X�g]��Ʀ�ZL>�b��`DD�b%U{�}��7{}�b�_]�'��oL�n����oQw��Fn���A)��?���Lo���Iq�A���/E�D�IT ^�S�Cm��Y���v�zl�u ��܋�_%��!9FWy/��b ��ss�s�����Ly��NLlM��~3L�pp��l�lo:Ydv&D�Ǌ*�ѹ|;@NȇR�e�c3��*�y�UU��_�(�X��L�M�U�N��h/�9d���Ѣ�F֕�w΃I�ҧK�r`rVJ_�e3���"&�F�F�Э�4=R��Fx:��T�AX|߇$%�za�~��S!�Q�L/lp�B5�=���I����6a�\����#��h���<�o�''��{b�W�jfm0���KgG����RaT+W��D��<v���h�E���F���L�E:$0o����c���������B��C'�^3�;N}G9&u�$�o,H��-��EL��m�㢳H/�E�����V�Ԏ���7։H����^�#x�˪��R�k_:㨩l�7�*�D��ⅫE3�`u��ܺ�Y�
���� F�"DLfTGA��L�������//�I�WKΩv��U�e�#4A��y���=S���?���0�f@7���n�$Xt�=�w�Q<߆+d��1�ֹ�b�il1��){EE�^�f�0-�����-,p>�Z��mh��QBX1�0��yZ쁀� ~p�,	�8��"ƟE�p����-����Fd%3�lWU�rHJ���m:/��Z��Jw��y:����=�?Z�@������g=�b��g�]�����I砭���>��I�fڽ�-+|�GS�9�QF�ZoS�d���$Q��\�&^�m�C�������vH���3���n��dr4��F���Y�����E����������h��|t�XH˚����fI�"y�|�Z��@�J��Oܢ�w��F���%��w)�G�/Vc�V	���j������9����|"�l��0s���1�ģ�m1�qO�!��qrd�
88�%�ϚR,wS<<�z�!	�
+m��i�.\��60�'���$#`���'�u�er��qsJh@g��G�[��:�>�b�i��V�[U�\f��[-<Ǜ׀@2��Ӝ��l�uR�
S��#J�C���V|��ߘ������M?3��[� ̝�Iz��[�Q�%A�����z6����}��4���]l"s��	�۴ρ�u�X�q)�H��C욻uVu��\^�ff�a���,W�ߗU�T�V�I7��:�a�B�&�%��B����.�ׂM���������(C����{<��i��҃�NG����9�g�|�L�mdA�~[�e�h :��ZQ��^=5O�CV����6�f����a�mB�kc��w�C�y?���g��,���.��St�+�(�8���o�]jS0����������g�9����1���1��y^lm�� E��B�	QY�@B3� �~Y��;0C�.ٳ�H϶�yc����� !|�F5�;��9l��Q�c�)܏%���xT�*D��%x.�	��K���4n_�iL�*�7��g��z!6II�k����U���R ?���-�� ����?���"�8�r�%
:D����8/�.�b	`�w�$���$CK���S�'��<iXGs�W�y�/�`�d��.���7�P�s��ڂ�|پ[;����A��J�PQhn�B?=+�vFg�?#AϿѤȵ=�"L��?��g&XW@��}��B;�R����F]S����Ǥ�^�o1�]������5/�cI���?�������B�i>�/���]bN��/���^r�]�7��,�0�su��ǳ�{���K)FPbya"�s��al0`0/{�)�s>-�����c�K�8=�����1�/���0�\��X�7��-��X68W*��p���mf���'�9`+�ߢ��ĥG�-������H�F���/�+i����|��M�@��@�g���lٍ��W���%2����Z^dQ�qS��9�ub.[$Kx�f`���=�mS#��j�Ԣ�o,\��g�4�-�`Z���Ҵw�V4g��������^l?.�|�mhp�m|@����l�%�/���(�Q��؍cjK��J�%�P���TC%o׽�_�9�y��q��C�^K�Q:��<Җ��g��Ԇɍ�h@ύq�W�K�y�`��yǉNn��l�WL0m;#Iޔ�1�)����n=b�#�nx��K�ĥ9���a�ܯ<UA��C�[�^�,Ol5��n���|�u���5ic�D��v��ѡ+"\�m�_f&�d63�����0K�|�"w�9kԢ�aU���o(���d�ޥ����M�n{$f�9%��vj��)�p��۵O�T@ه8�vm��Y�Mg:;ܶ�Rt4&��!Wsx���bҖ4f��bG ��߅�<���B+��bNyI�S��AOm�˾��(���VD��e�]��saꮷn�ݓ���B�Z�K�72�n����z����CA#��b�&R=3/�.R�����M�	/�#8=���/N)���a��mLg�-b�J���E%�&��g~��Aw��p$q��~�L�\\@]˚�0���z�bhHyֻT��������ڒ_�v��v@��|/�$��v