��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C��Oҷ�$�S�u��B=R0R�E����X{W�yh�)Y���ȷ[��Y94Z�|�cLP��!��U��se��\���?��C���k �:5\�,��I��l��:H���C����#RH�t"�qͿ�ǆJ���F�J��↫���������_��g0��?�/w��Y�?'�R���ئ�m�T��jmdK7O�0���\?�m5&ě�	��];��v*m_�#Z�M�{��f��ٜ��ʬ �&�5(�^=�V����kf�|Y��H��Lz�w��kD�4����4P_����ΐ�l�cS���x�W�pl���[��n9�{�dUp�2�߭b���G�~���A��?c�i!T�4Zd�$��'���.�v��g�y��;�g�r��j09t� d��*���\+�u�]��:&R\�Ji�Ml5p��8cNR˕������5��]htП��jC�ӥ��?����.
`���� �k�Kr���=��{��5��H���a�>X1#*7^�\w��+�kN�WR�nwq�Ir����nW�9	f�.Ġ��.R��x��ڨ!bI�`���ZN��1%C���U�Yv;��^u���!�gȡE0�O�aҥ�)��w	슚I;̷��V�q�dnMN/�,��CwUșne��H�\�B(�O~������C��\Bsd��i��������GϤ^���oc����y!�z$}\7>UM�0�,����R�;Ό*$�V�fO5��L��a��S�������r�.���B������U�m=e1�er��ʣY+�8��z���Ϟ-����(LX"s�0�{,�`Kn�GX��D~�|4�l��
��Y*'��V6 q�����!l��7o�u�M�4�r:"V�Y��SCA`M[��S����5B�����4�ld@�?P��d�B��*�͕�[�]�Hv�ߢc�2A�]d[�����=��@S��D�^�����?�J�'A�9�н؎�뜝��]����D�hgM�2� z�~��c������̭(���4�d7̆5+�g�]���L8��gW��9R��%�k��s(5�I$~#z��7�Y/�L��w�X5n�^��Pm�Й̓ϙ]���da���3���J�����J�#=%��;$�7*7@��a�ؙk�ȸ�{.u�f(�A�ܢ�p���g���U�p���lH�	
�u��M6��4�0����7���|ע�ύ㕴4rt�zD��r]e�FOw��&T�z�S��Cɹp0��(\�3S�ﲜ�2�xN��F����s�89(�00�7Q����ri�l�Z���8�"�	�=���#��zh�T�7�+�]Q�=Cr�p�@�ޒ��-҉z�����ipR��I��"GI;�a�������`v�`� |�SK��a�/ѯ3��7�L+je���X'4��
���Y�j4j���y�}	?V�1� &E�/r����x&��[{��<�"�R1m���t�(*�Xo4Je�c�A�*of�J��b�3J
��uB;��)��4(\�;���"���xZS!o^���N�'@�D���쨇�	y�N|�}��X���va΃�2�t>�K��?HW$�B4�b�7���H�-�cb��ہ�Sr0;�{������ ��6(m�,{wy� ��H&�W����)�w)��Ez��Yӌ��*���P׆����ҳ۸d�䋘*�=ê��fɱ�ܙ���-��]X�Pq�*�CQ�t�P�b������P˞�Њ�*����܄â��.�h�_z=Ҕ�G4�0^�Ui�i�;ʀ����E�J�L3H�j�i���� '���Z�/�*o�����T�/:^ڤ:����]����;�_o*|W���7n���k�]\,R�ܼ�XK�=��|~M��B�ǰ��)i�QR��7N]�JW��6ى�7�J��;��7����rb��D��gLJSc2�o���om��+����Ę:� �.��1�s�RR�(��;�l�.\ks|�#�#Ỳ:\IΉ�5�й@��P�5���\6�t�r�Or3�J���m�-4�q�u�xO�qjDAͽ���\�y/BcpVCZgZ9�G����A���
���9zܒ|a@��R,w�,�VC���Ժ������{@?��V*�;x��9u�%ϵ��ńE�ߧ���4	t�����OPA�󨪣^ڤ&T���a(�����&X�����D��6�E���q�mx���������@N��{{-}�7~G��!q��|8�kpC���W���A�q��h�FbQV���d�Y��\��L�R�t�x��˷r>st[`�\!N���E7�N��	z*6�i6��W�e	
rf�m
����6�1�R�Q{F'���y��Գ%nz)s�(� w� ��OESp&�ս�<�ʳcE�aq$UX�B�o� ��ʷ��J�Cw�{arI��@���>�saq��b��q�l�;'�0	�i��f[���O�����3
f4���i�b���:3РBp���y����B���r
�V7qŅ��ʯ���gL0��F�b [�@��y��wg�bk
EN����t4��kXEطkM� 5��R���y�eؖ�MOW|�%g�Wy�ч4��3ΩWm%��*�D��)�1c��B��Sy�T9�Oe1���K����6��	��l��a����r��w�Hm�>�������R%�g�t\��ʊ�}���r"Xo�/�b)��\>�sGz�ۤ�������a�MV�2 ��7��4��%�?i�~'T�^����5�U=c�B�9M��Rb!���$�YCy�H�|��\ ��n�e6���/�0o����M�����͗������*_x��Y�ڗ�BA��l��um�vosş}�}_|!R�M��]|����dͦ������P�V��Nus�-5I�RU�_8���f!��)�e�m��u��]�ڨ}U��|�@I��xhǧ���� ���-��\x�<Wר~�ܱ{@�7�UA�L��9����e(g~�k�95�z�T~��e\�=EW�-{���+���5��yLP�ߟ㮝��<=��>���6" �֤�� ��:GxY+E�29��3��)d���N�+�`�M�{0S,2� �����
R*t���@�ٟ����B�P���~jT���-��j�0PΓ	�צK��sZh�A����_}���קu�����La��R�X��3�B`w�/�㒺02_�m?)Wt,�y�#T����� �q�.�Б�k/Q�C����R}�<YKh�B2|���y־w1'�1#{V|�ľ��j%K��Q6;�'�@e$G+��:D�9�~�nV�?M|��4$��l�3ҡ>+�H�_�P��Q�zGƏ�x�vO/�l�q��Q�m
�
ś�ʫk�0ۓX�X>dߨ�`2���X��t�E���H6�����Y�L/���5c���Z�ћ��ӠĖ����N�?nǶnI)�1�K$}E��^ѓ/��=QТ��0�Ǌ,�O(/<�h���ѽ;���N��v�&��z��EQ���X<^��nX�!N��������
$�y��]e���P鑨��[�	�宽��6����o�gI�>1��g\��I�Qp�.����Gˉ�,jYTE>S��@>��"���I�޸{��g�]E�L3YٜD��ʚ�#T�1��ǒT07γj��"K/�t:#ܲMY�Qz���^�X�(X������7%54�P��&�R�M�Onk��:]k�c�A]���o�]f����py~0��<��q�����O&6���P�n��E&_�=�>��S�~�}֪u�`#�u�NR��%�o�SVh%��*vh��㹈L7k�-��Xn�K.٫;�c���#��{��=��xF�4>Z�H.FY�dPD9�x��%�P�j��vpϹo�����(�<D��S�:�1�F�~уT��:Y#���p��ÿ{���z;#/,��K�td�'h��O�9�P����+���i�30��2}���]��]@��yݏӘ�[�u�+��ґ�5+�����`��BcUD����F���\v�8D,�a��u�~	�UM.Xo'>
��2�Z�	YR)g�4�T��-Ղ�X�2ˮč���KhE�;�+ �H��6�E�ױ�h��%�f!\�y����~�0V���T�a�Kf��_r)��>lv��x�`�3k�J3J�b�\�3 N���N\��O ��μD� Pvғ%�Jc�ˉ}*�&-T�J�(��r�x��HG�_�*�Kw�$�[E�q+�`�)�a���y+h&��g��a�h�t�*`1�(�MX3z�a�>~}����S��(��v�����q�Ä���AD�NjqD!QEL�	�W�i���*g�!l���UX#QbG�Г]"h�tj�x �WJ���|||�@%���=P���� ,[������?3J|s%�$O�]6���jœVB����6n.�H��*%`Ɣ��J���*$�hG]K��pޢ�s, �������]z�U7*�p�^���W���im��S�����aS�P�j�pr�Q	``���܆���}1)�8k�/����mTtQIa
�Z�=BQ8}��ojlv���OK�')�b�Mf�Ml>8��)2���V���C�%G%I:�p�rG��q	G}/4d�@{۠|X��J�-(�sy�W%�}MK�.���b���#�ږ���iUm~���Co3ߍս'S/�uI�hء�a����7.��5I{��\�	O9� `��M��uc�'݂�T$���MZ��U0���'[�z�0��ڦ��^�:IoQ��C�%�b� ,{��y*ơ�}05U�*;7� �>s�h|���;('[1���pS������۪D0| "��;�+R����e������z ��G��8l丨�y��s��{b�����Ƽ	_�Z���Y�2�����������h�꨼��E0V�7�Tփc�M���8��-��\�y�Y��@����Ǟ7�:E�	�g�թ��!T	;���e$h�VӖ7{�Ǯ�"�*�;�y&����&���X����{U��xT�[<d�׵w��s6�]���ӓ�~j��0�������v����	�#��d��Q��{|����e�N� WR���h�0'I�v��Q�X�k"�{<��r #�w%�v�� �`�R�L�WM
�}�%�_�m�^���Rj��5��B�u�P���|�/��h$�0}���C�0���4�>��:(�f*4���5,��
���ǂNGѢo�)��l&��T��� px�6:F��T���a��¼�ٖ��V�b#_����}B�+���"R[�ixK���/�$�D$u�� ?|���#b}���0�?"�����bz�}������a�PĖ�~u%�����@E���J��'��w�U�);��p���l�\�T�l�)�R޶�8{�b�ҵ4Q9C�F�Tko����e���|�����0Č��8)?iJGp�.��ZJ<�#V)�O�a�i��)P6j�K�$��4)�=ҿx�d�]��;գ��p�.�t/�~$.�R澪�j~�C�,	n����b�]���V�t�S���,�7wP/�7սyB�O.=S)"T\�J�_vd��]��,(�����up�dcxo�4siް�Um��x��Go2���/Y�D�>h��,�������QK������m�ن��6:;U$B�!!�Ekw�/-�(��Y_0�i� �h9�2�QP�'T܉Rc�'/{�"�BBҼ�J�މ���n2=pi1�����/�9�7у�+��m���y���6���E�uRj�$������w���-�/���|*��Qu��d=��h<���9�f�g����6�@'��?���d>�ۃOh(3��¨�+A���OW��Nhߔ�~� ��PC2m�tU�9�I�#��C���>$��6P�0��a�a��Fc��-M�y��m�6/������a�b���e.ZZ�Y�����'�x����.RKK���d֏��Iu�yW�/:>�G�Uq4�@K�� @fP���o����;w����<���b���Cy��:N����p ��fR��`'��rvc��W�G̭jDT�3���X�O�Վ�\�el��#��K��&y寖���!�4��2��
����Q�x ñ�D�mZ�p�C0���ۋ#V�[Ǔ&A�s��P�1�� ��A�0��D��i�S(�t�e�^��@�Z�MN�XSea}6���\{2��nm�&>�O;�s~�*1�J��g�{���#�'mf1ͱ%�
�����+����̓N�zi�/��T	щ:��p�`�/�����@���Q_M��Μ����`�siJf �\w.5z���C�6Рy�=�>MV����1��~��3�W3MTH }��Sz�O.�v4�*�|p�-�:���d�F���3��M�=kj\��c��ysk�2�t�k;�O�r
5��ΌM�9��F
)xu�L�NE��)6�/��ku<*i
�P�Y@�qq��y� ���2�F��ʲ�sxv���|-�]��ob�Y���ߓ���0�zf����2����1.����(/�X��Hh!<�󴪊xl_�.�g��v��Ee��U�Ls��=sg��@�%��j�h��R(ބ��h5J�����C��%�_��΍4^����-8�KF��z_*��b�6$��k����t���E�hD,RC��HI�y�;������4E��?�O-#�AR�(r|u�.`�"����Q�#U�����J��
��%�f�}��t��|#gO��]{Ex���v��W �=�;��h����b�c��.[��v��>Ej8{i#v:Q�d#e�u"r����3�ۻ���
��zN�������9�7��d��3эqB�P��Q8���Ĥ��]oR�C0��G�o�l��z$Yo���ہn��)�
����h�J� �~< d�[1јEP�P��\���3�����jד�����D��,8�!4�|�|v��H�sY�2b[�N���V"p][w[?�����{��-s�G� ��+�RR��="�8G[USj�`;�xgBR_�����6�j�K���7��~0�k�/ViT��i"Z򼋮I�؆n��S��#[����,o��Nd`�&�~�e���������2��b�To�e]U���ZS�5I*%��� �T(k�<g���\K}u�4��a�ԉy������X7Ȭ���Y����K�=��`ej9h��R���,�O��<�5
J� �{����5`���T�1�������vJ�w�����Z����%����i�
��.6f���+���i�c
ݘ��Odp�����F}rjd�*/�&���h� x��]Ku��}�#6B�Fxi��j3��NWw����@���ss��L�n��c�����w]	67�Fozth��,x�-y����M�z�M�B���=n�kM�w�.��ӷ�%�I��8B�~{~gC���E�2@�'�_���Q�M^�ѡ��lJ��b�&���p.R?B�y��`�㏢A�9ծ�e�e�-[��	�XqEI�!��.Б ¡�Ҷg �e�2����78�8��4y��s�̤���J��86V �2�^��1_��5 $+6��1| 1�1��d �F[�g���zqφ�FX��[����H��p���]�l���ȏ�zb�~ZQ^uA(`���fl�op�.�2�����G-S��2K��C�8��;[��M`��B�6z���0���/%$S,��a�n=@�*4p$x��<�A�E�nV�.�%�K �-�2D:Z��p	�O8�M�dP��],�cu�1��(U΃}�]D���W��	Vq�/B��l�[���C�O$��>@����I������R<cU�j.4��GS?�.���ދ�?���a�q᫁⩮O���fv��!Rc��:��\�K���ߟ���y����jF���0%��~�/@ꫤ�tNp N|�	IT.�21ǒx��;x;w m'p����^�CG�+��3F/C��Z�n���,S����W��Ǖ#}X�'J=�G���C��E���_	��/��I�����Ai�%�.���)�L���g���;��he9��!�uӤ�^���F_���ɏ�D�H} �Њ�ݒ��4pf0E�D%��~�l����������r:�L��4��|��Z�K�P��d4�m!���vn�����H��~*VF��f?��뽖�����J�6���pS/�����O�������|�&n��L�WΣ���d_\�Դ<.X��6�h/�fK��9Ӷ�Ǹ�]���x�G�?db��⹳�f'�)��d�ߢy���=�3�����5S<�)��&�]��*��U��c�+��dl��_<}j�f�L�O3����+��Z���0J.q2U�����H�}a�@����O�eVg��`G*�-2�kK�e��!��̮9��i�&��Q?g��;�\!���G,���^�[/7�d�󤹤إ���U
���d�#�  \C��09�g�($\�<�S�%�7���]���4���	R�UI�/s�8Ɗ��_Q]^hq�2E��Ɏ}=���
Q�b�#C^?jJPyemá�q������t��؉�P�|��R�����+V�`��v��E��p�UK���TC�X&j�F`smk^ϊ�����*�g*G��S��.߽쥦��x��0�Y��t�#/ByBS�+J�Z���Z��X�S�o�K�� )��@.?�2�W���4�����������r�P�~h�S�7)*PS]�!�
k.��!gf �|�k:*�=J�M��|02C'�.��eZ^`������qل$|8�]�!�#��kS	X��u��W��>+P^&W���JӜ��yB"�(a�*.�]$U;y�+p�����`�{��x+{2�:9g*x?C7d4^���c���R4���w�I�C���q;�^��yԩ�g����y.�k�E��X":�������-2�M�}y���cjg�z���N�|[ q���j��z�n���!�P�KR@����:��3%J�'�t�z���Z�K���خ��b��@�n����;e���q�"o����_���O�	�U�񼇚��Jh0���xYQs�+���k��}0���Bm] 9(ޖ�7
u��~.AN�_H��<�Y.��u�N�~��(T�x�ΣܸN�w�T[}��u�FPR���`���𚵌�q` ��1�����)?
�J���{;���t���p����E<� � )Ef�;=�W���p�М��;�,�r�CZU#�g],��w�)N�c7�qIpӑZ~s ���8�+/7!p7,yR��7 ��چ�������G�Sb}݁�o�ْ��W4]{<�2d�J��E.S�."V�+Xl�&CyLG��)=��b��P_�� �4�{}R�5�ϡ�bA�?J��wLֻ������)��[�S	�ER��ò�`� FcCG�C�����V%\��&g�;��z%��Avx=E#���j&��FG�OO!$F�]�w��2�]��g�?x���$��Nv��i%�?����h'�n��`�2���F��,����˩������=�����[�1fc�+U�)G.�h��R6��!��cp�v��|��e<���{���&vtt��颚\d�/�0�{^Q���"p�� ������+XBHQ��2�]������f���̝��|�G��8�!*�o=r#����K;4�qw��y�\~o�J+��P��z���b0��+ �Y�\g�le��1+�Al�75t�V�#1 �9��Y��'n�l�Qfߴ?�Վ�����(�vKe���3q�n�3 f/�f5&)[:�4ɠ���,�p5�m7�J�U4�z���/K���.w�4c����לa�����|�{��D��3�9.�4��C����,y{wj�s���(-%�r�h]9�֍���4�@�9���L�_�&id@\T@�N �ў�))#��k�f)-���#�P�F�
�46!x��r���}m$�����"YH��-���%�楓v4���t֘Ӂ���ޣ\�X�d���;Wx�h窄�Xĩ��nF���cJ����r���7�D6�c��|�M��!�i����$�\��v��5��qC�w<6*���@���� 7y��S"�/Y6��c:X<.���6{LH(��d��v��>��`s����Ӗ�?�#����]�ƽ7@	�4��]:BL���ƀP=LT�@�ݗ,*�Ap`��[�VF�S� !+#�:,��N�*��8&T�,Ty�E��	�t��r�3@qlLeׅ�9��U�-�b���I�5�@�3=t�մl�y�����L���/��+�M�L��pI!�[_6�R�gmJ�����X�^c?���B�.�x�IDn�Υp����꒰��]mk�}qi}1�'_���8yo3�bܓ1���B�����P̎j�SƼ�ny_h�lq����(w��A�r�����;��Q��R4겝��vE�`�ft<���������A9����R�	�\���U�O���&�~-�����0�5',8!#f�Z.���Ev�qY"���u��D���|j.ĝ��f�A\�Z��>7"9�uz$�!+rx�z���r��O��<�$�rq�^��_��!vF.G�ޙ��s�l���=���I'dс1�H���H���7��=s��l�{�ߺ�.�rQ�p�q�hX7��� KdE{��A8�6"5�r�ô@	2���~�o�q��r��WK��c� �Z�`twR�(2M
]�S��X)�h1����r]��*�Slǆ��:rqj#wd�$W��)�I�{��«i,��Έ3T�ak�#L�d�&+����{�uVT���ҳ���MV��p ��m ���B�٥�
�iV���A��/��������%�v&Q1�v��s����B=��t�!ɯ�fԪ6jSR�o^;�Q�+��69�ֶl�������7m��x2P�**u��U�QE�ǲce=E�0>�/[�8���t�_t�uQ�g��1��F��Y{g���*9.�|9��N�da{��� ����Cp �|���:�y�ccV�����3B�d쏼��ۜH����6�����R�r�/���Ѽ��2qw�Is����%>���h�������-�����$�j�6��(08���Z����4�J#z��>T�G�Mr�����Tz @�W��*��5���������B�WT��z�-�P�j>��GΓ�OLkg֝w�%�3Q�~��ϫ�o�T�xk����ݻ#ɸ���&��iH���/d܄�w����{/��sC����͗��A ,�r��Zx�,Ɓ�jݩ��n7�L2�O�nd�-��%��ը�� �fl�bB��(��P��J���<{`�R�{m����h}դ�y����W<��%.�A^듵�"c`�ܽ����y���ݏ�h��� ���ZP�'��a�f��"X��bd?�ׁ2�]�h�da��J���d���^����T���h �]����t�8�d-f�S}>�?'�v*Ӊ��`�r%�;��H4�6ɼ�m��TZ�3�5��#>��-<���b�?���xTUHJ'qW!T{����?q��@�3xP���)�
����{z� 4�j���'ڿ	h�T/�1 �~p	���k�$oΈ�]���
���Z�R�n�hcZ�m
�Wd>~�(e۝#��XX�-�u��'L��J�q#��
�޹�k?#�ZK*琱z�M��`������Vڪ(fr�1X�P���������@C��"&����^�F��̵#F��.�4x��5�>��5���0]{>+�������F({�i�>�2.!ByX�&�2>S��s��V�d�ƨ�ݲ�N�GղSd�瓹��g��g���V	��?E����'��L�
~��,�ۙ^�$�L��qҍ���Ki��E 2�Q�=G�KI����u�\��K�v�f���-��31%�a�Q�,��4>\��_��	��*ܢ�ݪ��� ��ò��^H>�U�8��km�Q?�ћ���lx�:,9���xl�}R=S���2�޼�Hê�H9�KЅ���B �cF_Z���څJ�}���k1r���Y������*e���Y���XY�S�Ƕ����}��^�!��c�!��ϴ.� 4�R� Qg``�q�����nYr!�y��[g�OŔ��㢥�Cי����\���\pt���p3�\5A$prU�����$P��R� ��l(���wڬ�(`���̚E�p}!ѤsP�h#=H����X��b@���6�8�U뿘[D$u��mR�*��O�3�~����ǒS�j�i�������~���@��{~}#9�*0�'��
��-�r�:<Ye�P_]��-y_����Y}w���|�6x�?K��cM �=��u�i9�<���[g҅�q���`�5k�'���C"���\�l�]`�p���hk.��|�"��o����>)mkO��bL�_��4�V�g�ԋY���ޛ�u�bލ���^����M���;�HlR��<;����d-6����. ��}��Õ�fݰ�����{�zy�Fky�x��
_}�Y2�΃
\��v�U*����~|�P&f�,ˁ��.�em��y���RO=~롮���}� �1���� U��V_r�����A���.���!���s�&���Y!�hy4��<���X�y���ݵD8ǚ�?%Zn��faf��L��!�>5_N������!-(^f.4�)�-��~��H��ꄽYnX�#y'"����[��ٗK0�Hy��4��2�)��$�ė�ڱV�w�^/'�i�"�kE�\�~(£��n"���wV�������m����TP;ɓ�u��x�m�ޓ�y����R��dp.C`L�hL���=�j4�r ec�R{��꾨�'͟ߧcSj����Hdr0���
��BZ\V�b�$�����������&��)jx',�@K&L�[�������G�z��Ӫoa�NIכ^J^7v�/�d�����	������bC:��gϐ]�;�I\jܹp���J^����4�@l,� �F9t��Á?����������H6J<cI�0H}=,��u������~��&�����_R��ހ��E�����qqQޅt�����Z`H� �b$���ݛ�棱/�w��Kys�G\yr
f���f� �j+yT���RF'��(�C�x6��Km�ՒՌ��aa���Jpb�;�=��X�+%)Yũ�rCh��H.Hm���AJ��s�=Tx4�pHLU��P4�D����(&�b�L����ſrI��\S�u}8� ��ں�As߲�T�$]_�J�kum$.�Ҁ���U<Uw�W�x�H�˦�8�h�7�=A6}@��\Z���.h*���ʜCgn[�JƇX,!�X#��O���[�U�j������_�6��gt<� �9��ũ�b�䪬bZ�$/ؐN\�=�F#e�p����ɻ�d����}o���:aM3�������K���"}eN�
i�-�6!રi��&����#Ƹ���L?�ٗGK%��\��Vf~���pZY8�_����sj�*p�(2?�lh{ v�.�s;��ET ݏ�xko���.Kk�sӤ�觾(�y��K���B�'q<I#H֣�c���8;���@�r�P<�9�X��J�ʖ�4D�*��ԥ{��q��������ZOh"�?=�n��ٓ������ha�8S�Yx������� c��UY��V�Y��S��V7V���m
��į��υ%;K$:�2y��"�H6yx��Z;���G)z4!�Ƹ�;�v�jF�wЂ��ᤙŵ�Q2 �$Jբ����j��&���F4�<(���Tq���~w�Κ7�#�c��Y@j����娸W����ӽx]�F��<�@g��9��-z;b�;�aˋ'�1#Q�;�z�l��Z���Tԑ\ji��OP��<@� �Ŕ���
cR�z�[���Ω^A�W$,�fΛK�X׷�n���^!�~��Jgf�]Q�Ĭ'f_���NW;#�I��V�w���MQy�r�������Σ6�m�=@��s�H"�ô�g�;V�?�����+3?�-ѪRJ��.�>M��=B=�h�H��וg
KPqu��{�L�Y7kδ�^8sS�N���;�U"���1u����`��C��O��ۧ��&��`{�jh�(g�u|d��b�_�r�E�_q{�?q�l@�~7}�M!�g>!��Hʕ�]�1��:t/�f�D�3mpod�˔�!Kp���Ӏ|n��2s�ZA`6Z+��omoů�tb'¹=j�SIV<`�Ě�
�F��[�A?ۿo�)mI�.���y��&o�b�J��] b^ӿ��t�0'{�'m�4oߩ�NɰPN���GC�a<��:��$Xh�0G)��4Pa�wS�BD1��KeҜ.)����AI�\��"�m�`�,�Yf�Ajh8�I�iVڛ� �_�WЎ�����	����QD!��q�MP�/��4r�s�v����_̔���wwn�::(p'*eKN�֥�:T���tF��t�<⌮5�����X�����e����x��Ai�,,��w����xY}� �	� BYY�}J|�Q- є۝��'-�t5��d�O���a�h\ؔf7�nd/��у@�{�/�É��r��:"3z#�K��j�^��7!?mYy1
|7՜�=�7�hj���Nƛa�o�sb\�~���צs�b�K���i_�������ϖ;3I��.���iz	��C��Lg���b��n��w ��D��{{�<J�X�f�G��ۛ��x	��*Ң�:yu0m�_>�Ѽ��˚c��6zʙ��$�M� ^��;��$�G���7Z����o���Ɔ݈��X����yTn���ъ��#�ա����`���cѻ�D(��Ŵ�:!"c�r?F�Yt�^j��n�ɤ���K���yBe�EX�,?geÃ"��֦f0+�0j��F�}�&Q��!F�I����N^  5�
��:��8'6WWv4�t�O4F���WjP�G'��;(�Ҧ�+�1�/�rr�N,;k�5ܵ�c����䙽*����}�.2k�g�i�,�Aф�愲{Ecb���kGHT\���_��uHK���9�$لh������s�?��
F��P6?��v�9�k;�&�8�S�����rf�hd@�,!��)�y�@�m�a#T�V,���Eb^�S��,`�%�䧈s�r&;��ʮ�q�����zib�� C92�-Es��$��{gK?K����î���WL��;I�z��h\r����_�|)�ظ?b4:���ǳ��G镌� ��Jv��wm�8� �!�����nF��Ϙtx,�$0�z��WQ�s�)�Z�Dl�Dڃ�� eK�Ac�D5uV�޽Q_�X�)ӣ��5x�O�7��!{֕0�f��m��[�}��Ŏ�wneJF� K!�1�Nٯ��a���W���$ߊ'�ґ�2��T�B<X��?��;Ju�}vӍ#q�	T���ͳ�T�$!R��w*wi���X�ɮ�>���-�%=C�b�zo� 0=
�]��C��4�e��E���w8ᐎ��	~@������O�0���,Z��9�y��W^0��0���Q2�fc�Q��^��ۻ� �z|�7V�k���MHhV�QrWz�Tfً7Uz�/�;�|��
�2���B���B8��q>�]e��Ww����
��\6�v6����"�p�¦aP�N�St%{�x8Fb�r��咿Is{�op�A��Q<?P�7��ސO� ^�>D&M�dUm0���Z^�� �� �+p٩�؝�)�=J���z�t��z9ί��<ģ�EP�?�"�
��>� ��c(� |�"�*aPEk�*Ưke����JF�Z��&KCd�������.`���`~�-�c��`@��5��g�A�zծ��2s�t͂|�)��ײO=ub@Fw�^
6h��Ώ%�j�
��`�U�u��\��sjz+�����\�ޗq�S�Fp�+5����H?��ƙ��iI-��l/��Ċ9In~ai�k(=���^��һ���9��v��E���T����h�!]ӻ?�wL��MQ��< ��K-ifɏ!TjK��}	PB�����vVo�`T���:o��7�k�a������>���)��A8�,�j���c=Jc�\�_+X��E[��U��>�-z\a�/���:0��[0����C-�]�`�q8	(��&���>U����hwQK��k�9V�d��ƫ
���dj�`ub��^�qPQ��xy���r[���4!9�l��4�ʉ�����
K���ɇ�����y�nAc�}-_2)�%w�����9rzv�a͌Z�D����F�_<H�p��C�6��{&ME�mr3��f��8�HS!d$�������䬬\x�84�f�Z��K��Ʋ��b�3*���rlu��L�c���3�%d�Xg��������5��-��i!iؼ9�0)�,VW�A�<��Hf���Er)~����2�*�͞�
�=Z��Z��x��S���d�E�	�_1�
0ʠ�=GTMOǻn 0~l	�Ҝ���3�r���M��n=J��"9�[D�yV*���ѹy߷���Ա'�TFE��]�Pw�|�=�#ȁn�nV�_�}��n����uG���K����aT�}2�.��/KK�ͫ��S��|[	����op���\��[A*�p����p�l!�$tt���j]lm~rsl^�1j4�o��K��#�q��:z[��mvՓ��pQ��]H���ն�5�w�ȑ��Q�t��r;�)���_R������$� !&�<�\w�����c����l�x L��b�i������y��k�E�P���@����ה�3��M�}�)��
���u�F�i&T�r�jV�O]�3i)�#�,ڇ�����ܨyU2Ns�ˉ��Ɉ��h�CM��\O��~~'�5���(ݕ���?�^-ҕ���-���[	]�V ���o)6b,�F�<!�T�\>�Ƽ'�R�YD��e�K������t�R����7%��j�X�O$@�r�u�Ո��������$ 0��lԢ�-��\�@O�V��~O�b�2�=����u͒kk�Q����(ю���AuO:/����vl��T��!�������[��	+�\�}9��J[�4̍�i
!d�,1C��ē�_�Yx�Z�Ï��<�K�`>4كK�|[�-�K�y+b:J������Q�}$l�>@L-���p�H���Ȥ$E��k3�xR6�P5�wi����p�J{'��k{yCHn�6���?D�&h�ƕzZ8N�BS�d�J���M���tP�T�����P2��g�9���e��E	Y@:�O	�
���p�d�EQ�6��b��qE�<1�a"$����ٔ1��cS%C#8L��U��q�X<��� �ts����Ԏݽ߳~��a�0�]8O��J����+�%�nCG.�$�����?TJg��&ptQ���<>����������|"y�[2B
u��x��}{O�D�&�>f�W>�{I��P��C�p�%J�u!�m�o;�pYO�ڒ�	�_Z%f��q��?����S��P�{��i�(p�/V�҉��T��[0շ� w������[��¹�T߯�J�Ba0NuƁ��йl���|��%���)è�|3,�l�S�~]�񎊼Jx�Ai�����#��D��L[ޥ*�*e�Y�G(�:�\�d�]�C?:�b9�+�Zp�/���U���ߔ��cR5�G����w�َ�=)`u�~���)�w��,���'�E��ͥ�Q�Umఀ����s����}a�l�����P�*s���p���OS�@����s�!��G��.f�]��G��ț����.��i�Z���t����oW���s:6z@��?�0��,]��)4��k`.���&5��ZszÄ@���b�
>}p�\w�|%��!O�uu/<D�H�����{�������zH�&G�E�>�ӡ��yn҅�9�$�>��n�F��i߾a���0��}�����RG�-,��9AX-t&G�% �x��}H��Z�E� ��\�U��@F����M��'2�w7���Q�!��3-u���������b���h�"䘔ey*LΘE���Ը�YM�^�޵���|�B<[�qӦ���e�Ö��ě�qg=s<��A����%-y=�-"��e�e[��-A>�@w,��kA4�fVGD�@�q���?-H���jT�o��a$�3�Z~�1@��N�d�e8�A����-;�-pG���w)�,GC���!1�̷��h�MK66ؑ����EX;�i�ڮ����O8IM��5/���ZB�d�x2��Z�XXG�)U�$��n6���+�ދ���>��� ɪՖ	�	4��A�uJ�4W Z�����c���j��g(��{`�5=Gs ��r|%h��zȠj�y���5$��`F���/���^��*9ȧc��bD��'G$��+���KtwŠ��Whk:A�2�f�`F� �ê���^�]�\yN+��0pN��ڭ�2��z��&�%�~��|�^w�t8�L��,�F��
�9߈vt���N$4qH�רΏ�څ��z���o�}���E����iբ|�a�ң�$��c��q�<���RO�`�OMZ!�����p�Ǐ�[�B�\�	�	o�2D���B\JK�� ך�i�3t�����3���T����\ûU�:�� j�e��w�p�Ί:�v�������JJ-�o�L����l�� �@��6�q�(��F��V��8d�k��������sym��\�'7��tP$��u�!s|/�[ۚ:S�b�&�ך���j�G�T���!頽��g�{	fP?��^ӆ˪�S�A|�t{���8b����1��39�t���aFuM�iX.45�^�ը����� "u<!��2}���-��r��zV(��,Gyᷚ�h��`;{��P����s+�xÿp������
�Y��F�D�!��Af=���#��C&q�����l�H��
^ ��X�=Vv3�epE�?�G�P�F��O�8��b�u�)LU*A��QNƈ�����֯L��o@�as��3��)�	gvO�Qɩ�}�z�˟A?�L�e�z��a}�S��5��}z�f<�u�`_}�{П]&9)o <e�b�P�@߅��;����w@<�)y����~[��<pl��?d�U������Oi�W�V���4�73�i��=�a����%k�-�!��i�g��>�'�?TZ	�]m���c��WͰ�2j��W%�p���U���"����N3�dZ[��r�)+�y/g�J��2���'d����~J���*��ܟ�l;���FXa�<�$j0�Ń�.�˽í�O~�|����V ��p��f�o]�Ia�+��d#�,ʴ�X��ݜ6�*U�5��6�ePD_��(������ѕ���KH��>��e~:�.'#OǊ�e�*ǆ)Nzh�U����݄�(oϟ��%c�5�-�S�=��c�7�v�q|1/M���џo%�����ƌ���o�<��˞�U+����_FiH_���&�7w�O�L"��v90����󵕁�{r�j��:�������#����+�}��CA�)<^�d��O.1�M�Q���G3��O�����Q��ե�I;^�G-/�|��x�Q `���\w�(��ѓ0h�7:PJ6Hv��^W$��/�啟U��y7XB䥨�K� <��9GF��k5KwL1Fv���&�{�/ɷ�I��U��+�U[��N=�5P�z��
t4�ٟt��
Ld���%��OP��S����S��*1��vH��#��iKN?C�H~,m�:�I�O��N2
84�6T&+�VKV@�&؇�%&m�:����~������u��F�wb�s�_���Yn-��5D`�����;���N���L���iJ	"a�Q8����"ty)��e�&U���&��&��vB���6�n�&�$,�5���񑮼<����'p[��6��({�((���kQ���p@��6��#���y)��tu�u��P�~C���G��aF�c���} )����|�e�ܮ@���1:3t���'G1	-6̲=�b�"o"�e$�?16(���.�q:#~�D9�~f�\�c�T�ʚ T40���|R5rRc����n����g0��1	��d���w˹W�iLW�j�ٙ!��3*O�EmJ�E`C���^����������Z�/�1��8��=�҆A��)!�@��-��߳���O�ϧ<��U'�q
�<��O,}F�캨^�G@R�Q��~��xw��/BJ��D�&��:��u �:��V,u[3��y&��@�U�{�U8'�7��]��	xk�Xgt<gM~qϞ����׹+e��;7�8��Y�=�����5��%eհ'x�/��x���ڪ���2�~0���1��'O�l�!���o�W�c9M�7���,~�|uF��H:��h�����S��l�).��Qe ��a\yz�jI��
��(h�_f���H��N�^l�c��R�o�sE�?2�e��t:�l��g��3��b�&�v�A��r}Nx����>k���2���hs�Wf���3s�	�nn�˺M�,�5L�R`����X�Τ�=�g���c�Ҳ��(�o�jU���^��<����D��7-���<���&ԩMQ�_�|��c���>�㒹�G�.ߜ{���I�����g��7O���7��J;�3�E�
��B�u�K\�ᔜ'TݸD���kvOν���!  �(!D?��0���|J�卐��� �k-�؁h�v�|ưe&�?>�8������&+��y�.�V�\q�σ$Q�
��D�rC\�{�$�+���}��k�}���n��:�u���hME��T���I�@��73��\U����ȏd<$nq�e0-Y�+e3Z	���o��<O.��;V�I%q\��6v���l�#E�7�1�0�I��օ�}ι�ՙ���ErV���/�ihf�؍�9��(�*�#=��"���ڮT{�m�Ň��JM��D#�,]a%B�35����"�������{|��ח�:1�k��x�q�t�4%�	��O��\���z2I�xv����dY��X%]�~|��Ȕ��Zʁ�L�RQ��v��D���V��d5=��H�Po*�3�;�t��1��lb��L�\�Y�G���E��� $�`2�/��̃0���k;�C�XI�?�Рg��#=�?��ͩ:�����ʽ(��;�ȧϧ������_�J�๿Y*�Ы�%���N��1/%�o���������_Z��}���e(v�@�Sq0er����������!"R������^;�c���.��eG���͸�������(C���FP����w����F6SS8�4>�]�h��Sx�"'")I���"de�Md�,����D	���PG�8ic
P��Ҕp��q�LY2M�`��!��Ulw��D&][6
i��LM%=�s0t���ڝu��Ƌ�� �5���;�y?��8B�a��`��j��we����];؜B���10Ѹ1��b`�uLQ
'wj{�^74�{_>��c�OO���ݐ����|��E��'4��BX�Jz���,_N�Q;Gl������􌪲�a��AUTГ��8�����@�5�k�R�=�.;י����D�[?�Q&/��3]5���kn��d���9���-������0��힎�J��3���qc�۠�0��n�����#5O���3�E��p�O��6z5�'K�r�g����
���ޔu���&�|�r|#\���{<�� o��B�5�U$ooj2:d���_z������q���a�x{%i�dhx��X�o�3vFZ��[?� �JJ0�]Q֊},�9���<����<p����J�����5fd��	(=�y��k��n����x�J�LifXA��&&0(�S���vj�\]���ǌ�I$^���qG�O�������E��Ltn�#��<+�5cآ��~�T�0�)����gQ�ڃ�����R�R.箨��s��O��4�֧����N��u���	�ҙI[��a���%P(B�`~:x:$$��y�pp�h����f��4����`q\��zp���ьOAF��BN�?���u�i_�lfq���a��"⻢��>���ql+��"?	 ��3zK�kK�D@�^`�6B�:`�	u}���e��:r7�-���Y���Ȋo��(aeZ�Q����~QI�`:{=&��bA�*-^o��4�i����f�
� ��5����a2_��T�d�L3�I�K3���f4�S�����r<q"��;[�=��K�" ���U����)Q�5&G����clL�bʀo�0��
�~�C4����Ha�8���ӑ��^�U¤Տ���|�����U��ƕ^��D�����Q�#}�° Y��,��;AѮ)���;�ӛ�~�q`���zX�f~ _v ,m��bUx�7��:��F>�H��z�S�&aw������T���2]��Ɗ��VǸR��T��\�D�)▔����z|-3� �0+�)�g'�� =|_J`���V��rѡK�7����r&���<'bK���uX�3�|Kp_P�F�����g%-��~�6��ڲh{���g�x ]�=���-��~�}|.�@�8�ȡ�m�N;��4�ҍy��f����N�2�9��8��6dM��q���N◘\����˩8�1�=E�b}�W"]`F�.���oyȐN���/-��5x�n�V�eſP��Ǹq��w.���GY��L�YJ��NJ��I��i�<�᛹�D�p�G��CW����� U|�u&�����z�ǀKp<�9C�-��<���v5F<#�*��%6cE�w�*��uo�@��|�q3	��)��rN�4Qq�Rg0ǸX.��;y�[�,��凌ah
���=HXdBB�$2�!������d �ڌF&�`}Ef#�[��N��X�L0N�,��:�[�`����6���
z�%����ɂ,1m`*�5ÈJK��e��' ��H�4�g�0���h�������J�%R��d��)x?�S�·)���ͥ�����/4�W���Q)!��쒍�wf
[�?;h�#��ٱ~�1&J��l�-�$���2)")W�v�|./l����:f0��Z^5�eɸ�5�Rz�r�^�e=�xǱZ���aH{�0gRϴf%�n��8:�\�Eja�&6�+�m��@��.��ｲ�����������tߢBLx=��+���n�j7v�U�#;��d��%|p����6[
�π�o��cj��.���u�.��t�+��b@��-���K�"m��w�
˅�z:��g�4����!=�����u-�h������f[D��(�x�#��J^�.���-q���ҏ�da�lo��=�7��|�n�H�����U�M*8�B � ��L��.FqKrp�h*�;ތ� �ry�#z s�>�igQ,��*Q�)B�Ę��Y���gԳ'�&{�>|���t���<��CF��e3�*/�"�����;
]����`��nm�����y��
>șdi�b��4�R�O��$,���Q{V?��9�wg�D�ZMȋj��1�tf�\8S���,��湚��8���}�0�NQE漒�Q��1����c=kŬ,�d(�=���C�`�����|Lb��~��K׫�$�c�ߦ0:.HW�W)���
e@�n���Z����='(�O
�*�Vp�ٙ��;���P\ ��F�
Xc�z���D���� b"-��F�"|�Rb4�i��o����?!�ٞ\X�.�c�)��E:��]�l�p-�����7 ���//���X)y���\$���ob.�1CD�YN�&b�l��S�V�{g̕����i-����5���@�=����ʴs:*O�%��)�v��	�����X|kb���PO�bX����vU�s}����rN�fk�L$���޵S
�l�zç(�M������(�s+J�tҘd��k����/� �E���=�n�K)*\غf|>
�p�R|�������.�+!��fm��1h[)F]z����5�{$��}>]K�Ʀ�4��5]e�[�봘���9%j�gF�}�m���۟+��y��Q�W�x�$(��,l"ԑ/w�� \wy�l�׹!����I{>ӾN�fo��^zCj㉵i"W-��:HJ��>U�L~`��ި�fT�����z���=�5Cb;��ֱZ1�, ��Ji��fƺ�;/���l�����Yte���Ɠh�z�L��&Xr�iv7֝�<{�qZo\:��Cؼ֚j'fy� wB���p,I;�V��"qj�Ý���!D6driۇ�P�L�2�]6֟���L������_�~�����^�2Ok�N_���(��Y�VKe�"w��% ��F��F�V��=nՇ�8�}M���,V��9nP���r5?���Ė��g{��/I��do�]�B��"�ߪ��w���a����I7��:%3���D$t��B�Y#�\�������u�c:�v�P��~&����R���2ף�l�;PY�h�����1��b����v�RHF���57��*�j�pu��A*�s�!	��N���P���	����Lf�~��z��'��|�e'�N�>-���l�0I��k%���Ƀ�8{��Y炳���|O��N�4EZ�Q�\�{�At�E��z+0�q^�i#�O���:��G�@��ӬT[�	��3%~�,8}�:-�-f�V;%l�C;B޷Q�ט�S�y�0�m>3����bx�6��i��	Aªܟ.u57~m����&�:��1�Z �� �p��-�`&E	#��.�֧�����&"Y�g���������7ֵ;�QW��I��p�g�{�2Z���(BBJ�j��	7~c	�"�����C����b
����֍��撑Ց���=7�����Xa��B��l
��SnfE5��w�DQ�`����#հcNIg����^ۆܾ��1���:kL�&�n@)?D���]�B�T���v����䥬���U����`�OdF�0�?rg)�U�ҹ�&�L�9s�Flz�D����QtQ{ .�[E��k�Us����'2B�{7�J�n�l��Yd�����Q�k|{�$`�Fu�(LR�ijtDʎT����%��Љ���5~��V��23�^�^����ɘ��
B������ES˦e�[kW>�F��t�(	Q81���m��\��U���x�N����{@>"9C�`q�ޢ�:x����Ei�w���E��3�Bw���Bc�8���X)��Q\�K�\��35#k�%=�z�e���b'p��K��w7����5��,	�S��(�B��b�#���#������$�DZ�ꍞ�v5��G|jklO,���IA;�q�@sT��^tLO^�LO�Q��әIƳ�>}�KQ�ƍ�*\��H7�2�&M�Ϝ�z�n��Z<��k�j߯AW�7D__���%/�p�:�\�����g�L���N*/�,zl�?�5?�J���b����Y�߸�*T�3^>Q�7�* G�wIr�H{�u�M��<y�
MګL��H�)2s�5s�����M��-bUB,��mn��G�M%�vP�cY;�E���$C��S{���%��cg)h��E?��,f���OT�}�$�2jf"ߑ������}<�Z����5#%"D�Z78����qaA���U���O��3aBr��q%�A���0S�qQ8�ssВ�o�(a�,}��*ӢQ�sV�5��YX��t���H�������N����F��EK�s��U�+��ϴ��!ܫ~�b-�1\�������_����׼VyUT~n�S s&����sT�q��¯�.pZr���c��x���rץ�:���֠X��� ���M�Ԏ�����F`u�Ä�R�"?	� �z�^�:�d��*��N ���U>�����\�SK�C8��R:�R�L��^��"���55E�^�c��!���;	��W�<�.י��x.�r]"�64~��ߦ�\�+����m��^G�n���T̢��է�C�����`/$*��My�u��#5߼�4��pF/���`�S^ �������_vGo��d�2����%Dq���CG����^G��f�G^M��u��g��{�$�g��1��/������C$S��ԍ�W5"��j��6e�D1
���L#�;��i(?Q�9�G�������i����2���W��"|}�li�q��v���ӽQ�$�p!ח���"Y8x&"��k�ItO�I�;�;H.ѕ�)6��cz]��Ӭ&]m�m_��  �������{���/ �(�ck"Ta�Q:�~�$����%�a�pJƙ4�����W�����O.�#�6��ˏ�l*���F4�8������g��2��B!�ˉ[����\	�vF����Oh�z|Ƌ�������l�knGa��@5]c��f��
߅\��'�.�*��;<��#����E��#�;�,���{w���Q:�H5��^�΃�`C?]�IC�:0��6�(4}>�:�Ex�u�6��{%�Y����{^?�'���ҟ|"��?�rK;t�������R�L@D`r���50� ���o �zâg��������^A�vvKH2pl-/Ri�����d)���zuY,St��K�"Ӟ1u�ɼ��t�QP��Hi�{U���'���r�k�e�� �|�u�!\:����2�����R�{Ro=0F�$��E:>�������z�h5�R�>�yog4�����p9����h���fR��>r�$G��g<��k���?�0��h�ܑmt�c��RyY�~�Ż��mۃf4��` Yr�Ҭg
Y�hK�Y) �S>��Ve�\��o�`���3�A�x2�鸧�'�M���Y=�ϐ�/�@a��C�d�^y=V��N�l޶�'�#~'}����(�盿ߎ>R^4�/�_5aOr��bTrM�w�X+ �����H�`ϫ�5r#̟t�`]����p������Q��RD	�a,�����swn���\i��_,��zTΑ��_��^��w�5xEL�hCm��1�R��S��wlB���&Ev������E��s=���U��\�h$�;��74�0JJ�j<���b5���{�V����e���̶4r9�
�;�a��2���yt�~��\oF:M#,�PΉ�ϸ��LɺCR��Y*[���Jj��BFIO��
��=��Vxsë�SP��
���18�损����h8{Kj}�����t�$��Ĕ]�%�����w�vHhyA�5��	k+s���Yz�B�T��gLK����\p��h�S�Q���5����q�A8�j{�lZ8,��8����c�ƃ�׋���?Z� �X4��F�)�z 6g{��m5�[����J�1O�;�n�T��3�A��AX��Q^���!�^�Tsf)U+A�Ddu2���x�AdXd��J���F(�2�^�AJ��[ʏ#R����)��>k�ޒ@*���$)�+"�~/z2��7r2�BT��.鏨Ŭ��Jχga��� 
�U$��a6"�a� A��\�6���>X�b�l!n��G���Mxk��j]�k��C$�[`�?Qҍ5��yp�����}:&�{���'�o��صo/љ�a z�*#K+����n�y���v�a�V��T�!��X�!�aS?;��x�m��l�5�y;��h��oH��SՊ���P!H��:ȼ=�Q���OV����I��<��!��_���  Ե�Vl�<�#��(n}TD_D�B`�R�����9��(�p��*`�������Jt��"�щ%��h����!O�D�r�}0���vs�2����*I5:�s!�EL9[u�L`�cn�*NC�����֮Y "�U��"R�� �Kmp���KG������ߢ��u�����?E�Om���$B�P�C�����)��e�a7r�jT�X��(�D2H����s�G���{�`�8<R�ˋ]�&�h!A�B
H*w���2$��:������~���Q�Ǿns��L�R*l��8l�A]�e�u}�SÅ��u�9�����9��l�L-�!rA89��B��T���o�� �L��22��ݺ�za��Fbļ��vk��"<��4��qi��`�ü���^��/�e9g�8�-�k2�3z���p����n"�7�eb ���.R|�s{2;��Zma�? �V��tk2���`�Z!���7X`Z��Ӈ�J����No�:��YƊN�o#j��?�J�p)�t����d���[~�9 ]���M�O���Gɞ�4�.�;�����c�Urj�nܖ�6�F�屽�O�V�%�����&̜x���6o� Ԫ'u��=AY��/%s�m7�T*�
X ������D��Z|/�c����[�S���p 2f�4��x?s���_*~�K�|�i�O`ZG���t"Md�?���_[����!t�Iq�����_ҖN�
�\��Q��R/l��Tƌ��t���ck�;���lkHB7�+N�tC�������v��	�\{�o��T6�k��n(H�Ӯw��8�H�]�?oj���1q�`	T8ag"A�ބS�we�(C��d���ѩ���Ȓ1�[/s*D�Z��׵kJ��<������dD�w�."�%����D,������9��g+,���K�CA%�r���G<X��q������W�R����Y����u���!�^_�죐1جe�6�E�$���R&y
��BlE%P;%����r��\>3iY0
ҽ7�w��������K��&]���ZX��?�[�,0�]Z_���EB��/8:'It�d}�����*��{�� �<Xg��o��]�T8�~m8����xq�쥬�ŁI]U ��V��Vf��GMibg�zZнɋW�K6N����tq�����b�Mm�|b�(S�Q���Ũtp�]�_�L���3���B�i �0�;��Fx�
:��C�tҔ��G� T�M$t�13�|k:S9M�f����x-���A�~t%�n���7�� +�d���͵�0X{@ß�Sw���d��a�4�����xH�X�M��Q4�:*�tJ忆�l�x���<�XdZ�f|���T�,���qgK`�� 9Mdc�M4�.To�)4���#��M_S��������v�$�oԲ����ӛ�*"="%���Z`yRӈ�W��&5d�q��?҆ �ы��'�nm�5�g�
���?1��t�V�}�"�U�Ƿ%�ǲ��T����$Hb���n��p�S̫Ŝ\g�!�F��7w����;�v҈
;S��D�h���ƾv.��p�2O@���K����!+���˵E���ƻ<�N=��f������<*�%&��⋓\C ����78Y�M;�͵���wi��T�
�G�v����@�+�������������Nw!��Dz/ 
|�;���6N��I�����C�9�T�[�Z�\��<��������`�X(��4����0`���#l�QT�JG�7a�
�R�uސj��w�$z��v���E��^0��=d|iB�k��u�}�ke �}��7�^4m�z7�� ���AkHz4^(>M�S�aӨ?k3-��y�߀QG5�<gYfw�3����=(o;H!��k���wr�ޞ�{8&wƔ��u��F�O���L�_F�4<��m7����(󮅖UWo=@u2#ٕ���ޜ��s�?+pH:���S�� *�X;"R틀
a��dE�o^%���[�XI٦�հEM9Д��{6��#di���Ce]\����i{��?68,�m�>���j~���=˂x2�^���o�Wپ�9Y�ε3.* �;��.V����C3��Ra cJV[���>kN�Q�e�g	�<�{bq����b���`pd2aN��)k;@=�	�d��C�NS�Gl,����
~���֭d�7G\��U5���q�w���������B��G�bƕY�������������')�6I Diռbߢ˄��r�3�g��?��o�Wkޏ|�ij���bC�;n�l��>ymmH�#[�_�]��(4u��p�׻�et�����|u����îL��sA�"	�ߙ�Z�`�\�E�[8��>�e*�e�	�z�L�qo����:D��C.����ɾr��%^�uy\뜛�rc�Ȁ�?�E|}�=��鵳�
5����Z�r(�|>WSp�T��'NHN�V���'+1|}��ʈ�R�>� �1�82�?�011#v+�NR���(�v�t�M�@4M���L:]�L��ZA��H����Z���;��QN� N;"^3���d�3X9GF���b���!�v�R'e�X�sR�J��aN�kߞM�IU$���A�~µ�[�S�VI��7��K�6�D�*d"��:���
�FQ��1�m]����
����� 	;�t�GRPd��D� �
�5	F��}f�1�l��@qU��V�9�+�Z��%>�����È��1avm�J���q���>��w.�F�fo�jY�����;���Z�Ɠ��#AfCT��f��˰f��w=L��V&,`�Jr�(��0U�a#D��dǬ��LM���J�k���R(��/:W�%��/?dy"��ť`�z���	Σ�_�"AA�����J*&��h�ð�vȁ *e��4�شRØ��bb?��a��k�и��Ր��V�RMTj<�	j5�gؔ��[�LӒ ?�I=D�p{N*+������ԉ1�1���)��ÍÊ�Ȳॹ�k�]1?��k�.Ί�pOH����[²JPZ@�ك<|Q�Ҝd>P����~\l����2�t�\�fY(';���$R��.�ב#[����7�t5��ofIXٿ޼C�������Ȼt}7 -lHE}�d��9n#�?��Bl��;�/`$}�*
�*k@L�֪���O��0|�z��|����o+YS��r�f���R��7k�M���cMA�k���o�x��(P;��pD��V'4�+�Γ�B�4R�8�H��͠���ʑ�h�˅Tc�'߸�rP�N�S���e��怢>aޟ�]ކzz�ZY���) �ȶ��`���S�JT*{���E�U,�+�Pyk�F։%�6t5Ę�;��&�ܕ���%���R$I1mּ�X���l�m��0S�F'c�@m��ޔQ���5 ��O�s�hJ'.�L���>�y�J^c�$��l��Ui�T���.jn�RQj�����қx.X�P��1���XD��X�x��`�Yp.1�?���.PS��5�@Gl�g�&�n�z�{� y�o�ƘTgT����#�$�h����mU�B�VH�o��li�-�jZ�q�'�Q8ϴF)*-����'����:u5����*����CbS�#K�������(f�����e(������"�2F7��RUL�`:ʘ9NK��*��b�]�Z��#���41�U��GÂ<M�?�5����p8Ϥ�]]Uh�P ���;�j��Uj�K�9C�'��q���h�b�P�.��}�|�X�����a���='{�B�RɌ�8o���~������ ��.�:Ae5����J��u��+�!İ����F��T�,l��<��X	T��ok�`�i~8T�ѻjw�����8x�R�����C�0V�����|��l�Ȼ�65�q��2�<�c0�����5�\<��؀��`�_0�h�?�ŵ8��9��7]VԃĚ�S�a馧v0��/�~ە�{�B�0�}����2tU屹b�Th5x����lQ;��i���sTi��� ����||ψ��H�h�틸��$�Q�-eMb'��l*�,m߀�>��qX�t��%��c�����w�b���ޣ+ք�e�AP�cߋ@o�9����t& �(?��@��½(������_�nog��s��8�ߺ���1#>���Ej���y�t��k<$�e����Ӎ��_�+�u/��8/��,�����A/�~9�E
�G�U'	*��j��<8�?1���#Ɵ��*3��%�+)�>
���˱"�AՈb�!���+9��x>����X)�WjE&�.\���1�%��%�e'��Ysx����h�*���|��	�fR��rl�OɠZ��P�])���ȁ�jo|q��E��������^;�M8ci�����ޡͬ+�Plq+	D��|n)���R@��ƥ��˖��=V�]&�gT�x��^�(����:�ö��i���P�{v���ХL�&Æ�U_g�썮8_щ��[�1��cݧ����Ħ�R6��k�|e�Ȼ]8���V�"Ւ&��i�!>aeR�/HpN�G����[�
�T7t6��Σ���s�� U���^� ��ߪ�V�
:����. n0d-��E|"vƖ`���2	c��ll?LiW����s�(���r"�������q@Ԙ�s���Q�5�d��0�A?%�qS[�H^tg��L��<�T'O�F�HljѶ��A����O� 7^X�X��6��=T��f5	�|^(���g�
W;M$�jMr,�լ0�χ�?���Qx��8���v<y����4o��A#��z���R�͸�hA���2��*Tf;�k�ȃ�Lm���TT�IhvJ� �,2�3��S�qU���0��wRA��r]|D����<�o�	D��XӹC0�/k~)���!P�C�X�!���G�e�d�I��_�^`e,wvg�2��SY�0�`��zw� ��1��8�滛G�m��6�M�⃀�D��D��!<)7��2��%�aS�>�l�~���$!c��oA��b!UoNu[~ˆ����)�Qa�J�2�Bc��.�#�˰�E����|9���@qF���$�EQ��6i�p�L\���ȗ���w�V{*z
U8�+_��@E'.��n�O�J�M� ^%�x�x���o�m�&c�;޹*'.d@w�k�ξB����U�w�o�uo�On������Ǿ��֣��8x7��Pt�4���g���O^�ϳV�F�]�F?0��۵���/݇ �x8��
�8"w��e@���n"na�#PpXN�6��}���N�}fa�lU���ҬH&lCX,B�a���"� �?�a�]��P#ey1���LzDo;��S�D���l���������\��N��?,�	53o��Ey��]hE[�o^)I�E���*��;�zK#}�P�KX��X&ҺbGü�l �[}�SFT����0�C���!�
����p�66J2{@��4U���$��Úǔ��'X�Nc�J�N�ߌ���ąXҁ����>�r�Ty_�DqSZU�+��E�u�Z�T^t�$��+�R����7����c�Z�`ј�T�����2͸|'6P*�9�I�ۯ���`�R�GsYL��T�Ԥ�U��$	��`�t}�N��E��Al�\�
=�-�s�)�>��n��9��&C�5�.�P���p�K{Y,���mG�M�bCݦ!���Y�,+�J �L'��	�bm2��w�3�cu�jc�ɱsQd�Ed�͊�o3}yA��g��g�ӘS�d��}��,��[pt#*V�RQJ�ڡ9jF�����*�-�reS�� �U���b�]b�0� ��mݞ1
��]1{ŧ�,���d����WYYŮs�8:�v!7���
�.��l��G��)�U[��ˀ��r�4��d��_qK[���T��@]���H݋4�%��sd>��{���9M[�^n�"틤v�l2b��K��6Wm���F�B�m�b��Ğ������0�H+}p��{<f��d��]�@�\LY���{�1�b��y�-��wA#t[�(7WfX�)�!�д��{�VG^�x��j;���k����!W�j�[T��XE5�q�?�۝���N�0�ߞ����o�r���j!�w'+F�6���io2����&�B�R��%��L����"�?�|]����F"�`cc���y��ރp �ݭ]�e>�=�ގ�I&&a4<�����ޓA�"��le+C;�!Y���(���~;�~bk��.n����?�=���"�^�C_�o>@��X�~P_33��<�|�^:οk|V@�{?/�+I^D�g���刕���*&�ꄖWk�+	�!�-�z�%u����3�o���­�+�C���L4��C��.N��.�Zr��"5(�N����c��\} &��<���W��?�:HcM�lD��YA#�;o���0��K�nŏ�ӵ!|�>BH}Qg�fܒ�ݧ�*Q��،hMz��d-K��ҫ�R��):j�˅K�9C�su.�#���X�=�P�h�o�o��H�5� d�b�7���*�j�=�b�W�D�?�4k0��������E��s�HJ�t�]��]EV�co	r��/�"HĞj��K�|.Q�
�u9Ԋ׌�(�b��hڻcA��/�bI��($4�ƒ�l��x꯰ ����"���"�����C��l�4�!��i��a���o��ښ��v/��x��~�Fܵ��B�V���-�B3����XJ��^W#� �~'����W��F�?��Su�]ժb|Oa\��`%+/���.��Ux#�*`����w��@\����U��� �����}���0��ّ>36�E�!��?43���(�D���O���&�H᠖d#�iȵ����_J{}�j�{�,�>��f�Ht_ճ1���@���|萀�2}��ȽT�����N��n�Z����!Q⚋;��4F��HʓX'�7�&�Wd�.�W�p��i�Ɏ:r��`�Qj�ǜv�����y�z_̣ݚͺ�_C����V18k� �Qs)`c�i��3c��=�f�nIr�o0�%�� t�އ���x���a�l'O|�,1��
-��O`��2g���|v�<��%��	��T�f#D;��iȅ�9*�~L��s�c'X�l�
�G��	!9���R��Ή̑7�������}�,e>�z簝X?���1o�}G��9)u_m�r�9���W-�|V��*� 鸜Q`��X�c^��"��J��<͞.�V�mW�M$�{`����h`�:Z�Zvo���3���&����Q6D�9��=���*n�[�����B!
���lC���a�|�=�O`w���"q���B�'�
�[��	����Z͑���P��t��R����-��Q��Rd%�`����*���իe-/��� ��؎$�ij*�Q�SJ��1Io���'`+H^�x6{jaq���*psbV%9ɪ]���!���w����]&g��^�<�t���D���ź-E�cC�K����u����G��7��TO��N�C�?Q��󔂬���*9r��9�&m^h��E����! �O�����I�3��]f�1��ɒ��4Wu�0t
���S3`V����p�F��0P T���W�%��c�b��ۮQ[S�L2�������y6�,�QQn��S��s4$��Q����2������囷26T���ZmJ��+��1]�>0��z&*��EX��7j�b
�0v"��x���i��j�" ¶.�4�N�-�E�H�E������E<�6��L�H��"�:���)VHt��A�˃��-[8�пr�H]���G�\���Qfx�qf}�|º ����m���Z`/��\� �l�d}K�j��>�:�[�{h�';~$�u�4౸�N�R����x��*�̐(����y��Ζ oT-D��⢄��ֈ�!�a;, P"Y��^域QoP�j�.P-^�Ӗ*�Z��7ˠbp�L:�0�e�y��t�^��!�p����q=�v
(�.������߱�.Y�#�K�l#�����	��3hV]��8�s��k�����$��Q_�)��e�c�G�F�H�4�]ሢ�5B��T��93v\ӳ�J�CjtYr'��r1o%�#Ъ����l��x�Z�
5�������,�����%�{���1{-?Ē(��|�0��d���Z��#��wn"�>z��������o�a�h��3{z%�r_ڡ#&�����~` UJ'��5`y -Sez["�mE��0�*g�JB�c��!9p��K;u�*]�ٜZ��ڛ��)d��fț�죟��f��Ջ�I����S���5PC4+�ZHf��V�g�)������^�<��ߓ��eB��*��\5�b����Y��\�X^�=�$���5�o����<�+)����L�]㏩��H�8�lڎ &*�@2-P6�e̿n���*c6��|���i6������1��	z��v��4Ci�a'�K�&RC؛��B��SFKH�	�仔M;s��1�H�b�{`�޳n��k�[�܏ۇY�XD�6�T[ ���}��0+FiZYr��e��Y�P����f؄��՛�K��(��K?S�}2��䜠�Vt��M�{rzU,��9���r�8^�����R�i�d�(�-��[�����*W���bz��nE�Ɨ�����4ٻ��ХIs$�g�L�E;g<&�͝��n��	�N��]����������l���.��"�"�2s�O9���oJ%��ܖ���S��=��=8�ë�����TMT�tʕ�����X_H�Gn�g?��0k��r|m�j
9�h�э���xL��o�8�X8���k� !{s�h������pcAab)c
�D��Hσ��nE7�S���Vq�O��4�+%�N�h� }�cO�%OQ��F���6C�K#�����$� ��5��!��4��9����oDej�+��N�'=@?
��C��#c��@ur0V!zf���p�<-������Һ�d��/[�����PGK���L��"dO��������`�K���$ۘ&��CKzt�pB�K��x�`��^ີ]�?G܌�/��e8L{��e_��1Y�|+l�}9�'@�L�4�OP,����"���]L�BN��I_gWx�f���Iq����p(|���^,�X�Rl�1�cDr	1m�m�r�Q!i/[X�!��dU:0d+��O0xn��C���Tm�FN��:q��"٥^!�aIg�����`V���v��U�à��ب����%)b܀�W���8��F�T�Z�)����꺐���Y�������s�qD�
���5�xE�����LE㰍�.����@���{�M���P�X�ԬXӂZ����n��鈸쏠�c�y��ھ;��`�hr��*t���E�؍ĸ�G;q�v�]��~sP6�'B��M93[�W/�+���60B񴐪�n�B���H{�h��=)�l*��Ѫ �0R�7�D�Eq��h�9tGZ冧�Ǘ��L�Jy|�i���Iպ���v�CՄ���Y���ys�QS���H�[�FDs!9��D���+zb^L9Ɖ����o��<=�;�z{{X��	���_jݓ� l��˙\Sx��_^x�y�M���T�l�`0$�g�>�6�o��0�h���J�q�c@Ou~L8��szT!Az,>3�n�5��9f#bvY_�hњ4�$ʾ͏ޡ�U1����M�/��q��̮m��ʌ��vQ9$/���	$f�-������A�i��$�;�Rc��gu8�_�mu;H��)�Nc�]� �}=Z��������h�B��j@����2��m�A,݈���C�����A��ͯ�q�����m������#�\o�h���5���9̤�+Ǥ�$@�\g�
��`ϣ}����ee����&��e�7�O��B���Ϳ���*��\��x.�Ş�%Q���g�'�|��Խ��������ތ��tW��o��<z��Ol�X�65�R3۾�-��8��iއԩ�#<0��D���֡�7%H������0���=J/U�l^�^Z���x-��&��~�KK
�>���H��Ne����k�v�[��{(Z�#�&�'��u5ۨ>"4i�T=&��q���ɐ�ٶP�Σ�~5�d�6Q��aA�-zQ��H��q�!��~-g�#W��F^�U�}J�~� ĨS:Hɾ���pPe T��q���x�"��\X�PhP�,%*�C���R4Ԝ�ʜ�h��J��E\��㯵�<+�Ӑ�B�T�.�L��׉쾯`�ԡ�{�<��@FRL�hp4�o���o��.�=�]��,�_�?�f�昉�8��KK�R�ɤ����#�6�*lP�p]7�v��t�Tq����:F\b)��
<��W�1�P��$�B}�u�ա��i��޲H�7e3��
�c`���q�nބ�.PH\������c����Ii$j����R�����δ�@o��A���m�7R���XF�?�� y�µR؅evx!z]�� ֚@��?��7$�-E*H�$�3�5���U�^G���Xi��D��5m���W��(ǥc2�H<v��1/ wG��G�?�M#��dw����P��x���4�2�N���<X��\����8�p���K�78X,�JJ��15��G�s%���q�*
�_T�����l@��I+�P�Pw;oϗv��tn��y^5��G�$���bY������ ��x\`D�K���z"�������'@�ї���w��-��A@����`�(Ep%_���	��Pe�l����p^RM6�9ۑ�,�΍�9`a ĉ�Fy����x�P~h��:�DLԠ�7��zB��r�\&�c��܉:
S��`�F�gIH�5�,�=�{-{�@�d��
��SD��D)A��c(H��L���r"��IU¬I��Ў�-���.~��;۟5"�=�Bp�m���R����hU��s���cQR*����#Z�=�v���x�3⛛CH����Hz C.Jɮ�F�6fI�ay+ yS�#C	��R��ur��%��� g���Z�b�몮�fR!��;Mm�i�Y:��Ǝ��
�9Q)�M-�Q�Ϊ.�'"�������?��.�a]��P'��q�`�-vE�w����q��I�f�r�1����T�m��ꔀ�����v��v�5�zG
̺�=�� ��Sń�*�9zO&�ꄼ����
�!/N3&<�h��nSQ�u�x�S��\~�l ��q�{�+MM�cM�'��(KQ������{��9-��~�tzg��_�r
5T�}D�oOU&U4H�0-�i���]|'p5�V�e�,QB��~G��U`&Q���q~��2����hM�o��K���+��1̑��C?�R�Zm�lg�$���?V��1R��$`��c����W�y}ô��Kl��)�	�����N��nd:{-��b!��3ѣ�T�:x��K�G2;����13aC-�c���B���#��lLv&a5<�/�UC��9�ۄ��PV�%[me�7f���}M#�M$y�Se��)�O8�p��*�&v9Ϥ���n�DnF�7 �;|� j	�A��-���~�˷��
X�%i�G�o:,烫h&DI*Ԟ�����uS�L�yo�a5��	�vI���P���������5�#۾��K�ϲ�'�wrU��7H��i��P]m�*��p��KX���B�
I훛i�h)������.�� �eD�{�(��M�{ӯ]�٥���6غ�\�]i���kG�H,�%½��h��S�F�� }���h���N	�g�Wg�,!�"8���^E��+����O�����P2�f�����P���4wc�wܹ��4g�s\_֠��J���ʴ���C��7�]��-7ӷJx:0�w�mg[ �=�c�I$h^ڢ���=���>�A�-�?��
W��c��/B8a�F/��癕��kL�����:����J��n��똣�vk[c,����
��}:mlýK�mJAaY��t^��� �4fr\�6��<���d��v�h���R��[��&�6�rf���[C!e]Ep�19U��l;��q�����7���f����������"`�sv���`�V@�t��a��&˕ �����7�Ku�s���bD�KE�j��b	(إ�^�A:V����nQ`�%��}6�Ȱ
HB.��K�:��Èٚ�?�o;�@>@8��Ȓ�%B04~,�v����[����ک����-t�>��#-&�bzL3��B1N-Ǧ�=��Y�.���tr�����pݥH��S'�c2�X�/�G֊N~-iC��)����#�:_�F@Xʵ�+cYsL��x�~/?�2�@���
#��g_�-S 9-_��K��������tS~�A>�d��Q��(��� ��z=8����ҽ���=_@ݙ���������h!��~v{�I����=֯1�+]�_%��]5)t�1¹�P���}����_�,ܑ~si�&�8Ɲ�t�ƙ�c�Bka.��4�{�-Y�!JC[�}/`�S	��>�I	�]|�Å��e��.��OkG��D���>mX�ҙ'r�Eڊvj)�W�_v�u �dDV�����G�<wb�����*d��g����e��jM�bS��j�(����E%}̃�ުK��E�Tj�>��7_��r����PB����
���h����sb�|��P�W�M�8d�@���%�lX:6ʏ�Ja%��/�F ����������=��2���2t�dX��4c��G1��Es8����p�C� &��a��{��_���"�['N����5���q~�H��c:1�<aQ9�@����{Ğ���RǛ`�8D,X��u��` ����-�)����m����� �&�&�������H�<;��F��� �*��Č#	���$'>Ie�~���Ґ��+��LVԌ����i�<A��c�O�PCat�#s�n��b�wi�Iw��%΁�Nz,���84�ހ�vV;~i��٪�İlB�Q`� T~��j7ca�4M�$�--V�]եA]3� �LH[����S��$��s%Eb�:��a��h����,�;Z�B��K���<��Ҭ���c�|��애���B-s���`^�XѮN�.��WW0�r6*N&/���ڞ#po�Ǧ��P��(�j�?���t��0W5/*��R��)���z�$q_ӟ;W�1i��<��	%)oԶ(e�@���L�������p��3mF�IJ�U@�ܴ����0�=	J81�Q�+�g�~�T?ǒ��}�E`�`3���z�M��$w�)�/���jyIP�Sb����P��_���/�嫍m����:��f�(��&٬�[H����qL��Nf�y��u�b�Z"8^Az�_�f�_�τ����I>
l�h�h�U($���m�$+��7�= ��R�	����l��_6���yDH�jK�K@P@����VrAx�¹�+?�l0lK9'IZ������:�k��rȉ���w��ݜ�*���C�U�R��o�M&��dg9��n��{o� >�o'Z{���f�Ä��؊6�����8�����1��j���/�
GF�{��L_h��i8�DM*m�P�RF��}م	Q��꡶�Ls�cSr���u�/,+�N����3>�����-AN��F.������}Z��Xd}�qZ�Q�>�~�L�5��P�8��M���r6��������
��T�s'A�z6��b"��pO�=VM?A��{t��|���X�9P�Y���|�۰ߜ�X%�L��ɍg�� K�3Q f���6�4�{X�����J��^G���ۿ�/��\I��6�,�ƥ�klo�8�$tZ��馌a��b-�����;��M0?�M��S(������Р���/��v�W��9p.�s�2�$�Pa±�����j�U�s�˪�"���(S�ğ��~C���}Tv4d�
T-��~+!���8c2Nݳ9��
le�p�Q;�_T�qﾵz������֩����cA�R�k4�M� ���J����Kb��	��0�]�X��b����i�p7�|nݰ�_^H��Q���>|c�a�A-�6y �?ByS���xt�W'1����q�P��PB:ǂߔU��p��6��γc��Y�v��U��:��n�~b �(?�xc.C��Uz��Y�JS�0� �6�Zd�"��X��|ZG�,���.>"5�h���s�Q����wo�G-�`��SkSV�m`,a��\��l{/�����;��H)�5%,�&����?ؤ\�y�ߙ||MP4<72C�����A������P{�Rk��|<���;nc���e�*���5���%[��z�:�R��]6[�k�>�}{s���vC�����eS�������}N���J�� �מ��O�Q�Z���2L�f�+��t��Z[i����j9���s���Ŗ^����z7d��V��/e{�������`I�^��i���	��ʩL87x�C-���m�[';q�R����O��#����ed��n8@4��W

�����~nL��s�͂�1�h0*�f2�`�a�yב����v�˓�4�L�w�e�Jߦa6���q��v�r����+���mS�-v�N��r���(����� ^K@�q1/��5�d/�nE�<�!]�K�����j.4ǅ��)!�ǚN;謆�B!̎�~(����J�*c�R��VxQ�,�N:7���)�lD��W��R��b�&:}n>�[�9N��A���$ j�>iEh �wS��^�����-pT���5c�Z=`��Y*���������c��f�{�C����s��喃d=ֹR!�aX�4���cNTB�@=[�(��\~@�n���b��{g��"X�������&�}�SQ?����L���Ғ���KO6N&%�>�����b�1$�%`�'�ߪ}�U����j�m�{	�����a�ѣ\�|큌wP���#�x���-x_�YPj\��P�rUӯ!r�6ѡ�F�7"<n�@����� �$ѐ,�@p�bQ�o���]4�')��_��@�m�d�o�܀`לo�)JsiU0��O����L�-�'z�{�C��͖���dW|�8�n��#���H:���������z̼��$ml��lI��G��Զ��B��5]6�G��K�*��u:�NjԬ���
c��'GR�qu��ڢ���<ǘ��se�S���ל"O�� ���Yj�l|?�W*5�U�| �]�Xh|v�l��Vt��8>�=S%w����:�"��B��Wˆ�'��%���>}���H��D�C�4G�j\T��b�T{/�fbj�N�K�� ����CP"�p��ף�R<X��R�6��Z�w��iE�0]�g�M�T˝Ⱥڪ�Y�r���~ �td�4&���]��Ġ�}����+j��
i��}�iL������xV2������l���k�o�6�Ǜ4��J¦���S��ϋ����|��u����	�C�~���T�W��Ps���#�����xͦ)��b-�ݪ���#�JZ2�9�� ��U�kJO\�?(���#C��pD����_�fO�o㮨�a9���f�b��)����s�E(��DY!��;)[�<]�uM"�VEn'����JX}�RJ���6����U��B�B���,�3(L����E �MC�G3lK߈���t_0g��T	t%}�Lp��wwai�N4*̇�n���ȟ�
G]���L���
�:-Y�)��iy�/��U�scq�4ə���ƹr^�����o�ҕDINN��մK���X;ZOM���_F0d�:�Ta�����9�^��H��燚RS�_�MmBR�R㎏Qk	lx���	8�i2�5%^q�������9���}}�S�5�y:!�*R�Ɇ:��,s��J�U��*9𡚾��]�8WҺ�C�<tP�A*g7���g��5;��y��xBk6��@t��v��
_�!��ԑojp�}��(N�ğ4T�Ak��y��˚-��W����