��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O� ` ��h��#!`"^��aP��v�P�"W�<!���B�|hG�'��g�G�h��6Y|Ia�$�]{��^]��6�N����THFn�Ū��X��u��'�HJȌ��k�ܨ�>7xD��x��~�X�erVG���a�1`�r~#�e7'�G�ge^�X�¢z�L������H?����Ώ��BP$�d>�GǙ�@E�*���j���W��N$�é���=a,�;0]�x�d�!eco�OZi�*o������2�A�s�����'1D���2���F�u(�!���*���C)�1��i�&������I�BB��_��BO$ob~�zd�TP5n�㝞����G��oX���ʩ=N=<qؒ�;M2����"�J2}�I*�}�gTZ#��f��(����z�}g:="P����������α��N��Q���x��������ǂ������Z�2��i,�_��,n��������?���6~;$�u�p���Y���<���9W!���(R��S���s;=�*f ��_�����}����,� }N�H]�va�^����s�8�"�zDP�h�1���(]|^��BO%�QG�3��U�D5� ^	�sJɕ"���8zMݷLLm`+$��:�7�A�?^y>�#�q�������ys�/�j��泻��͆�[���g������V� ���3���^ơ���E�ha�r�s��K�N� ��xlRcj"��<��&���.��7x'x�޳�@X9�@��	\`SPQ�g�h�|^�JY�� � r�-eW*��hiE}��5&�Ea>�e��q������O�)o�K�ј�Wa<���Ci��a��dJ���a����NmrM�P���`tL͹{���w5�d�I����t�����Q�#�珌{�.2�8=�4�V{u���`p��yQ�K��.T�W�n�{�����ҟ��T��G�j��M��$�:9��%=��Q�R:�O��XN�@bޙ�P��6���Z{�fF:!%7����z,R~��!����7TU)�}�u"PyPĭK���\q�!�����6��e�8R^�Y�C>���?�wqW�V��z,g%(D1����ݽ����fDϻ2p�<9��4��7����S����{�8��cr\���$M���WT4���gr��y;Y�F'����,f�$m�� ��)������f~�7���p#�<q��\9�F+o����EP6��>ݲ#I�ƛ���YMS�7�+��lM:�c�e2��׾/�T!]���v���� �M�J@����d������q)u�Q����y�ċ})���A���#�U��X$��Vt�D�Rn)͈���/D���3��#w�B��/�=�S-����:����u#9i��>ut���X*gݩ��,d[�>�lK�K��\��G"�(Ȥ��)~HH�YN�v��d)�2㿝Ub?U�+7���
$zb��l9_t��ĭ��o���D�PS�M�#ͤa5�NS�Z{�	rh�v�jϸ����p;�r56�,ӧ�&N�͗#�fNϿ�k!>��P�P��%T��\0Z��w���(�yu�<?J
�c`�y6Ov�9 X����IW�>Q�M��H�:��H\	P�J��䂿 ����C���g���h��p�0&�Wf��;�с�A��=�Ё"������Ⱥi�~d�'����a&��2��X�w���0���A���6
`�&X�n��"�7\<���W?��)B4��qi�P�~J�je��3�42���HFR���:�ی�%�Y���(�j"H��V1f��n[_���A