��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l��Hf����T�d�aF�ܾ� �1�1gā��T-x[h��E��edȇh��>ʄ���hPT㍖��l�U�=^��fw��BȎ.�<NV`����L����:źΖ@�ր ������*&���[�E�o�0Q����g$ʔ��L��ލ<-��~��_Ը�3I����]�cF�)��+�K0�d��xJsQ�&�g�Q�A�a\��͆���X~|�Uf�5qѸ�K�����!�>�6�����8�W��\x|}�X�'�W�Kn�f��R����S$k��JOW��80[��A� a����=���K���>\i��H_C2/KOB{g�r�z�ϭ���۰2��,�� ���L-�T��& "]�	f`3��y��o�ۓ�a�qr������Ǝ��dX���O�r *��3�$%63V�`�Y}U�r��m+䉄5=چc�!��\o��v���%jO\�_߽}!%��M���)�CO�ص�>�:�%;���kD�sd��A<�n5�s���Er��4��ߙ��
�G��T�u����f>�IEļ>��2~�pkCȤ�0Lj9��v��I9��=$�a�xa�N �4x�u��P}��BY��,ѽ��b��On~>�
n�	�x�\(�7��4�6]����Pn��F��xm6�ֹUW�׋$�T��ZY��m�\�E��v�b��.0�%ee] ��xg5lf�9m�$�|���
&��b���Ūh;�fJ1�3�T7/ֶ��q����>-�ÖB4@��?��B�UгG:.kk ��Z+�f�=Ơ�Y����J�oN/���)˃m
P�@��|��`b���8J�h��h˫�G���9q�ɛ�,W���I
��y��Q����T+�!l�eN