��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�3,ESA����ٯ�+��Ӳ�eHS� ���CD�,�eY<T�0?� 9G�ӑ~�7C�M�=6"h.w6K�����=e%�_ّ�L�'k3�؋U��³M�)UV0!.�c�f9!;��0?t�5�3D�X�[���.��?Di�
V ��4;��3�VFj�C����@����z;���8flG"�9�'bK�ǽŹ@_���2�b(tc�ӟJ�Yg��k~Dm&{�+t�.C�A��x����BZ9%�	��mvãR��HiY"�-D�-���cJ����)=��n�����/$�m���)�}��+prAaJb)Ĺ!􍎃�2�:
`d*�Y�]������M���ٍ�������n�AC���{s�����}⺩G#SHm|�3�����Xo��A~K�֙L����'��!�����gC43��t���Z���-f�-�UV߀F���\{娬6}w�D��>�����O^�1g1�S�4�T���L9��J���[,_�y�+ňwE�0�g��|���k!�-�����ZiRװ��lSӴ����۞̌�˥g`l4������)��SiMMy�r6�3O�N����ۧ\���3f󕘱�P������8�+^���b�'�`Y|��-�Ps ,O+����������C��}��U�,���i�jz�In"$�}���Zֳ�@3��5�R.f��?u,�]#`�ė��<ߍ���2��vn5���,��f#֬���������>~
/g��`b%�	�?�k�xT��)�� �n+�Ţf{���>gY�G���N�|��J�����-��p7�GQCk��f��N�-@s�o��^Ď̴�;S������g�c�g�#�'��>H��-��i���o��Y�X����F�y��� R��W�Q �O	b�Hq���� 7���c�x�F�*[��D�~}#����+�vە1�D8R��BȄ����P3������t�Z*�'�?�Ţ�����Y'�X���F�I�9���C������lծl��!�H�a:��a�0�Fmf[�/v�ŉCl�î#��_P=	(�c��Z2����Ec�ay�F�s��dA�Z�V��2P�����!e�v+�N�9^e��0��Q!��8Ӹ��8e�]��t����&Ak� ��B�����d˺f�s&Q��&..Kn��q�ޜ3���i��8��3���y瘀ύA,�~�8�N6l����ѱ܆�v�.��2��IN_���.��TY}Ը��d�9�[���qu[���|wВ�n�O+�ř�Ҁ�Q,������u�J�H�	�Q�:\�.D5|�դ{��y��6﬉�Vn�?�ޑ��x�����P/��V{o#���W6�F'�e8_b��;�g����7_:c:��!������(�q�����m&޵>':�Q�}=��5:}�OIp�XF�㍿�r�h�#��M�I*Cf����+"逑��t�IҎe`dI���W��KA���i�'�s���w�A���r,6���z�µ��k�%р��>����9����=�Q*�����p����^�W!t�F���-uE2L��G:_��/���.)�����FA���e�l��γn�V ���n�У�0�p��[��n�~Ԉ�I�=��I�B=A@V\H�pt�|���jU��,�R���8#� ���  ��;X:'k�a�ț>�7_$C���&��j�+%?h��X��������b^��I��h_E��I���&���t�b��4����HHr�B�;9b�.�=͙���>��s�CI��R$��̳�J0ĕS�4U��@_��;�\,[�g<�a��A6�Z)��Y�s+$��;u��vV�v����y�� �ӡi(��Q\9<p]��AeϷ�p���u��>e}����+2S�
�c:?�ǄW�Yc��3�Y�58�k/;o���k5�����"Df�h��ӇJ�q���MW�ݮ7-<<[z�p��I��E����lu�'�J*!�r#�H-__�e�H}\�S��a��B�a�ڤ6M.���[O�Z�n�g��e�f{��ﾻ��;E�����m�VC�mc����6�o[�/��1a�ZY��]i���f:���D��F�D���f׏b>�@,u���)8�.�՗`�c��� �/��6�9+�p��!��v��������B��Mg��Ys��r����O�����,����Y#�%7�㩡�c���R���$@���AB�Z^���]�F������C�ºyOv�(-`��i8�:�d��yˤs���JC��u�ыG�,a`o�H�\+��s2Z6ޛDr����u�`-ot��A�ymU��O�!�;�3u�1u�tr]�y�d3i
��\�I�WT�F~�^�]�{��) �#A�|�凪��k51E���H��c}�e�bM�RC�\�طzW���;x
�.K-��+S��#��L�F��{���bv�T9B	�Y�/+u\�^����Ы߅�7�8~*ӧ�R�J��a�hZ��������Ɏ2f�-��P�����l����5���!��%��eȋ:َ�� ]ǳ~��:^mt���J"]L)�<5v�U����:�<ޓbw*����QI����v�-I��V�aj/����D@��t�*���
���"'�n��>���Ldh{ ����=���tsu�{����zV��f!�_�A�O�w۠��o�@s����˖���o�e��dd��Ym �I��JޓS�?hW�<�������@��8�ʵ��*�/"$a��)#�Ph�!?����
��|S�t����qUf,=��c��gɕ_#DL��΍'K�=G��x)ۇ��q��#���gT���S%m@��hQmh(��$��>�z�T-��j5�O�����̿5�f��Y�i��A왿eN
���m���=��j~��wMy�s�vb�\7����וּ�ˮ|�
WB�ݻ����Ծx��iy~�c�o���c���\��O�H�ުf�y��/Lּ\�c)T������-�����Cs�^2�nyl��8b ���bM�(��:�d�1��6�Q4l����M���4�����Xt����h��0��﭅�Y�$���� �`�0EG�]�p�Ý�h�L�7��Hΰ0�h{�:��:E�n����F?���ʢ~l�1����x,��+��`��e���גx�5�꿣����>ic�B$�H���'2�M3b��F�.;��G-3���W	��d��$�BD�#p��+���YUN@�6��9�.�'�9\2��q�Z��z��I-A�=!�)��x�)e��}B,���cT&������V&�Y�ީ.k�9e�!=��}��jU�|5fm�D����4*��%�INog��B���IA:{�C}� ��k�Nw�0$JڥC#G"&�����D�̷�U1VG(4}"  3J�6ż�PF	�xk!r��������4m��eK�K�xvд�e?��}�����n�M�hC���Y:c�����e���̴���\p��)�8�u5}q�G:�j'��9�Ef�0|F�w��aQ(�;S\x���Nw��l@��1r̩?L��8���&D�ܡV��5)8�m��g�� ����؇��f���qI�W�"�yz53]{(kV�Tg�Y��:Z�Hd���/�T05��4�Åc�C��F$�jNfN�j��T-b	���w"�� �H��&٢�͡?���V#��|y	��Tڤ7wъ��8e�B��$}w�V����$��5���.nhn�X��6ړ�εE�-.n��Cg���-�����y_}�D�,�]�HGE�|A��O=�FTa@M۴ࠧ��N��w]c��p�.3˱�:�@;�ϥ�w�5�t]Y��hG$1����ʬ�z�~�:5|۽O����3�3�Zf�m]�����W�.�P$�5��c �'��yҾ������"Ԝ��:�6rfM������0����}"��pSI�psG�)fW[z{Hx�'�?�^�g�f_|���h�\����E����F���_���ᥠ�0V�"��,��IwO\�B&?N�J�HU�
��6�?JC��r{i��JX����l�Nhw� �W��@n�x��P�2�m����p����ֆ��E(fS�Tƚ��S���jI��ŝ��U>����?��Uv��i`,�N�Ed���>��A=�y�}voB(P0�DN$aC�4<��m�4�H���6; Zh�;�a���{���J�Ka�O1���ԡ��d~�hVy?v.B�X��!�[|���ccd�ή�uc�����A�n��%�[5<њ�EON$ԕO#�0������%鏖0�_/�[�Xz4r�W�Fw�M�����jZ���G.p�Uqڴc�S`�4�c|;�5�� y>
�<�Pql�ʐ'a�c?��EOĸ�
�}�
,q�x��0ہ�����*fM���G����ۺy�e�VՅJ(��̤�[b�XtN��[�:���ſ=���亁>��,J�
s�v��"G������M`י��-�L�NR@�ч%G�Ĭ�aV�*�D#��hr�
&���WG�1��W��!(B���\����C��W��8��F��?���~;��33���%7�rI�B?�g��3y���������"Lu#�1��{XˮG2k��=�z��\i�>.���Rfo�����!M��ZP�Y����iy��!��&/G�e�jLS�s?�J�Ī�(����?�xĐ��$���1<��<�2sLR��`9~�j\x6bI�)t�j�Ԉ��O��n�a��!���6��V���K�]�Ɗ|�s��!�닔p#,��<x�	��n���^�DKI{#W��'�|N�m�2���v���V7�[�d�� Ž[�h=�E��	��l{��&��L��<ۊg�4Zul�N�����H� ����L��D&�G΂�l4
��R'pU�5Q��}a���T2�N�)0R};�g<T�0,
�&@Y4s�;�
�#��!pm�����6rW���,�Q��j�/��­��ӧBLĞޔ�m�{��>��~���,���8�Y$��<�V�e�'����A�N���ĝ@���^��kOG�'쉿[/N��꠸�{���l"J�B.��k�h$�xi�Ta��6%�՚�Q��W���y��|Sn��v��0�YE$��)Lw���dx`�������d=Bt,�:$p��Rj�����2e&��N�E�okbh(k[����I�g�/}3��+��1�/�g �,�Γ���Q@���6@E�ѿuU܅i�j�!
���qwEK��e�Ps
]�y$lV2�\�I�ܫ��*��� ���H����['J�㿋$DYoӘ��w,�+k2L�|���`��e���~t07�;Ik�o��˝�����W�:/G%W�u�V�~�$)�8
u��R�#�]�;������Eצܽ7�@m�}-7>��}���z�V�_a���_�����3�m�⡆9�$����)��7����9�L]�h>�t2�>*H�?�)�4�2��������Lc�n�i���8$x}�_�m�l����4��љE����
	��#�QJ��� �e�������1�P�碻��F�mS8Jc�LP����}A�2�Ȉ]+fX���<��t3�W�H��{:�?�x�}�<��P�ϕ8}������Pn��W�v�����S����C�W�M~^�҅FA�XX;�:���b��u��o�t�q�(am.HZ���{ �/�M��~h�O��G,}�JS`g�ݼE9'=+䭳=��������AT��,v���U��ƹ^��F�����e�K{MF�����D��B1;����=�G���bړG�-�-�<��d`v�_!940ɐ#4]M{Qud�&�4�5��nZ�����QO���e6L�L�w��:(2��#�;��u)e�Pd�������Kkq�P�nJ��9�)���ئ��+&Ȃ����˙��tr��,��o��^��GIIr�p: �����ȺA�v�A`)��u*�`= ��\�<���&e�0U_�`�/&Z��.����`�O�o�RCP�d�)��ps����V�Q�����A���T�E)aW�"e�죌�)=r;�?���|�腪7��%n��ۧ���'�v���
x�MD�;fu���3�F);�;U0F�v�x)��(r!����I����@m��y+��:�H��>�����ꤛ"CK%ϻ��N�k1�tP�����8x����:����M{\����~Ol�� �.k��'W�c곊T�H���:\]���p��}Wx�.a�I�e���Hu�	d",c��C�� ����^1�1��k؃�k��i�X5�DӮQ��:���OY�e���jVC�?�_h"��/�A%��>�������`a�~�C�J$�mDKq��gU�7mU��9t��9J�����䩮�m}�?! ��j��ƁS z�]�K"s���l�������w��`�oS��M1��~�n�}�]�RZ�Lp�:�E(�Ă���+(B� <S�07zxdyst[�)����>x�\�YcnC �Z`4���9|�kT�qE���\+�*�E
`@�?1�&	��Ԯ0-A���u�~��h�I�ܷ�45��<��A�?~δ8�h�z�|�>ȗ��d$&>ț�����z��"��-�Ho��8bY��,�R\��8�1��ک�W��=�ܺO�~
��"}�*��臥�rG�G���i����u��ֵЉ�5qǭ���H/���$�
o��B�tmB���cH�()�6Hl��EԋD�(6[��� mՒ�}r]���b������֛ �觔fU�|�v��*��!�p(35��:��o��U7oۡ�u'�b�� ��x��BbG�}w?W.��k�R�B���k��:]MX��pB��yO~!W�Br�C��4�{h�`�q@��(2��E�����D���ox��2B�z�@[9=��X'D������9'$�)�P���q���J�3||�C��H.Zܡ�PM�ݠ]�i����B��2&?�^�Mk�t
��Óc1�Y	#����ƁN�AF�H�}�d�QO#I��e9E�4凉}�E%x���ʩh:�~�g�{BV��,�� J4�'>\a�!SHE求�P��	'�r����g}���� W�2�y�A�M��O�d)�ު�6�$�[�0�Y(�*���̺������>���f��&��z\��`��������h�����&�E9w��C�n� ��f�� T��B�&�#T �5�i}x(�ܓ���6�T���wj5��3�Q�Z��0�>���z��}AdEԬ.�WC�g�N�c�RLv:��%��\���7-"��~@)��0i���z]��C��yRgb�{C��U�������� 7����vkU���.L3�LS�~������6�w��DW���쒡C��Oz�����W�җ򳑳���:+C�6l�Xw/T7��,yWc�́�Uh<?�Ԡ~A�vG$�%[�@	��T�K��M�Wʩ�:n?|Ld�x�8����$]z�T�|�u���a������NE�&�t>NC���9'ȫ��W`��V�TO=(��hy��T䨄@|�p�#@(��eՖ�Su�� �a��;