��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��E���������ڄ�p,�)��Y*����H�	�W���!r/����V&�
I����k���W	�Ś}���`Td�lh��N?o���翿g>�4�2�α9��E�ƭA��J湅Uk5��$���Q' �������� �9bZK�������w�k�����B�6�9�F���R� qDv릁��T?���P�H$���8/����ȗWG�M:f/V�]�,��x��໛����H��_GJ�^/n����~��hP��5y	O�8�)b����d�.�7��n�EL��H��"&�0��8(�1����<Oj�r���R-h��M|�NHd�W�b�kYތ���7X^���(�BH,�i�Z���}���<b��Oy�h=4��R�f�I�P.><��J��c����K���=��=^wlkFƋA��h.�}@�% Â���f�z�]Y/������Zx,�w:[�;5���>�c�-OwL@��LAva��ټTB2�ݟ���&{[i�jP�Ai�.,����WFv���@o�d��᪝!@�����>�z#�\
�ĭ�-��Y��D��+��rԳ=���ʅ�To܍]o/���o��yC[d�fH�?��Z��=�Hj�����Tp]XHip]IKp�\w�-Y�w�IF���%Ps*�����v.g�ٗ m'1m� f�@���?Zn�s���pD��]�m_�=l�j�za˴>$��>fQ��h�x�+� �6T�)�� %Z��V&V���@�X�����q�v�.?<�}�<ٮo� ����-�gC% G������[O��e���Σ��;U�ĸ����踼ŃA�v^#k��<ZyQ��G"� |�q� S���ݪ�|�CZI�M����D,�4��E("IAi��7X�fV��_јR��K���e�&�E&��T~NՔ�;�k�H���c����䡛`�Y�+���+i��K"S~�kzD��ݩkX��ӵ�La��5Z6�P@/���+2ꉽp���ƚ"p�G0��_��ښ�/3ժ���o����N��.1��T�����������r���hP�c��ȫV��+��DM���I���� K��]tQ�0�I ����L[��=r����&yi@2 ��#>�89kQ���Լ�ݎl��H�Azf����Jh3��]�`kPE~#ӍU=�<Uv�g�#��Z����9eS�(d�$�N�6�hQ��S��'�8��qo�3;Kn�!Z���[���̒#�9N�v�;��e�bo�Uz�F���s[�����
ݽ$�hO�*&:��J?�yc�>�mad���+si�m��� F�h<R�r0B�k v��t�@�!m���;�4�V|�q��Q�H[I>��_�t0%�(�ҟ�"����P]L]{El�<�4���8�J��љ�S��.3Oo�'�N��QSh��3HX�撦um=��?���1r��D�LN{_I,��֌�^R��rP�KuQg����Rs�}8X^�6BC�n�2�C���fs^J�m�?BۂAh��׬�,տ+��=��!*��xm�W<Ę����O�5\Fx���9������,��3�-P�,��x�B�o�?�&-͑!�C�G������F�B�wԬdp��iϡI�2Č4֤��rʄ
࠷�<��y���8=�K�x��N�G\'g�;%ׇP&���@I�4F"�6��O�V�U#�^�/r�_1}2�R��B�> ��Έ;��'
@��r�^�"���n�7��>X�!�������6i�U%�;_��\��ά%E����D~Ūv]�dC�xt4~�>z�a��.�a��2ߦI�
��q���$*#�Ę�UDS��U�u�ʞ���ץ�Oj���g�����O�I<9Ac�ܮ����#���;�x�#
�S��4�'\�V.(��r�e�5�
'-_@Z
l$jJ��<�%������I��tI�Z�㉔���
�0@Pw��
�V���rA�PV|+mDlƫǛ��8�]$!r%�rݢ~C¯X�z������~�[`U�ӝކy[	���!�Nt7?B�LV	��L&��a��ow�gI�ۦ�O�RY��/O	}*o�՞]�����tJ?q}ş�еgU�-�K�l��"/�ո�i�m+�m�\r�GQ<�w�.f.` ��y<}��v�$[�N�]sڭq� oJn�r�oW@�	$�E�>�:�s�i�! 'g[��R8aj��@�wi�GM�&U������B�����-�t�9����<�|z�R<G�Y�(�IV���
J��n]�y����
Ɇ�Xi�At�:�tƨ��&er��V�J=C$s��t!}謉i.
����n�0>���]9s؋�����2�����>/���PJM�P)���I�]'?�ք*��{k��ǒ��z>w��J��ث��V�t'b'����s�(w9P{Z���%iJ�7rЙ�R��Esi5aqrŁ'�!µ[QZv1 \��5)���t1o)����%CC:\be��13pr)č�o�릮����D#�M'�����ұ+8}^��hT�&b�'m���*Y��6T���� �qe�̎G7c@�π��x��/��|���Ttz:e�����1���`�|D}� ɟ��M2j�/L8)32U�&8�e�O�;k�׍�i�j�=�~jmz?��:�l<۠�9$�EjGEn�v����߸�l�2.�cxY'�YF�/��a�n�
	ȋ�������:c��)�����ٽ�~�)�d�'��ϖv;2a��0*��)���YAdN��!�8A��3��'r��G�������������:���w K;{���N�[�=)m���L�T���W|Lv�b@���T�����zR���퀳p(�pÏ��sCS>.g���7�{`F���0��+Ф�%%��J[U��>l?8b�.�����aGz~�,oDh#d���<.��[l[r��s�����g�9���^`����?�ɺ����9�?C9�`����ܷ��`2���
���s��Ph1@���	@S�����Kfg˻}���0��L� ��|�&'���B�}�	�u^����&��&X-�hrK4H�:�����c��B�M�Ԅ@Vjk
�z�ĩ:��r7{�H�2�]�$g���F�;�(�%fT�'v7��u�J��<x@ԖqC�zaY�}
��L�7Z��cvٍ|�6V^�̪/�hiA'���,�^�	��e��s��S��D��3Fso�+��7'�b�����C��Z$��Ѵ"�@�Rt#�M�ws��_@&�Z��ع��V��q]��:��Ɠx{`������M�,8��r�IQ<e[��-��u�b`0-Q�V�;��o�M*�@��\� �;�R�hx�@�C��'� =�.T��v�b^�=ձEn�|�L���}=`8���6LÄ�{�����\ɑ�N_P8Y���@j%�J����'�M�r��d8�cF��m�Ȧr��"�t�����$�l��[�5G_��G�[#�o��&��QB�G�0e���!G���=ڣ�!�4�܆wڷ��S�U�;
�R�xM�y����W`��nM����]�a�h�E��*r�T�\��C��œyC���ص�A�Ƈ���W�SG�Q������@�;���r{Q^u�趨����1Js �<����ʈҏن��h<6��UW�%���]�^�.;�_�#�J���B�LF�'�&yC�k�`����X1�a��-��~�tw����DС��Yl,�m�p�FW�E�vbh�4�`��0��.`�/q�mL���p/-�q.�+n-,�>�NV�[
�-�GQM�m��H��p��+U�[�aUU��	����:���P���`�
��b�������R
ګ�����n���d-!�Jϖ� 7��̓�&�\f?�(�s�$��&�L���p���l:	C�hQ��>wV��"!��*�{����9�I��)7��l���H��C�'����I �n>MWH>s����#�l�Y~��͝�1(�����ċ4�ꑡs��6vx�]hAh�P�j���Q?� sE�A��l:��x%���q��T2����6��O�[HNM#	^�7`��rjO���BZ3�����O�2���N&�3q?���)R��|�Z��V<~Hņ��˝�"�J�J���.n��$��į6�g�D"��=Xc���
��-��A>w�^\0����B:��#��-��i�)qa���˻{(c��?f�Lt�ӧu�I��|$V?"�Fd��Q3+u���7p4������?x/_��}�;OE�#�.n�W��/?ع�;mޚ�@��3�`l؊��>���9'.�+���n��9���8Y�,��J4]�1F8	}c1ɿ}��F��F����u�~j�f!X�u|�N}rd��{���k^eQ�`StX�<���iI��g�͒8�.��H����V@?������P��r�R�0�ǖ�5�(RW�E�頜�Sè����q�n��U_Xv�e�|�C�6ö��r�ʬP���P�)�2'N*B$h �� ���a�jh-e��[�R����0�d�1�69�^��uܲg�Xy�M��/�k<W�������/u
�\�����SW)�@�m�H׺��Ԋ'�q�D�F�m�Ļ�D�wd� �Ih�T���Ã��?b�)騒�m�=_c
2�<�H�lx��_e�,7C�Yqj\vVU>��.,�#-J<�^�~��|��e#�"q�@���>���K̎��.���.�{� ��q�`��^��ʻk���gq���*GE�Z��4������nk�^�;�WU��ͨ���(���LbYZe��U�>��#Q���d�2s �Z�z���$`�,n�~���� Jg�;T�L���;-�~�蹄�18T�w'�˦Ydu�7��/�ń,)�r�_%|3!��LJ=��$���'��)��Ev�]����Ƌ�!Yz�D�� T�f���2���
��J�O� �<,{���P�8�MF�FGHnL�c������&\�?��	$)��f�����R[\�Y�����5�����<B�+�O���*�th�י�ʶ�Q�v/~�C���	X=�0�i�-��U(���M�'\%����x�)�L]|be����G�)���,�S�qШ�o��J1�T��Xw�J�S��ľ�#3qo��;��V��λכ^׭n�A��?s���7~׃6K��4��˭�����л7-��A�b�K��AH44�χ{���ʙ���>��Xn�.(5�f��$\iK]x���|�i{�l9�'�(��,���8�r��T���i���C�Q��Ȉ��4\l=@�s�֊��g�Վ'.g��!�"lS�4���6�-N�ǋ�qc�gh������T�*_����&�X+Sz2AP�*����e��&����_|�&�j�nxǟ3�y}���	���"�����	1���	���=qh����# v��A���z^�U�/�q�`�#c�;d�<aU:�(s� 8�Jչ�Wo]��k?^^fX/������5���i�������6��=1rq��֏�P�[P1�<��XgH������]�A��*�/�k��~}d��Y9kť4[ذ[��=�l嗭j��X��^3��}�1�Y�d1�tb&26y��^|��ӌP����W��)�Pw���n�v�<4h� k�+x��waxC9�\�;��H�b��E����G�ǭ[�� "*^�:,����쪪��-��Ѝi�m]K�-����5q�)0�H,x�xN�ױ�+�;/�7X���5�O�N4Mt�� ���~g���������dzbǉ�����Y�Fq���gpnG��q즒��nʹ�m�0e�,tF�q�Nt�P�r)�_��>:�u�Yn��T�l�a)��8�0Θ@F(۬��+�M���ۋϷ��F�k�kdG��/s��!�j�3>�]�s*%����ar$�E��S�Չ�d6���:�����'��H���D缗1V6�Dr�oؠ(���`؏�?	�w�݋K���T��ZkgtƤ2̉
���+�'���=G�̓M�����M�k.Bm) ���Ɲ>>���+�ڄ݅߅a8!��9V�dɊ<�����p�O����u|�$ �%
/�N*�@��Q��S,��u��À1l�%���Z��V��X�G����=���\��0 6{;c�����d��Oڹ�ܕ��}���x)<�fE< #����rު�mg�։
��D�zb��[L\I�F'�9����xy��́��~*B{
��yb��jg%��0�w{�!�F^�viR�u,�|Q��&��4\3$ �)w+}����}�N?
x;��h��(`�x�S��6�_� *�aLD$��l"�� �E��ˠ?�7���Ľ<�>ca����l��hNX�6+7e��������zm�F� �"�KJ�X�(+`���LR��Ј�R݇�=S���k�K���0�,4���o����#����,ξ�v���!\&������~�jv��v~��G`:}B)w���b�PѶb�w*�M��GEOM�����蚄_w@���,� �it��({)��!�&P�`�ýɮ�����k�����)�x��Io��pc��� ﹶ��vE��7��~9�5@8�2��M��)�CE}^���i�w��-��ŎNWQ��,*P%<�U�n��l��w;�&��D��YW��B^Qo$����� k��׀|��.|����F������/i�@�����3��SigoPį!���3��rx<�;������U6'��m�#+A5G�y�-�<U���� zPة������� #0��}�.��!ƃ�`i�\�`	��2j*�Ȃ�J3�J�T����Ӛ{�7�ŋa<V��1T�$�����cH��eܚC�=��Ǚ���Ln�/�<!Xp���xb��]z���,�W��`Y��ݺ�do��NN��h��GG��$�s���sط�m��>׺>3!�!DEJ�g��U�4NtҀ�#�ϋ�м*��(��Hh�&�1]���z��"-|y�N
-2\	���	%.���k�Y)��zg:��M�u-Ed�	�����F@$˴2�'�i^�K2@��w�ދ�*<�S�����(Xv����/���p�$^Q�H
�qeɀ��#(�e��x^:7�4L�k�V�=�#X�@֐��ѽO���l�7`��2�W̰��:r�)'����_ʞj��Mlz�}ȡ�-�qFvZ��Y������&m@�o����Cq�ΡC�9��ssIn0WЁê3��]��Zoz��mS7���?~U�5Ў@�翧=�`��4:P��k�K�����=",#ʼkr�Q��a{��η4;GL��y���\*�W�`�m];�eI"V`����Z�I"�L6@���zuB�iFtqO���
3C	Q�	|(�)�f�2�f�b���emp{�H?Vz�e�>`�2-z�^��������W�+x,G(�s�RY����u���^U>��O[�2^\������6�VO1>И0��ǍgT�ɲn�zT�1�V��x	{�P�Xz�w��Y��V�il`$�گ�0�R
�0��@�KI})N��D�i���j��H�A WjtX�K�0Xc����W��yY�郂����Ez�J�s!��n���{��"ue�Th�v����� NC��$�'$yhD�-3�Ro+��J_��GYO�O0<3Te�����5A�[()�F�w���3�≆
Cm��и�WXӕ��N����ARP��Ot���,�=�ٴ�x�(�H�U�W~��(���M�c��,T���?�s�7��	Ty���aX0ý���]�&tFD����pd�$!P����<cWd�[K7Δu~b��Z���R�����%��=�F������L�6D�w�/U�7����U��~[�T����T��JK$�4\:"���5�����3 |�&��d���_�J������p����q��`�Q	�}���څM������]gL����Gz�}z�]tUV�:������W�AɿB8�;�S���.��@�/ѤV^��ߩ@)����*T����������{W��6穄4����Yu}=��Oj�Q(��zE@��
i�){}��m�EؑXX�4
�
�B��:�!7���G�]�#`�ݗȩ�����9���;G�d� ��H��/`v�s��F���pW8��޵�1.��|�8dm$���2�fI� k�Q$�I{�y�bދD-Ӄ�ȋ�x(�^/h�-v����(�_���/��[��ڭ�%��R�۱���5Nm�'����Z��~VI�J*7��<�[����Zo[T`[!����پ�X�^$ߟם�r�����I��/vSo�NUϺC� ��%3@ڊ���ݡQ�HW�S� ��wHX���-�o1�QU,ߖA��,�//O�b@�������Q�^��J׷\0*x�U�9)��iQq`�!K�ӂS� =��H�	�i�4�t�2Z�Ѱ��6#`/���؏D[M��]�hg��!ӆ�w�d~�\)X�>y�'Ǟ��Yя@�(�~��I�ޑ )f0-��H�&`��r.�dGMciz&���
a��ʹ0���Q��C��᣶z�8©����G�_�[�WK�nRc�������Na�
�F�b�B�3DC(b>�}����Xm���X) C1�/�8��3&�X�mΆ�V���z�)�Ĉ��Ye���53#yׂ�d���u	C�|m�s5��m+�Ƃ�ڻiK��[��SK�-g.ϞvT��F�X���]\Jv*òӢ�� �u�R(�G�3 ��Ï|�{ǭuS�b!���),%݋ �k�NmDw�󐟙�oXq���D]�a��q�Bͩټ��2��,��M
r�V0-Mһ%)�\��yA�8!�u���P&d?�k�S'=hW��ҝ�7����B�0���AC��r*�� �)�D*B�H�K:��z��,��֚�f(�є9�!�P�a}��DŘ<��]l|��=u\`)S(�ql��
V�)�A6�Sk��U~��mmx6~��mG�N���pW�!iXF�^ۊ2����4�C�\L�X��$�π�LR���������n��ZQ[�� 8:d�����P/���g�mE��7���*34e�� �c6��a���*����DP�x"G��/�.���q�_p�n4լ_��������̻vaHd6M��tqƑpe�����B����R�~%nH��'r��c�Z��M��?�[5y��(�����`X,�#�6M�h�d��.��e��JoJ)\,��,��Y�]�ij�5��Տ@�&����wa��~�7�5G��R��˭��}�H�|�;�"��Ř��|�t�齆��9RVHǳ�9�#-<�zN]㊻�w~.�mB��^��cw�e�)���o�ϭ��cÂH�].3	�Ѣ�3[���+�f��e�M���(�W��	�	5$�1#'s�	X����v���͂pF2���������E_���5b蒍�n�l���e˜3���O�ڹ�;����z]�?�#��0@����˭Ň���6�M�@Y���吣�Ok�6{R�aM�"s�� q�3� .��#rL{TU�W�qut��V��{My		��;C��X�Jo�s�,!U:����እfJ�U�h�VK�A�������:���g��U�E�Caz��6̌�BJ����o��Fa�@��	#8Zۈo��Ӧ�)�/C0�	ά��V&x�n��.�'���3^���}YȮ7�cí� ��jT2
x1�J���猹�![�tG��`q��QM�ܓ��@;����6~�k��pK>j����-Z	�Ff	I��t���T�QH'�Ei�s �¨eh �W|��:���^��=�w.}g��a��K��'K04�gmß
S���҅0��(�#be�Y�h�L��}Z��I�}KMB�D��mm`�hn��F�6�������?�Uވ|L ƹ�1���|�t��f$(�����kr�nS�w��=�51�����(K�Dc��t������y���Z�e}*M�.d���Ω�6sZ��^L�%�AH ��-J��8��)w-�+z����.�4�X��W��>vh���VYتAX,7��o����/�ǻ<mA���?|d�Yw�F8n�-���X;д-�A[-q�V5��~��QNNm��@��O)y����͸��s�dZ�B����6��O�J�P�ƣ>`�EeF�"��b��W¬��;t���3�RY���&OW���$pڐoZ��MS���oD�Q6<���f>�Ҫ����Ώ�}�7��QwRI��AX$_fʘ�,*���;1�jD��/�0�<D3~�0m�'���s�TXQ5ٟ����|���N���a��m��SŨ
SR�a�"����\����@q�ܡ��/�*�}l�E����ِ�v~���z[����X�?]���5��NGI[�$W����
����|��$\��i�F9�72��vu`�H@,��H���W�eǪ�W�@���u��2c�,CB��n ���δւ�9�.\|���Bf}l�+��$���\�A6/�碽J�������ĸfn��#�6��sU����$c.��A"���}m(����D\���X5|�����/�۹.�R�� �:X�d{��9Ri8k�u�Mw'�����#�=�^�������tr�FC!�/�M���3��� �na�W�B7�>�8��s�-��MN)�����
�l'�7,�]z�V�׿�H�G��}1��
��L�k5%WƳ/��Mh�����x�bmJØ��ҚU�x��[�oC׈��F���8O�b�e=E�X��/vNM
�[���p��OGB�"K�C�<$@L �uQd��)�w ��mӞq�pl9ƥu������T�;���-A{�*�*���2�,��c�G���+p��i3뎚�<��͜�HW��)X�}&w���V�5�{�%py�[�t\�U@�P�:z�H�� ?`�0����#-��t�o=ɔ����C�ַ:�_/�D�4�d�?�Mxn����3��4�&Cڝ�n�8�e5:��C�Z��]L�lhF�1��=X���9[�����t4�X�%0V����G�=U���E�"?�'}k̈́#=nԐm-oG
a~��T2�.bϟ$���}��_GY�F4��`]�}��^��1�,�$�����7�#���|e11�A(Р��y�R��Z�7�KK�-zr�؟��l��bk��o��b̹܋7+uP���yjv�-O���IFAo���G��f/�Gk�3���\'�e�ۣ��A�T'`�h�6�����i,5�JV����`�uA�(����&��a��ھ��F����Z�4
"�+ߝ]�sl� G!?'��^�����-nm��Rq��qKv藫�;�2������EϹܤeUw��]���^y��߱�7�o�yb�b�g撑�0�1J�+�A�|x72evt���8[��)�����a��Mި��iH 4�\��p�z�����"4E���m�Q�p��0u����rs��ե6�K?m%|����\��㾋��,�Bx����/X*BZ�p"?ɄEx����;��24��#�TD�&�ɝ��ո^����D���/B���Fo�#U9����.c��/5uƭR&.�A��W_~Ƌ�X�(UԈoE�����$>(����	�C��c��X��//y,����^�xL�S3{����6��wy����,�9!5�?$�|��k�;�lԓ���3����)c[�øǡ����s+5C7zq�Y��
�nZ�3��E��j����P/;���%��� Zo��DYd�����R��UV^w��&����n����+{E������|is0����!��q>d
��ɔ�>	�v_�j�{j�cB�E2����Y'F��/��+�+뽀��X1ۀ�>h��u+�Q�Nk"��N�0I�@���s:��>�T��y�3i�3'�
?�q6��qG�Ɨ�=A�.bH�T1]��{�471U��v��#�5��LG}g�oNMX�0&7��y��8��D/�< $���TGt���t�q}i������շ~ �n%��3Y���lNs�x��6U��|#9���Ύm�u��v%����GAW��G9B���V��0Z�7��(�o꽅�$�O�	� �f,�;�Ic�����p#8+
V0xy�6��g-�_L d�1��� ����ߟ�?r�6��:>q� �w����5r$k�CH��"���f'�h�î gC��|ʢ(�3�>�]]PLˊ2p"�w�}1�����X?�����\~7
�DK���"�K��tm�5N��6"(����j�u�Y�n��KI<�6Fl��&�}'"pB��!�P�;G��o�RR�����v!�G0.Z��s�6=Y�H4�gjk2ט��=4�5�B��+��ys�vs����z&%��:�X.�q�3U[{�s=[n"���|vS?�'��\���>�%P����ȭ��J���)��� )�R�C+P�<	�tĔ	��zWZǍJ#����1τRW!ީ%���'�=�eZ*��'�Ԓ u��,p}�4y|�@耸�����Q�}�%��vK��pOoo�gD�d��x��#ښ�[0��1졺�V�-�Z�����v���h���~��t�����7��S���C:5q2�z� ���_5f���� �b�NUrL�vמ^->`@��=��Ɵ��v��/?z�魡iZ�}�,i�����S��+W§CoT�����܍�@'���Z��5�oZV� �{uBUS�oa��[�V�G�B���Y���߶�8�?��9�p<�֑�]Эl�q����Ĺ�@��2����{��N��MZc�j|�a
��x��/�rv~mhٳ:&�q(��-a4�������w�!�����v���杨V��*)ZF�2H��%����-��vVՊ<b�ds"z��Uk揲:r��|S�4�6Q�l�J{��[�顨=�%��|��<U�3�Z����VWU����f���I��|-�զ�	1n��c��$��b<������O��-�~m+���w���6������g@?~�s-���E~ͣ!r�����7t��7Kt��R�o�Y��i�\ͧ���������5'������!�ut��Z�(���P�1[�ۂ.!�Bsf(gYg���`��,"/D��)S�nx��ͲxP�w`qG��0H%Y"�<,e��T����iw���J�f��`5�(a��M	�h:wJK�8�z:2�?v�������N!�h�s~��Z��^Qix<1~�)�V������(j4��� �?��Fe�c@���{�M��w�f�����4��l_+e�Ů��5wZ�w(�RW���SyЗ�f�X�f��[� B���7-a�Jj�TDo*-=���/]]$Q\�-^xX�2sYÁ�IC���@+ມ󭛤ڍ�K��C/�@���X�y���!EkC5��J�����v��"e�����)S����&�'���Q��78�·�~h���>	;�*{�&+����5���4�A�B�C(=C����z��ؒf�-W�GOaq$WN��R�"�_Po��f%��i�i12Ia^�i�	��3��ϓx������[UG�Mm�Da9�)�z5�D��&�g���A4��N-�nw�`��T3��o�����n
j 9�>��9\�d'��&,鎇s�?ֲ��x.D������䌐�
�A+��(��X$z#� �/ o�F�b�T�?��?�)���.m��u���,S���Ik�����W�b�F��D(X�:\��p@C�� �L<F�;�GW߸�e����x�.� !F�k|�s-�p�s��q�q�k"{�ˈV�L%Wn.D��׷�����h�Z^ 7�c�j�xl�؜�4�K.<�*R�56�i>E�kW��@2��r�Ô�,�k�n �;�Bkp�۷j(45�*/�����' B�(&��G�#���JR��G���v�z���$����
4�I����s�=Q9~ 0�I:k�7U�?|y�')W���:N������B�IJo��|�@2�*<9���lQ�)D�l�V������EK��C�ޒ͑d�um�Dh���w׳�_]�q��_~G��u�.����7�����?g��e�~�r�P���S����?�O��<�O�$�����e�@��C��l���`CV�'n's�r��7�Z��M>�'�|�K���n��-�����^ �ph���3���ny����Db��K7'p���$۽�8�u��I6N�i�2�I�܊P�o�;���<#��yk�.�r�>d��q����{H�م�n�9�i�Z�&���AT���9�����GL��R|,��-kX7�B�׾I0�NC����%�����0�!�V1���N-������������ ��V�T�������l:.d_JʣY�S����I~��=��1`8������������<��q?�*��C�x��^Z��8��3��D��q%���%�
n��nf��k�E.�6����v`S�I�/���1��q½*�̤Oj�fP<Ik��}��M�4�׸A{B�A��Y�pD<����Z�ܘ�Nh���]��c��L&X(G5%�d�����}��:�����}]�߈r�8��Ȗ� Ҟ""Zn�)�>����Z(�GZ�Md+Zlz�O��%a�7��YD�K�_r�n��ȝ�(V�U@-���3�h
�X2��e����V��ާ.��<�|��:��H:��u��p�� ��a�"��fL~��Fxa�k8�34t��u�r�7�%��`ƃ}�<�o0�~��s��Rm�ః9�6Ed�m���h*��3��N��m��MM,)W_��`�����.7gWn��Ȫ�Էdk��~���
��:��l~�xE��{A��� �Qل
��;��jkr����"3�5��*kB�*�[ Í�,|��N�J�ֹ�oS�_x���A� h@0|�|z��޽|����J����u�}��#h����_��h�$��Z��(���?���P���Ƙ��9Le(s���'^Kf|&����^����"Б=�w���a=��3�ke�2��Ģ&p���ӟA��F�N�tZ� �S5pF?�����
���V����þ�b�Õ���H2h�K�:F&Ij�y��ӭN����@��#,J��m��o����yj�|}N��/Oh�va�0hd;�[6(���$�����f�J�	���F����`�����Z�X	(���qsͥ��.eˤ堖�a�ʟ�sD{q��P
�2�0b-I�?�?}G��p��v�s�͵}S�L��	��@-�~v�n��A�],nR�u]��S `
ѶNY�Ps<>�8G�'�{q��[��4��m���H�R�5F>t�����������\g�o��4@K��ze�-��w[��M�PG.��u���!q�m�X�I�����+8�k�{��Cw�ak��0v��'Ds,H� �/�)�K����IB�8�\JJB�ܸ��uk�3#=�{����+�,�/�j�n���9�>�\-Q�� E�������
�|�\&�7�E;jU�ٖ+yU%����_��RQ���P��󡛌S��ծP��u�-t���U� U�6�\$�2'���;������ű�6ODۉ)���4L\�Ӽ1���Y<;����
.���Ncq�gT��1�{+֮�qxO����=TB8� �K�Z�<"��p,�Lv"��N����o �Tj!l?)p$���e�e����d����o���EQ���y�ӝf;�+q�BI�h,!q���w&kW�ށ'G�G����윸B��9�֍Ky��N�T��f\zf|�`z�_n@l�5G2��K��5XE���� @f�?F�Z�[lb~�.!F�z���^��GJ&�氦�i���S�"��2�w�NƘ�t轐�df?ܑ��Ω���\W�W���Z�;t��� �\c*���<�`n�^���G���	5�n���5����݌�q�P�h�qH9a��0����&�P��4�؄�L��v�#�`���|�e��������&un�k˒PJ ��3���ys+��U��<}G\���Q>�Sn~���f�F{U�^�m8���쏆N�{"����V��^�lR��"�("�Q*h"�q_�"��H���O*u�]���MM� J��\��� p\o��'�׼�5���)���O���|�U�;��	xP�7)d(w���&I�Ș-F����6�U��8x��'� rMe[������uE7���"Z������=�9m�#�v~�ѢUO�#�3���K���>�Cq����Us�w�>��SF�q�0�m[Uq�f1�qnb�r�r�G�770[�tW[��}%���릤��V�")���ȭٽA�����k�"B����j
zUj�WY>�&K>�4F��8$?w�f-v�ՄS�<�;L�Vyo�)�aA�,9�ϔc�Om�����s��`�L�Vl.(�;����Vn��g�s ��d�-�'7GP�+�1S!����kZ�`/&�-�Ƙ0R;���y�u;B����V�2���!�6�a_�%U����`�p������$Ֆ�!��;�KB$�p���w��F%�܆}�Y�9)�\Լ���磔�m�S�cx��߹�C�[�(���K�$/��`��W�f�la�b�S��m� ��խ\�e��+��޳�&�ѽH�&!�&�����1NY�?��E���*2b�O���|g�^�7���Q�`u_a`=����E�vs~(��h'dB�ͤx��@�n2Aph��񇩗$g�Cs�L��^��l�kދ����3��֨���g%ݷ�:fMt��E�.�d��k�=��;W� ���͞�,N���_��d�O�?ɩ����ؽ��4A������4°�*rސ���Up vvH�J��l&�c~T �y�+yp�Iva4�N��gǫlZ���� ��K��e�O�⥗�l���S�ފ�LָE9b���v�k�#�(��A9ϓ}3�=�xrݯ�A�����ο?�^`���H]sBRȾp��fn��ʫ �$ԍ�z��|���đ�.1ݘ�~-T�Y�K�m@�L�i!���{��?L��/e m��Ӂ������'�vؗ{�a�~�|m�3%��k.�(,-����x�$�L����]�p&~��VrXhd�!���(2awJ��4�Uzp��D����8<w!m�wm ��g��eO�ޑ	+�M��1u���j;���ޠ^,�⽸;�B�g��?h��`���Z�U \�q����Z�dn �u����ʯ��*�����.t�é}I�T!��e^�3���N��3� Wh[^�*�Gj��GPI����}��[x�]J�(5p���(~�6�M�o-BP����<����>���	��:��g1�S#px�?�	~c��!��} g�C~'�����5!F�5�H��>w�������.N$����Df�J��2�X!.�Z�O�ep�v������
��X/���my&��nkq_��e��n/�	cċ�S1�!4�d��G!�d,'[�"UP�S��,V�U>�0.�hR��&ni�DҊD�yN-�1�3��R�#�Ԥ)����9�R�u3� 	����kf&����=�g
�0|+�b��P�v3
ᕶ�pM7cH杀�#����H�E�1wpK�}$]�l��o�ԉ���'н������%UN���|���
��
�F���*c��&8P\iw\�֡��..b��3�bś�{�²6ۆ��5D�ýqRŭ�J��b��r��?��م�,��;J��"}Ejӻ ӆ��y�2�n��!2'�{v��䕳�v�T������"{��oW�9�Bn�60�g��;��N�Vwj!����c��f]G�I.�=�����7�t���r��_2�� ��i��+�$�r@�ok�uJ�S���`d�C�_�C?��ܥ<�C<���HxP;�L�J�3;kaW61��Sj�_@��h$GM6�z�zI������+���(,��M�]}[��˨����t��݌�C��f�H���Wq���$$�&[C$� [�}�u