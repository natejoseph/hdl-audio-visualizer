��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���֪F���[2D���DU���|��'"�2-S�T/��tp����8���5�V�:�ǝ.A�%x�%��R݈�,P�L��ԕ;oJ9�����B'?@�S����U�����[3G��+ӣ��C�>�XWx����/u�����4����^�#�E���}�]%�:p�Hy�����W�F��2:�\��D͒�����8�v&ia�7s�g�ג����#�Zs���c���/�a��v84��1�krl>�q�)��zY����}�|��˫-xI&�����iC��q��M�*w*��QM�{��כy���"�+���� ���8�TD>0�tDDUFN�sYK	�M���ь|ơ/:��M=�^��{����?���V#pi�^aڂ�0����52����q�@T�]��_�����J��ʠ���0�v�;i9Y���%�L(�@�Ap^�U��ik�L���{�}J��$�,�����3�}�U�L&A��'�^=���ŦR��[2k	r��Z��W�����ꊊ|O��kd�L5J�ϘVE�Z&�{��U�����C�ϼ���˝���퀛)�ߐ�[]�����M=B��5յly��£t�>��!	��Xi,;��~��vћ_��7�M�gʇ�f#R��k��2qBf[R��{
���NI2_� �ee�w�	B&�&}�'��l;�tǉ�br=#�5Au=[�Ч�g$@���_��k�h\��	&��a�7$��^@e��|ƨ�l6"���6V ��q��K� 9m���=+vм$�wJ+kԽ(�!!'�r4��ӟ^�t���=�e:��[8gI��ˇڄ���g�x\U���%2�J+��W+�d�J_�yˠ���"�q��'��;pn�R4��x�o`�s)z�$����}��6|,�y��P�Ļ�Y�zU	hO�T{�+TUǂ}�<�ff[[����''�O��q߾6�%<��..�~0�̠��+�ӇlN!�$�h����{-����%��{�R1�>8�B�m��1�s��}�废��"v��C�0U(��M!�N��V�b(�w|�k�o�a���ɹ�GW��v���r���g̔���*�R�. dl�1/��U�72��P/8u��& 14a���$t]ڛ�zF�4o�<���WE�r��I��^�5h��GLo~;'%`��:׳H\����Xf��G�¨�νtBm�	��Q�M��C�\T�l�$w�mD����k����2g;�i�~|��Sb�L�/�NB�h8ܻ���>ꈢ��u*�nR�q5����<i?�4b��EU���?Ux0�:���O�4$���\mf̜�:��5$�%��h^��qV]F�f[��G�ݚ�"��=kP�`�\�l��1���$Agұ��=4��5���	�Ƈs:d�4@���챝��q�;�^n�~�婑�W�}<ym�,�������1y�_f�;���� D,�(�o��B!�x�B񫪠uX��R#a��գz&j�+����"-���δk{���0�@��P�s얶E|�x姼�R	Yk�w+��=�Z"}�a�?�$��2��W+� �� �C?��v�m_։��!�0J�bF�g�\�tJJ��.tدa��ᫌg#�� p�m"�W���u�ʎ��hH%US�z]�@<�L���&7ȝ�2���<Ap,�bʾO�\�D�7��E>��[��'�����MSJ����?@�(�^�x�{�4w�H��F�*�iB5�s�]�LT���E@s��d"R���~�}e%v��5���Ȍ}��!�v�d��w�g��tEt@�e$G���D^?�	^(�j����^ֲ�Z�:��˗4���K\|�.]?+���,�2�[y���h((��噂VKUy�)ً�jiH��!d.��fM"� �9Ȝ>�AN>�R���������.�)�l��ڸ�9,�I��V�%MTҩ�݉�ϺW���D��2@n���";Zƙ���;ߘ{%�߆���o�
s�P�.u�h/"�ł��������c?�񍩹�ρ	t���=2����9�LT�
�IႦv��.�k��M���g�ٻ693B11���v���֖�omW`��[.�{�nKŕhQ�m�D��fG��x4�y�l�'��:H���,ɮ����ݩAsT����!s�-�Q�uT��=B-�.�X�#ј���
B��J�P'{�^���-&y���"�qt_(�j�h�qʃx�X´�4�]B/�ZX��c���5{��I��k���������3�	$���T��	��?�H�����M~s��
�ެF5Y��d�IV ڪ�-������o�7�}���J����f�{����)�hu�W5Yo}��=���S�xU >�r^�=��@�u%�q��)�fA��W#���opE�2�)i�^��+30���ѹ>
�D�H�uPەz\_��96�^n4gLl^��놫��|������[�Ri��+��(�jӉ��h���-��^�M�;��sSu~�qں{ULH�F����o>L��:\�2
��^9G�$��
����;�ǲ��,�E�x	��B�S�Pnv�t�D˻�W��	��/\��h�yK-��]8����7����<YE�z�3�Ε�����P�(�D����{y��nN7,���t)����NvgIK_?�B(�B��g��l=�Ω��a�i�0�3xT�8
��]�l������~�`w2�A�F� 唝��dPP\�S�ڹv�e(U*sw����-�YE��/�2�� 
J�J����%�$ā�F���Y������JnlO����?�?l� ǅ�S�ڈ��N"p�Ud1�YK����La3Dc��X.�4I�@�+z) CT�jzg���'��J�Q���&݉�P�Bd�����mU�t�1Ԋ�l��"wj;2!�b�K�#|�j�jĦ7R'���n��Jl�-X���dɌ��z���<�����4`k�K�	���ߠ�܎�T����X�<���r�ͅ��򔨑+�:_���KZ����ࢣG��>�i��ނ��f���)Kf���aߋ/�OO!ҡ��h�P_EJ�5cg�0�ɚ(eK};���LO��&��9?O��L=_["�D�I^V܀z������PC&�~�E�Hx^�cM���u�-���Ub�K��)�*�k?�9)������8��T��@�8B���|�F{��'�/��1�Q��m,v���MyڕG�]�g��s�2,rTߗ�;����-y%�q�� �6���Vw�֨����"W\��l�T�e�j���+c�گ�g��|@>��єG�q�����4f)�c�����`��o':��%���N�r�	�n���Xa�X�RMg�u�'�W�����K���M��!L�CK��}���e�ſ"�!�j*gi�wX(f<�_���(f���`�UM_CF�5^X�Tv�؄R\�r`���!R�U��mn��z2Չ�5�u=m<��6��j�J�)�=�j���
m��s��Z�<}U_�^	��wG�k&&�y�>�d��+�(ҐCl In��\���e�κ�����͈�+�o�e��A�Y@7{���ف��:�b[�n��lfKT&]��G��\�k%b6�J�8�$f^�}t5��)�՚W&`��&ɨ[�9{q@NgQrLߠ^B�5��W��on�����6�BQ�Q��b<"��|�un��e�����c=϶C�݌i����/fGR<�L���qo�}�������h%-��]�K$4�Ƕ%Zr.����[�������##|�b= %Z_���\􄶃r���O��s��&`�I��
R[��c��s؅`̗���*p��RX�~�-��'Z���ha~��C�d��LX�Ҋ�_�]�ň���W/M�r������7���>���G�0,�k�L%�|�Pw���$��S}�U&2���f����6�r:7wV��ڪ�?Ki��i]���f<🇆�������!���k(��u��yx��R�yD�<��F}�To,"���N �k��m"{[.��ݔ��y؍��̛�!�4�w��YB�s���n��n�'/�G0x��V)�B\���-m<2�P�9U�T�:���R/�gs::ᔍґ��<���>�����_��X��~Q�5^<�7]ұp�w���.��𤹣�!�����\߆��������������ގ�N�8��ͱ��# m�{l�6�A����,�i5��]� V���{����<���O��m�uFT���[ݍկ(d���\�R�J��i�:|Z��#¸iE�B�1�ON��J�[��Ti�����L?��@4�H��?%��f��� NԬ�Ƅ�M�|~�uk$T�w�������Z���8���p�V6�3j4�?�/��>)!
����)+�Y
�8Q�
K��UF�|ާ;@�$a+����kYa��Hżb�v7#313Q�Lz��IIk�%"� ���3ƀ��,m]��Th����_I�!���|�O�	�Zd�V�+�o��t	�c�p���fc�18�@?W��=p�Zrx�az�.��,�R��vM:�]I�K��5,j2���-8��$d�Hl�Q�
b��ڒ{ɡ��^1CTA���F�_�gJu�x.4Rɯ*9��q��v�vUH}o��:KU����N�Զ|r�_ڈ�=��~��I�P3��&��Ȱk��� ��l�-�����ڽ��n�ْ��2l�.dV���Um�Z�)�_��/�����Z��|-Y����f}��jh�o�e�&3pq�e75̱�̗�p��?SB�Ɇ���G#x�&Pr�p�޺<8<o*��=!�x� 2�tTE�-w�Xs��t�K-�  ��)Z����F	�P��li���eC��N�Q��Q){,Dw0���麬�^/��!q����(iK���%W�+&�jD![M�=��\=3EU�CG2���Y�e)���J�n��#G��;0B۪M�l\��>��N�d���h!g�k�<o ��������	څ�tԷp#���2��J?��&�c��^����K����̳[)<Go4��ďm�.�PC���]�Q#m�lH�Q�Y�����5�b�{�c�Æ���zԠ�B5Lר�����ow�Yb��ftL���׷^�	ݜv�e�W�=�ϱ�����b���;ι�;�yM�⯱g�g\��������U�-�]8V�#���1�TlB���݇��q7�qFz;��E@�f̐cK��L�2�dؙUke���Y������a��`�	s��d���]�`_�z&��v��LF/q��3���K)��p�|�a���3���C)���k���P��5љ�ax��%�#�CV�JrjwvsƗL0����V�Y7����Յ+
C�>�7q'���\W6��Ȝ� ��j>E��.mY��lӂ���2^�=�U���\�8ە�����F��'E�ml�����ὖh���8]��Ic�.�1k����������Y�f�F��� �_�N�h�z\��z�n�`���eА0�_�Q�	��L��o��9�� �u�����A���z����� �]���ZEn�N��Z�|ĵ�yyh��C��M��&��J{��z,k��i����"��h�D@{*6��P�3��DKS8Z����y�M�3�z�n��K-��r��łf`��R�b�A�
O�{����h��4hF�:O�a���%z��>�L2���?�޸<X2*䅻�����ٮ����%�] 3�������D�94A�Bˡ������R����gR;E&����u��`2�OX��K.�}�	E_��g��r��A[d�&�օ���馟������n�3����F�!�G�|�rR�o��G���_��d��SO�$��њ��aO��������ʁF�ӳ<m$�$�ё3R��������@�(*(i���k��Ns�b�2��T��w뗰����C6Ҁ���"敂X��%R�Z���QW ҭ��6�ê��v|��"�r��l�r�BkX������ӳ���u
9�SX3��TN�&��k����|y:���u��w��T�S9/:g��\���bµ\EJ�J���8�fOَ�˰�I���mHv	���ߏ���Ԏt�㼼g�
g�1y����<�	���n��ڻ��f�Z���_�Ln��Ѐ?����;��?w�Da�e n<��uk�M3D�l6Sqx��N�Jk��|�6֊����;��2�G�|�4*I:��W��Z��Q�FW��7�k�0A��[�
w&�����=a-��^L�15/�Բ�ƺ�_+򍌪����ְ@�<���]ÌڧJ�fټBX+���n�ZߤZ��=M�������b�N���[H��/{J#40� h�j!�_1�r�2�=����5�� �_�A��3�ǅ	ᴌL�F�����]K+,+7�Z���E��,'��(�H���Q��^A���.x^-kVΡf�.��^�I���18�l�OG�߅�%�[;�~2ԉ�?X�t�8��Kߋ�LK��?���7<�������.?2k����?��׊��ߝ'z�@n��ߪ�먞!�P���z�Y��<��S2]ܪ��'�ݔgP��#��P�"�:�s�K%��b5 4�P�gN:��LJ�b(x�Ү��KCݞ�!`z���T�0`j�I��޼,|�N��'?&�98���舘x[7�xM�p�»Ql��8�# �����9�)�ql�S��g~Y^vƓ��j���W�� F��]pۊe���)��Zg#�a����(����(�˗�=;/F��h"���'t�@�0�Su?9�׹��u�]?mif�?W,�9Bj͛?��|(&�=l�NUR
���C}�A�DU3�۟�@� �d�b���ҭ�tzA'��!,�"�,+��Bo�M���4�z��M6���Ov5l'�d/BJm� ?Č30�B����:dd=f�O&��	b.�5�j:�N�QF���m���f�r��x ����� r{�I}.�Ψ����F���RGo�?\�����Q���V!�?�;���D����v x��S�n��mQu���9����_�e3�ȀW�9ݪ!ϥL7��N���S�I5�e���.s�|M}lex{�F��N��+�b[rp�l��I�� cI~�x�#���o��8�R��AM]�7��F�wz��EI��ݙ�Ol>P5O��� �-k'�o�=h��o�
76�hl�IQ�F�z�e�T��(��.[�~�cD��� )�F��
�=�M9���K�?�������*wW�)׸�>em�k���d� _p�l"4��SVj���7�f��M*s��O�K��a3�:7��'�^?W�g�z��U_�vG=w���i�6���j\8^Uj�T���AlT��^�"��';��ɨ�_��v����l�,�	�Í�Z�cL��:s�ʇ�Ec�����7�E���YI�<X�NlvjH��5���>%��Fw�'X��m���!,�~��(%�Y��^ �����'*����ın��K��1v$]���p��Q�^[��C� n���q5��������v��G1\�+s|䈜�(��تC���W!��tmc�A�±r�8P�g��W\N�9+GH�e��؀�Q���J>�4]y�-k��߹G�:!"�^ꝸ:��X�<:Mw�S��L���|x@Ys7?��:�b�}s�CVX�n�26�1���%}�"���+I�M}��`���B��ۏBZF��49���
�w��a�hT��]�̢�Gg1Z
�	��ZF�P�J�b�w�!}�
:>�5y��ɢ���D��Fu�}�Ե�mK���Q�G�_�o��4W�<�w�}��/��\6HJN=��7(�S~���=+Kh�����DY��{'>K�̑21�dd�pv6�fY� &�B����`��D���
v��x�,~����30�%�*��������	�5�?c!�� ���Y��?�8F�cN,�ȁWn.��;c\p�à�-�o�)��cr����8c��3�W(�:�`�Vg�� uuq�E.�~��C� ��Mi��{�	�h� ~�l�=��*\6|�6(N�z��J�XJ�����@����!6�g��Q�� ?�9mk"���hK�u��z�f�R~�j�-ڼ��s}b� �]7�������Fa׭'������BEm��_}��z���X3�B�d��&������:�I.����_����]W=!����W�
h1��|�w~̓b�k��?�q 〣W�F�kj|̰�z� Y�\�5�}D�� �^$��:�e��.e���0�W�?=��I��0@re"����Z���6֝g4&DX�΋Dn��g�C�Y��QߨSl����9F�V����A �ٺM�c��C��:��a����6:p13nU̝=��y��ɔ���<�5���z��9�)�)�� �3P>^Xa;5Rt�#���f��V�{��y�Őt|�7��e��]�t�5��b<����l�-�h���8Z� ��9
fo/�������(Z-�.���>V�z�+�����B��,hy� �XQ��A�V`1��j��.��hGe�%U}�(s}�c�,���nz�@s�z��`���V<y������C��� ,`�k�Z�&))}���\^l�������4�=�Ɉ�P~�爝$+0�AÈ�*��|��f��ۂ�it��ƦJ��)C�߈�9U; �آ;@������� qA6�����m���B�j� ���}��Uf¶��v�xr73��&cc���,>�6͓̓�l�۪�/�.�/�qS`�1B�����0*Z�iJ�}V�+ѻi.�3a�W��%�-�͇�R��2�JJ��Yھ�_����g�!�[�V������K͞�;�p��== �A���u #��=V�����M2k�a���J�c (�UǵE�Q�Yv;!%�O^Xg�9e��u��˹:��I��؈X~��������e2w;��
>�>��5����趩/v&I�G3:&&�E,��za��;R�\�����������|cY���F���uI�����\��ax�ޖF�}���Y��v��y'�0��O�p����@���נ�������@�zG������bu!c�nfh��/���H��u�R�I�N�Ֆ�0��� �+ʥ���_'Q�p=l�����N6�e���.�?�S��r/lIR��Y[�b^��Y
U�����C��>Vj�PM�9Bd\b��#���X���D�[�$�=Vd;xlm�Jx��&�zE��R^$���U|�4�`�H�X�'�w�_-��BnG`��j0�j}��04TMz��W�����XVG����]��eF�ԃ����]���X��r�]io�>ף+	�v�2ǳ�QU��y�"�����,,.��w:�r��O
)"Ո����xJ�ƹMD�C�N��ؕ�B���ڟ�B�?�"&b*��;^��Q�&�c�� ��hssgVG�Bx"^0�����r�ط]��vGC5���Sb�dNw3Yq50Y���m.�<j���\f�
���w���W��u�*�h聜5ӝC�K���6�g�n=*}QĀ>�!ϛ�\���n'?V�0�7��� ��w����8�44��n�`��&w� �;���^����׆�Ė(�`g��e/���i)�w�:�L+WFΚ�B�G¸�>Iy�Z�Wƭ>�! ����Ip��_Bn/hT��� B�.O4�-գ�}�׹(�Fi�y����*m R\�h�&��iR�a���a��_�'�B��[{�W�ӂ������u����׶Y�Q��U��@t!�0B��m����
>A��vU��J�9�`+�}R�ʟ�[@�^X�p��+�{<�P�'�=|�#q�%!٨����,p&#a�B#��g�i��!�a��2�ug��rƊ{W�L~r��?�Y��c8b�hf=�xöu�S�"m�I�ڒ��d4�_˳E9Fg����
��6�� bi��8iQ�����}̈́�tZ�~�@���%�`�
���йp�*�C�̜y���@%%�EG1�?�zo���t�Z!O��J����Ǳ����� �o�����&��Wn��R�ǫ���Q�FJ�o=zN�#���Ca�,���^*�S�k��Q��v[��Z*;d��Z <�7�a��ڑ��"#�?�FY�|�x��5ޮX�r�E��U�u�@Cݕ�y�Œ��'m�B+dJH5�T��7)����n
��,����X��mшOd}���`�_�Gf�X���P[�y�=EG�M�ڷ����ۤ8��g�sg|��R�@�w�	�����U�0i�0��'�m����I���L_��<5���l �?��D�w��s.lU�����}��d�-`�.G��C�h\!w`�XJOH���b_�g��I~�.{X�@�������
���[���#���EOt�~f^l5&�X�L�bm��1O�E?������p��^�[��K�p���,P��`�~����D�\䄺h?ѐX��1
��#��D}\��
��;�����:�����(-�\tϞ���X($�E"����\
�"9¯����^��J��u��Z���w��(J��q*eсH-xU/���k�� ��6���{{ί�H�4�g�#�JX|t��-�
:�#��6�^���a�L�������p�r�fR�*C��~e �$k�J��r��d��β��{F�ֶyC����,�H��w^��H]��A�۰g`ʿ�H�9�����+j����3E��"��ß"��&���tX�X��L��][�}2�_<��MV£�`i�
�3D=���
����̯�:�^M��~'�0���/����9�`��KΆ4�JޕK7'�<;Рm�αX���Y)�c��?�#�V�gqtx�H,*�i�7\U�#�n�At0c3Ikd5V�U�Ϯ����N���g}��{��P&�G��XC���� �d�z�P����Hp�WTJK��'�(F�(ZixͿ���ɉ��Pm0��^d���v�`A���i�B��IUe�QÖ́�t��G�y�����BV�۔�y�v�K��@������=m҈���.��z�*Q&ڡtj�O7�'dƂ�}�J�OC��|bxs��D�op>�T4* �����4��"B�E]B$Õ��(�g6�˾���E¾��#;��b�Y�
�t�qY	O5'�PF_P�0	�S¶ϕ�9�빹�Ps���Q��@L����/����2.�{��&������GG����e6E�͡�	OW�xY��]f7�
�����������*�ݱ=9�k�����J����F>�٫Q2);cd��}tĳWqh�Ѳ�#&yT*$nta��ٴ�$����*4��ʏ�T&Ӗʳ$��m��%5Q�h���rw5�<��>N�� jJ����*4B%��	TWp�ECUL��y��^Iv)���pe��A`�3e&s�&��'!e��u:�V�$�&������w�J�����?e�g�IJ�>,��uԞ>3���qqё�@��j�u��hF�QߩL�T�?P��?���W��۫W��ؖ���}6f���Le+D�cF2�l�T]4A� 2�_S5�@>�8%��քRϥ��$�hZ� ��ر�[;&,+�e�q�Ҽ'�	S�sN�z1�$�c��Q��ҭp���78��}u���x��v[��8&��g6����v�L���ρ~�Қ��Y3��=�!�ȹ,
�s�-39�(�2�0;�X�7V��G��o$���ϲ?�"��H�Q	���2��B_=DQB(������Ș����e����;��zT�\��wwv�"��C��7(� q�I��:w>���o���6oT>vN��3}�ѥ�>d�i����q���Z��Ƿ�w�|Fɹogr�16��V����$$<�_�ץ53"��z��m9�N�z��:��ZK��&^���A��I�+�������@�X���x�6���(!�JՋ��w�V@*]�nE�F��寽���І��R�����.���*�ϋ����T��$X0۱��4�2&,ᆒR����4ag�.��1�>����U�sKQ)�G/ C#l�X���g��	�f����<i�{�kx]w0�ziG-c-�od�Kzm{�;WUC�Q-�D�3L�XU����1�Q6e��j#qc����3��Td��7|��5��űY�wc�ޗ�����k�z�cE7]�*�w��P1�+��%�g0�K�pI��@�����C���X=���U��J�V��x��ϕ�K3�5ݹbY`��4z�m~���N�(-x��uc/���ѱ��������l;�UR�>��g�"�
T�"
X�G�#h<WB�MF��#S�0��鿂(S~�i@һ7spλՏ%p�����w�t.�u�z�1d-P�}7�p1�[�f��_��g�/�R�Q��:��`X.�������
 `��z��,��c<�T2��v/|����>���*V��Z�
'|#�$0�
��U��Ir0��* v6����?@�����[��
��
ͻa�	�P�Dd_�A��"n�sB&�V���aגgO����4��-@�$w
7�nG���
�Dȳ��*��rT ����h6�0�R��aϿ�_;_�E����rv��@���mِ4��=�Vl��TC4�/���g{��P?���{�Y����k`�3ɒ�}@�i{��ӈj&�q��j�8��~�W�Yi��t��m�zp�NN�L =沮92��+	F7�����'uv��k܅�r�.(�ssc/���2~���is�X�W�HƐ;�B�0ʯ��2�FeIh�����]��+����p�.F��>�@���-H4��5��W��u>�Y��W`W�h�#�V�l|�����SH���7�?h;&��kuBC[dvq��~��|ܜ�X"Bn�����#��@��B!��"�я��9�hL�����bX7a�%��U�:ٟ[Q��j@q�PeBT"��t������[����=⨠êx�Nc**�/��
��h�y�Ă�H���B�-�#`n3�g���(c�4j<��y�_�l)�tʨ4���!������(j��m�� -;�%H'!�c��yd}�թ56���,�>]Ԓ�펢z�1�6|>��j��H�0�,��?j�:dT��AP�=Ѩ��Q���pØɯ�@�{pj]Sl���ބF3g�!+3�d�nɬ ������-s�r!�3] �u��ԫ'�8�粵�{:kaC^���;^�o �ί���p{P�ׇ:Ѵ����Ty�G$�W�.Ik�;о~������wz ���Q(���/a���K��b��Ch���PՆ�.D�h�,�|�1�k����&a���V�q$���ʗ;1�H���I݊~�����=�(-��!9�������`��ޟ�lB����Xs^+H/�o�qU��+ ����姅�ؚ���E(���庉b�g������#e�^;72�P�w���\"g�W�����u���B�HX�ׅ�̋�}����r��,�^|/ȍ��q�{ܲ���x������L{�� B�J�h��39�c-h����s�l,�1^��eލ_akY}]�DF�%��1�j�aOE�n*��2H��ݮ1԰�n�-���͈��;���=_\z0Y����'t�Q��ڔ�u�Y�ŵ�:v=��������2e�a*�:u��6C���l��#\�xC��^)ԸQ�;M���ϱ��.�Ǝt�0�X$M}�y���7-H XK_��1��Y����]'��a�	����jr���p�8��b5V�<�4=$�Rk3qJ�]2�,����K5�V/u�u��B��x�-�����B�-�ݼ ו:�?��\�'��j�X��pgmآa�������|�s���	7�(�0�w�/��>�ݔ�D�d���+/R���׍W-����K!vƚ�;�V�A,ͬ�n\�5:��l$���v�-(ygy��p����Jm���8A/C�	<䎹O^s�{*E0�=$���	\N��_�y�WbLyb�)3숄eXDܤɉO��j5a~�q������I��>��Tu�¡o���/$�Wⴘ�p�r�ۓ�*��W�.�R��2}__���Q����
�)�PL��\�/{T�E T�LYz{�1J��&��x�y@�� ���t�4���@O�i5ݜ�@���l�x�� v��A.
��ljȬ2�f���?a�N_n����ζ�7�DֱȐ3�80S8u��L"5�?�i�?�H��0�M$z�t�x�(v��;�����/��� K�\��\9��c��1-��.):·�G�HuP���f��|��5�G��ɫ	
j�Q�J�����X�KeW:�h���P��)�wꚑ	fj���rPV#�?ul�0�eq�����*
�1�ƢC��V��eysISSʜ��2.�q,��zq�9�t��m�A�ޒKf;��?�v4 ����������Hk�#^��2�!�H�������c������rQ2��6f݃�M,�&�1 "�;yu2"լx�
b~��'�� �9��&����������w���#4�J���b �=F�~��=�\.	V/��.�8׈⤋����Mg�� F����ZƘm��VR�^O32{fF�i�Rz<�����1�`�ሡ�l�A#*�� J�����r��/�1��CWG[�g���nr�sW�UV<�,]���a��S�ֿO|M�NSo?��ҳ)>��'�4��󩻶��%�b�Id�.�/5������*��ou'Ƅ��l�!
Vu���r���u�]�/�%�7/DH��'�֣Es�v����.�9$a����T$a�E�z��2���y~�Yv�b�O-*O�Y"��<'�� L	f,9�Q�2�ctT�.��"�k�dZ<n�^vU�a�l��e�
�
�=1���Z)Ȝ�X�(�Z���h]���swQ�؛ڎ��ah3�mxt�f���C���#b�/�^�����6�бȪ
����8��;ry�Y�w�Z�B8�%c�g�M�1�8ȷ���a�~J9�{�i���f��$��;U�j�'r*d&�['��.��6�O�R00��R�Żmy`���I�+���|�',�7ѫ�B�Ӯ=AW��;q��F�G��-�,�2D��2�R3���S��a+ױ/�x�a��E1Գ����=���J!U�i���J��X�U5k7�;(P�΍�O��z%���e��5a[sl���rsd
;F;+8^~]�i!ZM>9mM\�x��q��t��i�ˌ�)��֍�8�׫�JE���ם����h�~��������!	��WEj`��ĉ`�9ېWǽi�&��; 2�J��6�&�H*�{�t�1�7%�����L�������U���Euh�_���=����t�yϥB�p� �ޓI���x����)�7B�T���sS����J�?	ѳ�Ҋ�$
�CaMf��(p�Y
�O���K��JN&���6����"��_��ۼDr"ea,�����c"~ j��s���⁈��3zǫ������N�y-������Tr��]�f�nʄʍo�M�N��jq����mY
�CG�ʠdr�>����Մ���EXQR�����qL�������TS���	�7pr�"��z��A�i������̕��!�ժE�F�����k��9U��=����_�
q���F��ϟ�u�c���7$�2���@��JZx6^D[��3��,x��~-�A�cT�E3���S���ᵮ3@l�J���	Qд���ۮI,|�6g���s��q�Uٗ�=���3ul��*�y�l+{�o�(>E1����
p-=�7�2">�m)�h`D�b�����>�Xφu���K S�׬5P���JQ��E�*�'=��y�v��[;cg��>�U�@<�v��M�C���d�����;�FQ���q�!�9e��R������Qjp�՛�y�'�&Z�X¦��V@1)[&da��T���C �&Sc_�ܔ�;G�F���8��6�D` �?>����8�|��{�8Gb�Y��e]c����-�6�����S�2�uP�~�k!�믋�7�Q�ϑG�A:��Y�P�i�L�l�=x�.W�M����H%{��\�'H�w�͜�a�?��t������+c1	�t{��);��(�zj�\�M!���Wo��2���/����0�OM�$��S\��K���1�;�o!�\Ǹ��,���\��0v���ğ�VG�=<v������BXc_Y �[�I%Fn�A�6��kf4D��r �]p]aVtlux�T�b:��*�ن�Y@�E���o��,���Ihj���Xқ)E�W��y�5�et�`/�d�R��mvN��u�	;pGnΑ&Չb�a��n�䳝�%j�>ioAÓ�'�iG���7x�h�@��K�o�W�O���Rc�J�i$��@bȝs�^����A�8ᜏ��w�hga��Ȕ@g+�Հ&�H8ڒe暁����vH��q�
a\A7��՚"+]r�
SSا����P�:Ⱥ��������mW��y�9Ϫ����n�v����a+7�>}������^�Y�XD-��ώ�۔�7ː��U2r<(g#�ާ��"o�.H�~-�G`��釚Z	H/r��e���,�-щ	F+���%���� cyEr�A����=5�)������u�q#W���D1i9:�x���)j��c!��U>���C�E�j,_?'m5�ڥ3�DX����7�XO�T"����)��mr ��y�a�e}zC�(��SGs���w�Yg����X1����ߜ~�#�g�q�ђn���(DlvI�����⽥Y�Eb��2�9�5�ׯ����(y���Y��
�E��~Y�<�T����.sJN�fɊy_��K0F�CV=���r%�-�4&�G�a��sN&2��'ExNt����B������/���C�LH!2i�S��Jm��2�~�\�/��`7��$�os��"��k�e[A�o0٪�y��c�⬒�Q�?L�6�3�1	���RK7,��x�3.�\^d���̣��6����P(b�V��ؚ��>�g=](��;�0E�� ͓sywj��8AZ�۔���#�2�H��ҫ�GPZ倮���Ȓ������(��lG���i<B�d|o���aӌ�:YjL� V�{	�K�vZ]7�$�e��>)���S���0��y �7��v&�����p=��d$��sT��4� �1KEи���`��S�c�U-��s/�����2���F���L�|�G�?�ӫ$&�Nh2� DVHqm�RYlw+m�r�.9� �i��E������Q��&�B�w&B�2���}pIG8	=��4�R��K�d�� �H�.eL�!�����_��,1|\3��T~��ds���\�3�u�Kvn�V���X�HɌX��Ⱥ�3�`q�����JKUJ�X���\�F0��v����m\v��}��Ie{�c��#T� ��u^Y�9��;`��O ���>W�x7H)��;?
�9�k�Jg5)H�Lf���+��b(��l�7����d��"+>c����B�"���)o˧i?�[�������N�ں�ɀT}���֘�w�f��R�p��lL%���6���h���f�~��Cȼ.��ܭi�{m���o��1�u[r,��@Y�%.:>��mA�77���������h��UN�Z�������+2�Y=}"��S�y�$�2��s'��0I��6���-TW,Ύ�>:���z�$cb�H�_ɥq���D��2��W@���P�SO=i�T�[h�+έ�lS/D���уq�iϱ3�ćx�V���f�H���'`t����|C��ЮJ&ePk]c}w=�w�6擭���$��,"�x>hr�X�Ȋ��φT�ĭ�c��0���w�]�\a�P��Q-�[ᦆ�i.�J���P��/� ��0��I�	�Fq� x��B��l�H^���t�S�qq��B� �UH!�x
���b%�$���4M���I���wZ�G��<������!ц/MN����8�9b��-Ռ�;G�S�+PW���;��w�[��P�^S�`7ܟ�)��EHYd�a�� jٓ��o��4�v/dW�.5��^5u����{�3+�w�u��&��Ւ�=k0��䀥]���z�v_)���8pxж�C��GƯ^V�0j�r(BY�7
frp�L�~��x}h>(M�CWM�~+�H���>�Tt����]�sO��^��T��%my��������{���g:&O��D��]��2ʀU r��@��h�lΦ>�_}O0+��g� Qb!��q�~�i�$��E�[cc�����"����E9Wgv�B�,t����=�W�y�-��I9�p�� "_iu[y-�:��;1���������� �����6aـA�:Ay3cr��W���1�!ʨ� �4H�d�X |�BH�S\��_��_,N���	*�\��)s��R<�ƄI���c���`���Kw��f,Z�t����q/�Z�!��K[Ǵ��~AP���J�[β�����.��h�{׀.��!��[�����F@��V�Y��Q�o<�+���s~�{��6��l�S�L$���;ݳ�t� n/�:��S�ٙoV:�O'i�\�"��݅�a�YP�}"����cآ��js��(���dk��d��.h�R�ѝ�<��]�T�V`�&)y=�A�&&����d��@���[+� \�o���g/��D�/��[~�L��K*����ҷ�Xo,v{��M��H�t ��;@�֋�C��2?����@i��X
,��(+�~?E	y/�_b[C�(�wA�HN�NȤl�sMl�o�`(���~-��y�8Ī��*�#~���� ����3�]��<m�c����ƯAqp~�^q��U[b#UOE&���g�3�!�"'�zk.��|#۷�C�]�E��m!���Ì�Er�H�1G{3�m��٦�3�X�����1����1��D��tcgJ�^HA��ӀK����Wq����H�Q3�܏uK3	������b�3�QH����Y!����(�rm�*��{8-�ڥ@�VE�WT�K�5{�}���������U;����H2��\�\�R�;�����ԢUŜd����;v��ϸt�����ȇ
��~>X61�"~���#�/S�D$ޓ�X�ݕD�P�N ����9��2�9w��R".٠�6���ܜ��'�7��d_�l��'���a�$��
U�_����R��q~����)~���$��)��
��"<����>�
��k��ojI�s�i�֦?�����7Q��Z�A*uQ��4�V#��o���� �yd��"Q�U�.(n{Ő|��1OΟ-762���q�-=�լu�R�ZHw�r��'W��d�8`t�|#m�r���$\��ײ"�NQJf|��"��p5c���C��B�N*0A�Ω�e%Ƭ�*Ѧu?���B�mjw�,�;i�!���u���t���Oo������ʇ�45����v��sTt�m0<���05@���Dp�����X�~� Q+�7E2��K���:p�٫����rm�܊4���p�t%@y���?�Lr�����c�qM �䛷����~�h׍�!;���]���*����%k/1���\+E� �)dI���)�5l�$qT����,�7�q��^�Ó�u�]79�b{S�Ľ�U��'�m?�w��i���Q� ^�;��)�ߊ��zҝ�T�� ]՞�|77Q8-I��̈́J�v+�W����n]��"��A�O㰳VVH�LB�v?iJ��F2��r��E��j���BJt%�3� �p;`��@�JB4 I�[�SK������?�Қ���ހz y��Y�5!7м\p�1X!��!ߏ�8��O�Y�7��o���_��)˕��,~&=� �T��<��s8�G�'�����V@�xS߂�&�	�v����R�F���u��N�"{ߺ1�$2i�0�������b*��P*
B�@�D����#f-�H�����t�n��2��k�2����ĨRu��B�h:�8Β�s�PD�-z�+�l3�MV�Z&���Mx�b�
����E�!oI�Ꮗ���J�X�g���1�A��0����%i�D����g�i=8�9Ê���b`�v�<����xZP2h�/�ݼ�Ug�ƑDB;��W˗�:���;�7t5=Y����9��28v��ru?x����K֩fF|X��R͟�b:�]��4.��d'�����k�v����o�5�,�{s��*h�f?��t2o��b�,J�$JO-�}�~t�6����� x�X�T���P��l�c�ż���V7hT�A4Cˋ][��ϫ�=�o�� ^+oz��}����rѬ�әq��t{�QC��zu.Ǿ�WH�Pt��m���po�P�
j�m?��M�6�{�=��S4b�*"_4Pb��K��e��
�t��.��l' �YV���K��
�D(i�b5t�Su�=X홬x�p��Ix��2.~�42ԞѲNS�ә���ȆN�3�����ቆ�%0#G� m�]�RV�2!��=�m �G|���������Ӑi�n2�;_��B;��i�ccI+�Qi�]�8�OY��R�[���ҳ�i�3���BᤌXz�c��	�nv�����[-�	]�6K��sfܮ�\E���;��P���}HHB�{p���S�J�K#�2ya+��ƾ�=��`v��Xٔ�^d�&Ԩ�)��u���iqjg}g��KT͓�J�cqdi����4�)��2�uA�F<,k��Tl�H_Ȳ�y	6b��I&ͻ����L��r��<wp���ޭ��ǁr+�'���(]@��B��hJKD����^e�p��S*��E)��GC�`m���9�p�A'�<c\�V�un�4jM��f���^�=hϫ��D%c{������+ގM��J��������� �+��dg-M#妆[lS���	W���<z���O?����(n�2ʾ���d{��Y"!�-/���G�WH@q:wb=�>�U���F��I��c��
�'Sو�4�<� �2p�R�4�3�K$�v�F7/��$�1Q������-bd���W/���F�{u��N��Q&R��<��G��#����?;�F���o���Ek5�|)/�$���'ĝ�b�n筏����^�JI���U)"��k)�L7��Ң�D߭7����R�Ƕ�z�"q��m>��ΰ�UX��nOg�--,^�A8��1yl�����!��~�t����ǵ��${b����J="%�����Z��b���R��V˟�����Es�0���r�j�wG�e-o�X��ݮ'@����-Q�����&aS5�i��z*�o�WxiUH�W<x�7�;����q@c����0����ݻ-QJ�wK�%i?>D$d��F�d��qy�-���B΀�F=}��c����2g���(7t5��l���*��j?�=M:���3j�!.�*�Ѫ	R_��hPވU�q�Mna��ʘx{�QpA���2J��;o�\���:%L�N.�j��	}�pp�e��٬>�'2����F��/Xo֢���ӧ������&�<ٳH��(��$��3�H<Zx�ΐ�PCr�F������Z���(0�5Y�i�|OL�v��Y{�/�1�&,�L���펹8�V�SkZ�\�H*Z*A�����l�ь�
�Wfn~�a"��"Җ.۩�f�@�\?�(T�H�*|̡�L�W�6�9�6���J�T�(��8�x� �7����cㆣZ��]����fy��ee)���CK�����ܫ��Q|��'
�.�)�P����aä�N��'��:��y}b��>��:>�o'S2!��|��%����m�6<
���O!pw��7wfV�S����m�?p�����������f>eާ%�� ��V'[V��������T���qb~��K3k��]��:!��-JV�N��^5(H�=��@׬r���\0h�n6ˑ�P�"���nu�<�w�#�rj�춺>�""�����C�vҖ�1�g��&/Ln��3�@7$6UA:�͊r9�{d�pIo	�����\G�`T�EN�P����<��`�t�8�<"!nȤ�qZr�6P�t	�h���$э������fT��Z@��������Y�y_�,�%��
��҅SD��8?�|�4臂�y?�dG���}��"�c�1q[��Z�zEyz3�e�k{"K��u�9tL6�Q~�BL����	^�?n�+~tC����F�b]�/��
����O��x�[1&��U�R�d��uCw��<�|G���/���ʵL���3n$�pl����4�#L���K�V��P���qQ4�/cƾ�N�)	U��F&;�g��
�qk����˱���4���}� H�,� �:m8Fe/�:����Ӛ}Hm>�L�5�R=W��҇�Ȕ2���T0��z�2x_8��fHh}��H�j���	�\���֠����B��*s�(�ݠ9�ƛQ��������ҹ���p�����d�G7y2u�����aB7�zq���`|�v�+�|�+:V�{'Dl�4K�V�Dja����+��5q���1x3y�ږ��M��F����s#�>X��B\N�OD��+�&���H�,3�΄�/.���M�ߞe�T%w��2�Ժ.���A)�e��}5u��B���TA��=H�2�WL�gc4zU���hP�P�/�<ic&�nI��vb��R�g)�<Y�X���^Q*�9V��Y��Wm'�����>���]�򢊺Ҋ<e� �7{��5�5݉���3��
�}�eGbZZ^�P���%��S��b/�Uc�ޟ��	�zGج9(2"�7���*�>�K�� w2�n86���-J
P���������f�<���BEL���=�,q�X�V�&АL��.,��a�	��1��h���0/ȊW��?�*��y�ٴ��e�����. a�~Ľ���w�#�Kj��/�v����@�������i�s�TL�S���d��J��(�;��t�'i�7��&!�Q.b�� �վ8G��;t�!.�����{\6�H��6�O"B�zk�%$�~�T��S�,.��5dX��a,�t i��E��o!�N�-�<E���>�H7:8�i;6�3��{���s�@U�|�nё�HzO�3�m6_��/G-����cn��6��g3� ��*s��L\�g���f� ��`�4����s
�gj���o�S~��r�7"�4��h<�1����!Pa{�0�I�_�����Z٠7J����M�� ��N(��cS�烼iI�>�_p;߫i���4���J�j�=��֛�%�����Y�u@��(��(��VuMZ[F�$��+4*�zy��c��L���� '��5�*��88K�p=ʘb�_����fc�y
x:6�.�st���g��Z���08&I�7�q��%�.�U��i��~B��'�r�D�_�"2�9�g�G�������A�����δ�_����$�O����JN�KIJ?2�v��q����DJP�M�Y9f� ��}��F��s�#��ş6�J2��c�.�����[{�v�sR�d�c �_B �+'ao��`eF<lI=�
m׸l�|P�?ʡ?*á�?
=)ZM! �v�^�t����Q9!�w�Q-a����E�ͻ��C�݁��z�v���(��e57�-���G�ڑ"t����4^2�
��F�i���w��;��W�p�fX�W9��/$�M�Ԕ�+W��+=
<z� ��n�z���>���$�줓�[��t�rZ���c�}/���Y���H��QTp����??����=v�'�����+����4$��'D%�r9�e�(��oM?7�Jxg�C�����h��^�;(�T	�����$3L��.��T�v��D�-s]���7�2R�`y��Z����M�x�,H���Y�{���ƚ_��b1��b�i��#b�^��[��ӟ ad6}�&}���-Ƅ�}<f{$ ��<!���gਧ?�C�(�4{i�常�!��=��1�Q��Ԅ��	n��B��tL����m� ��Fvc�G���Sv��!�5�����$�ڑXp���l`���P�����/�R��'\N�J���Y��s�P��X��x铹K͙�e̽����Ѥ�?�%���� �p�l\�S�ד���C�V���Z4��v+�[�6���a�c���!2�ų������_�y�	S�Lv�ue��4�m����1zU'����]Y�G�˒�0�]d3=�Ơ�ƛ��	7�0����;2�����B+�Gt���?J݄[�]�5KV=�v�� ��n���>a����R��)M5�f��m���,�@W>^:#p֫��$G�lڈ��<����T�#㩫��!KDS"���V<G�ɉ�p��s(e��E8~ �,6UJ�P�E�Ye�1���0h�,'o�Q�9��==�����.����L,3#΢ّk��
�n��l�]�1�8�n'�$yĽH˿pܮ���!}�Cf3���X�A���/���@�s��bڊ$�SG~� ��Z�ox���BԭaSH���d^�'�Î�`�u����yW�O����e�46�#�X>6���=X���h����B�H��'���:��g�������ïJ��m����xՠ��wq�'������`F&���!������#�m�{�w�r���7�1�� �|�d��Z�m(�ϩ�b��ڹ�&is�n��M�	歞 �[��m� Ǌ�6z2TP�#�G�
wsrʀ}��xQ-�sA+;)
��i!�]�To��S������[Ԍ���ۦ.^׫,j{��,�����{l���9�֬�����4�EG����Ys�N���	�����]�<�]����$��Lrl�{�E�j�2�e�:�)�J�k��{��-'D��x�����L��jm� �b^R�~[���'~����l� ꦭq�˳��gDMj3�^�s�%c�2�� 8��}�O�FA�?��*d�)g\	���G>�j��#ذ���z����M*�o�s*�O�C�eF:Vo�D�hW���#��ˬ=l�8f�.��bW�e��H�$Y��΢KcP$٤�O^bۧ.��`a�cD�*���Ǻ>
��������X��A:s�Tdpw�\�%��z��YK��.��0x���W5��`��-����f�?�l�{�7���J¼��\��_��T�oř��������;��=I��Ѻr^ �6���	]��,��)3H뾷��y����F��Ha��l���M�qc�֓�y���6�y�-߂�h`d��u�V -����AN9@se��Z�Ƹ,"�7���F�bP�H��b��!,����L�:�w�ҍOU����V��䗲��-> ����}�x\�z��x��ڋr�Th"��:؍�\�n�U5(��>��o#WS��x��#�^b�lJ+$�����YT�\0�;��-���Q���z�S�;���AA]X���8��������j�n�R�l�=����Ose�Fk66����T�+7AF�ԓ�6 �l��N�o"�g�!g����eI����=b��qjn���B9��K'�9,i"�ZZ��B952N�����)@ k���!3}�������a\�(K����#�}�_���� ]�4J�8��WЕͼ#0���eE�%J��I��%.������/�B&����`S������$C���Z��t�E�Bߖ�c.F�E�0 �Zj���Eh���Ald���:q����7�p}�&Io��Od�d0�|�&b^��̈́V�'#���1ErSŔm;Ҕ"%;#f���S�;��t��5��^�h�.f��R۾���~��i�˼_6����kW�'��-p�[y56r�]"�An
פn,P���Qm&8-��U���O�0�\�2���0��S��;O�D���h]�S_����@(\��	6�bC�r�.�Zq[O�q���S��Џ��΋ٵ����TKГ���V5ԣ�s���*�^#\_S��9����ІPUY0��H	8���/����2��.ηע7*'9G�WyM�\�J܏�ofW��B8��/�6-����f�	m��#s�x�ϰ������؇�`��~��_�H�C�	Y�[n��9����ȃ��"��[��w���j�]T�~`�|��M2�}d<��Dr꺜^�N�� ����j�fY�N�N��[⨥���Og_�<<(����+��)@ڽ�?��JT���XpO�RC>�k�׫&�T N#?�_�:Y��+��#�����Շ�������:�8g,/����G���|T�?�"ʹ�xպ���u��F����G�0�y�do���u3b!(0(|im'�1y�k{X\�ѪB�Ͼ.=��� :jR���?+�y7����i\��E��:2l���ܪ�ԑ���H��z��赱��섕�d�騣��e�иzsM	I��k�E8� \�޴�O�˿�`=F��i��`��,�7���>��an�9{�=��l؟�٢,a�w����Wɋ��������n�#o0���D��./�@O��\��/�Ph���FM���Z��&(V��$n�R"�m��t�C/?�r�-�v�V��B���
� �q䕞�ٽ^�X�R�1u'b��-����C�t@����q �nY��+4\d �W>_u7��>oĿ�-�~g���J���c�<��@|?|�c����oD���녞�]��8��E����hs����X�wJZ9}��2�N�)��/�������zw�r	��֞g!�MG��ryӔSRpY��G�P|!�&��ͽx�>L9�շ�+d�̋R[�}�*�l��Ujl�Ѩ�ϵd�������W{,��@k�Z�E�_`�5i�&n�At��¹��xϓ����7���f���r���Qz&����3}�GnHɜR�տ�ȃ�}gga�9Y5��� x�V�F���$��Ƙ�%��R�����ea�Y���g;KT�S5H?��zu��sI���UE�9_�-��s�y4��跛;���^M7��l�'�u��[����#��}�pw�o���������}&-B=��+�仏���/�!.��CƗ�e��A���˧�l�I_��b���!�>��qE_d�k4��s�dK��9��0ܺ��+n�h/8p
Ź��3ѵ�7��U%5&��Z����غ�:��s_��T[|��a���Qu ���+��'T=�=��ԫp�[K�w���G��z9-\�+`��S~f��D�G��U����fE��Px�����<��Óc�v=�֫�I���
A�Q�5�I13�l�mX'��nW�	��L���=��y v~�fvV�f��PcL���Q�ti.{�pf[�x�.�HW�GhT�y�̭m�8Z���9�pr����:�ƞ�D�`뮻�Ea~�sgr%�;����%��G퀘o�XN�Q
te�Fx �MG���ç�	6&�4*
_+h�tF���Zz��qlh~�B�͍���&�b�ޏh�@��Z�\
#��,�\�m�`�0������a~>T!PQ�T)��Z]Tp�!*��S'� `��kj��_ٺ>��u�����O;J8����
��ɢO��_��_��ܓ���z؟�[n�h`:�u�r���s[�X�J�	1���7�}���WK_����)�I�����&�}�%��V�݋.��u���+%ä��α�-6���󡐊Í�t��Q����T.EJ�ۧ�CG��F��O,����C]���g;-%Q R^�d�w���u�J��&��W��^�zܴ�+4�[qcR�akI��W(�,X�V�@p��J�v#C���Ƙ�Lq�%���������A�/�BT� ��8_9U��=�{w���|�Z��5?�j<��v͍(@���y�������q}+��y5d����/yV�T<�0���k�~���<��ˤ$ћ�X��JL?���o���4	1t�k�6��3ո�8�~�A�Qsב�'"c��b���`;Ag�u���z�͒��H����mu�{W[A��%_�X!2|}�p��~r�%���0d˴�4�nq����Ӝ�1�6������=��Q,\��loc}�9'(a�)v4��!��#����R�,EG�a_D�5%;�1A�7񤑖V���M��	�	c��}rV����K`�{R�&(�e��Y�,��o�!/��t0�z�CU!���x�$Oa�e�>�voNb�x��ijDg>��J�VZ�S�F��ĝ�����!$�.j�T��BX5̻99���9���B�㗿^Q���|�̭�	ʩalx�$UN�P�s��]7Bcc�418���� ��mv��)��JVJ����R�UǷ�˖� `�� �@;W��˛�=-�0��m����]�d)�E���H�O����r=��!z[,�U+z�3X��̄�ے�mG�WZ�䢋
�U��.>��f޵'o�?�?�&���8}�U/8�Hp�1Q1Q6_Hmo�Y}P�6�-����l��;��N���絍�&�y��ւ�.��-^�w�;=Qq�o������L��W DPr�p�W3�h��A�یm��={�`D�G��F��s�� ۪�,7]#F�Ʉ�w���k
*D'�Ee��HTרun$ԕ��� 8<����5q���I��~��� qze^2�a��)4����/�fߠ��C���u��Z���	ˬȘ8�F��/��]��Z�D����v"��B��Δ��͏��G�I�=���tkrE�L^�7<�c�[}[1�j"���Y����Kq��T�}k_��p%C�P�$xs��t��v>�W����>���"m���k����o�Z��/��8����L��C���������Mc��ԡ����j����~�[�q�=V�����w�����X�-��̌��c&���j�i���+�!���U'H�G��nu��q* �S!s�ꪜڅkϽvj�_Z���=X�4�Oݴ�����>wƏ��ե�~��^C���dF�d��;g�)_�(4���>��ٻ�Rԝ�-���98�%J.Kwlx����?�S�%@�OI�@�ㄓ�'@���M���`�Bд�6�+�m6�pL�Օ�4�K$�����r��4��;��&@��=�2��*hn�?_o�O����qw�\��@�Ѵ����#��2*O���3�/�M4�EQ�b1�y��?T�����&���:��8>zNA�>�!�ݽB&kٝ<�/��HgA��
!'�74>C����|��O?�UJ��/!�dE#��`="�;&������ 
��\��p0�X��1�xy}�Q���|@3l*�D6�������}��^6f���
�$_��=S}��;��T|j7��}��g+�07��Wb���`�n*��v%�����[��u`ٚ[�յ�g"@ѥiD�4�=�����Ŭ�V�A�I���9f�R�����q?X�J[�O2Sn��Kb�֗CW�X��I���/�1N�=9��8��H��\7<\:�rY�=���#����m�����z�M"NO��w)/II=j��/�э���"wi�)@&֒GQ	�u�ЕI�P�D�n�x��X����b��f���)�_�;��綱��_�v�u7�[j�S/��qK7�a���Ox�g�6�w���
��́OS�$�4n�g��)	�)��7*�?���dX�I'O(��G�$
L1��;WY�R��ˆ���cn��:)㣯�"��9t����~v��N�'d`�=��H:.���.��k���'A�7��9}����yF�� ��ELբ[�ו����ͱ�lu��Cny�&B����rh�~6�ͨ*���Ԝ��el�� 9����n���]W�,��6��6`i<]��Q���ҟ�`�PI�d2)�`�d�*����Gh�dwc`i�H�F�%�f�����Zг%�^�l��v8�ZJ�g����0dN��H��_���ސ�_.=w���Q�Iڰ���nLw���q��Ch�����,T|��[r�(�����H���ᑄ�
4��`�,W���F#�v�f(4��С��t������]��;�D��Ռ��d�z�ڐ[NL��#G�����&|�L=V�\�͔��|�N	�^��*�W2I#���t\���zv`	�I��M��àȡ���M �O��e^u.z��#�C �I�&�P�D�RQ��c9���辁��J��0ɇ�W����Z2}��7�f�vm�j�;��{*��N���2q�i��ԃi[N����|E�D�F�NNC[�aMj���I��l�hc����A�D��;]��Z�K5)� t�[>�"+���c����M;0�v	���7B~ڈ�
��B�6:B���mmG0� 0����=�aՊT^�{��;HX`gO��p�w�i�w� �� ���{ϋ"��R�&�X���KjÂ��.C 3�2�J�t�R�5��N��<�(�ҳ��'��.�suL�	��Px�^���
?i����aF�B�2��U��(F{"`t��B�ށR��{��#.�Jnr����1?ݫ'c ?����Y�	�������1ժ��Ru� �![M��{���J���y�|V�4��jP?ߓy�Ab���@��W�����A�!C��xƇ��Q�_?<���b��֌������D�����T��C��#����n19g��	��+DT�S`�/�D-᭷1��aw��Cg����	_5��P�%A����u�O� �8�~�S�a�<�� ��I�9,J(d�����х��r�>i���[�3^���̱�nd�,���oBӅ.��]�%��h�h<rwl�7?~Of�\��4��9�a�����ܿ�-.XE4���F:�<�v�a\r��X�I�۵/@q�+���<1Z����m�L�
�)K��ZʆT�b�*C)��K�%��sQ�
)��x�`{��D!_��	t6]����e��]ři�c'�T�.��������^)���r��e�<O?ך$wI���4�������l�e�Y�<���A,')���
�d@�R�+鐘L����T����-���iCS�04r��+�`N&L&���5:S�������L����Oˌ|$w�
��bC�F�����E`T8$�4�Y�_m��x�	-:+ٱ3��$����[�E�<���u���^��������?�kn��J`^ɬ�M�lLW�������'�;/]���l�kU#�KLW��E�Cͪ����\�b�;�"׮���:���݈���O/Y���2�.O��c�\Vl��n��6���\��-OZX{/zMg���(�2р�rg1L��B�=�����������\��b���_2�#j���_�u9a�t�������!�2� ��+�T����t��N2V0=	���rr���VTd<�6��6֣��:>sa�^`+xOH�h2 ��/~1�8^V�����R���1�-�`1�m�#�r��yf�C�2ngd���B vfXP����$#9�E���5Bv#�IW�5��_��Q�a���G�&]u�y��n,��>Q�m�b%Xq���ݡ�M#�5���]�]m��Zqh�4@< [�]Lu�����v!e���6l��vl�Z�rp������g���}]��Buy��%�K2pI���j�S,��R� �=��aZ-:[H+UԵ�%L�Tpbr�ӀUZ�F����M���O�8�M�淞�\lh	7+M��\fO������2�h��n�Ef�ӣJcuЦ�1DI4��~�� ���^u���3���B��k#� �+#���*(���0���N��Z�����<�?��U�`4`0� �gΘ��i6�NѾ�!���ގH�_�ۍ��]\��߻�����^!��UH�[���CPr���0�a �+���M�'��^��F�9�Թ<KS,��58Y��g��b2CSy�Mu�<�!-@1��y��7ͦ��5�Mc_��C6��sgh���3W� �y�gXp|�'ͱ���G-�i�&��otfA>x�J�yZ!pٽP�(�	���J�kE`D.3_�nxz4J��wv����k���+5*�RGt�W_8�I�wRTE`�d��C�Sh�r��=~6�[��
 ���#	Z�C�4�OCGDD�yΪP��Q%8Ӵ��6B�0�)a������0�:���:Wѧ��N��f ��
F9Á�^-4�|��=�T�>s����*L�j�4ԑ��SE�T�@3J�Ae����
N���q�L�ϖ���E���#D����/��oI2�.����܈�����%1���.,��=�v-A$��)6��n���5]�x,�����ڭy�?'q�4��R��C8���P��BY�p%[_�2���G����
��A����vD�N�KiV��h�V�C6��<!�����%x~<j�� u���WW�B��|���Fnʯ��=�nG\� �^:��}o��љ�\�Ht͈��=��E,
�i
�e>́��U$Vo�]N�K�B�_O�^xa�1\/�����D�/󳅬��c?L�3��=; ����~j���nR�N���-�Q1,�3 W�������%0������[,8}��D?$=��u��*������a)�F���v1?�|�U���Pz��0�S��y��_0�?V��^�@v����Og؞+kp��Ϙ�K0� w%Y;G�,�u�w��ݩM�
tK+:����b��hǁq	����G;�Ƶ@[x�5P�m;X���9�}�vK��O�Ȭ�yaD�Շ��e�A�#	�{�:�y�z��\���P�E����<�^�ݶ��'��KË�Uk��2|UZ��֞�&2,��T�N��"�����0�w^�rÁ��^�5�P����8�^�O���;��+c��OC�UҦ�u�0oIH糄ͷSbE�l��z��z�t��h�Q%vT+ɸf�`G�Z�N���4����P�s�8
�s�&{Uvk�6t�!-ÐCM��Bf�n�c��.��լ�rd7X���8@EY��@�Ai�T9�^��5ʃ8ئa3C"E�5�����v��\��T�߇/�����GX�0Y��;�4�k���o�m�L>�
�S׎�"�lS֗r|I���V~s4ڤ��J���$����U����sDNΗ���E���x#.�dQ�-�QំD)��x�$\b�%C���)B��ټj�9��M]��	O{� \ ��MI���p�� �6w��K���O(hS֐�Y��V���:��v��D�H^h�[�{�N����grU����t�_4�<�iS����X�5ԓ��OP��kN$���XA��ɔ,<Է����!7��^K�����XX�;�OO�0� ���?���[� ���k4������A���g�lo����79]ٶ�!L�rP��za����_\�v��s�խ!$"��cJ)�^��3��4�bM�-�'�x�y��*��A�����q�~���k!G,��+Γ�g ����5ˠ̎\r��L�I��JW�ρsm8Tdc��S�+,�Ƅ!�<n�jLM8��T�繓�2z+����CϖKU����l6n"v���ئ�m�������wi)�gm����i �@뀈��ϖ7>���ͥ=a��,#�.�t,*N�9D�P4Mc��&�v�Ht����aH���ǥ���fcS��y*��V�I.�ń��3ӵ|�֣�w�E��v��"����7�Ҳ������̜m�7rV�/�hLt�BT6W�!�Q�t{���Nke~W�θ��x���V�8����c�Q�c_(�g	�KJ�g�o>ģ$�/�Y3�,�^B�B���y�3������s��L��bИ�E�*�7�/Me䬺�zrh@l�m���ͥ[4���5���� �2j�hb6G�[�'w�:��i���Z��vk�0
F;e��� �	��v�������.��"x$�B�(�@���&��y�����r�G�[t�Ю��v�I�w����qs|�cw�\��2�ʼń&�6�Z,[S��Jѧ��x��zb�b❟+p���P�;��}�F�����;i�\!��ڜt�#OL4�$�U�J�V�+f�ǵ�4X�W}�����،ܱ�'���G�0�ie����u�_�����Æ����W2�N<��D�о5fHj�W��J0�ʑ|[!G�,����k�c��J��.-A8K����P�y}�z;s�K��=�X�	��N� �ޗR*�c0z�+�Y�-�� �|2i�.���ni���8 ��?���$���ћ��_M`Cx2o��@;g�Z1���\9��cNcM�^aP슆鶚y!��8rVg5��_�@�'A5K�w5ϝ(ZU�_�b��J$LϤ�k���q�~mKW��B�5����$���86`�Y�{�JT�=/�'�|^I�Zd���X�b���Pc�����t:��QR���*� �OlD77C�ЋR4M�gzx�8$�C�X�NP/4�)�%�#{$^7�g�tp�pi���� ��4cE��|�.�����J?D���7q�uu1�e�J��5���>�H+��Va"��0��u�}��nJ}%MIh�� �F�l�-����6�O��Z���"EBq��eD��b�����;�h������a�6�/�T��P(nt*E�{�K��?��L�p����1 � �1��@Re;'�\[�l�C�U��#N��#��Y����o�P����'�9#�{�@My�݅�v.(��j�&�����o�e�yBA�|����T��5=�D��*fY����8�A)N��'�\_��zӻ8�x�M�s-l�qD��Ðc�F��#=�m�^�+�MmA�}:1�Ȧ!U�Q8��b�^Gn��hC�\\���	�����q��� 0|���G�N��o��N��>A;Z�9}��s}����S&7�r7O����I$��&�°S���3�*���ʡ$��ج�^��^]��~ aP�Ԡ��	��\��F�i��uLA�a%�S%c{~�������8��M�Co����!IY0"C8��D4�'Iޕ���bAq��6�q�n�CO�ә��X9�Z��fE�偮�5����u���ݔc4��,���J�t/v|����*|iOөCM�>�TؑԺd�y��`�F%��-�dHi��V0j6���3�#H1�(Li8�.�Wt���R�]���%��`�O���h_ܶ:3��b�ʏ
�6
�����X?�B ��-Wp'	@Ա8 e�⿒�ZM�g
�I�����O�I�X�\Ip)h��mjP��;A���4Ok;Ȓ��$Orh�˴���J健�M
\i��6�E����R��2P8��ho�p�&�k��� ����Bs?ԟ����l�E�%.��Y�L�چ���k�_��	�g�u�V��67s4�N3���v3�{���pby뇒�$#8�K������@�]��\�#I�~lZ��)�HG���3��g�8l�-H��U(/?i�X2�f���8�5s�7z�J	�/��Cz��in�12}���/q��?MI��#��=�D�;)qjJS�d#x�X�W�-�9_�U&��k�g���	�רm��k�˦�xq�^�%�E�O<?GcW��?���ZOu��4S�^���v<�U�s�?��RS���9�k"Nx�ШFD�J,O�9`�a�}?�<�̗8���SR�ɾ���36���C҄���%�k�g�nJ��%�ˍ��CW����� x�^"��f�:+���8l��@��战�x��;�n��$��L�����j �?��P�Ӽ���j
�m�tQ6v"ʖ�����3�7��t:E�&�� ��'�*X��P'ݾ]9@�3���^�՜�cjڣ'���S�)�C�V���I��ݚ�v!H 6�e����b�MBX�Cǘ��F�����G�G���{:V�9K�e�_<�u�+��չaxU���rֶ�J$}���v�<�ⰹ����ɛOy� �2H�}���%�:żo�}Igi�+c/F�g���]q�����-�]����zS�t,�X�t�$q�R�El�p���Rk��σ\�8�*��g'�7�XȈ"�N'��g��+L���_O��oP�$�=S�&#x�5Wa������λ'56�d�_��_�u���������fV�gE��,.1�Sz�-6@j���/g���1�᧷41�@8��vM&{�0I�&d�ӳ�z�?��
k��8�:�=�H{g��#Ѵ-�j�X �Wi�F�Ň*���&^@)���=&▽�31(
���	L�f���Af��X�6����кzJY��;�}k[��L���驟���g�QT���D+���v	�~�����»�e�-;�㣐Q����rZ�G�Q��|���� ے/�&�+�|�O@VO 2���,m�G���Bބ���G�dE�sb>.c�^���{���k=�����c�O`	����q�a���^��}����+�L�W�I�۱ƅ7���=0^�'��7��\EH�.W@	zk�è'�M�yB�#��K���v�y�-�	i23R�U�CA����o�=W��)�K����|�kf���>��/�_a�w���?�:|��O���sF�=�٧���"C�a�JLiT2r��j��8lDIĪ�_Ә�1��h�6���k�������9�Q_�Sv� �a>5^g9xS�v�)n��U_���R=���,����q��w��k(,�6���Uy�[w�2�{������(`Tm^��2ʜ�l��{�tί���|�K(5��ch(1�KR����pk�M�e�ʧt�R��r�8��hB�G��m�[���YbA�#my��z��g���&e�[O!o�%d��Qf!O��_�2��d���Ʋl���ue��T�m�&��b]�$�k4ā��(�<@�11EE�Ee��(�����2�jAb���]w�'����^�.�A���l�����]�q�/��b��2 0�''�mtr�L���C@Wcv�i�
��Ƽ
*����z�P�rA(lB���L��䉜����!؞��sEɀ�6ia���E���.��� ���lu_�eatWi燒�^�S&���J��>hÙ�F���px���^{�[��zj�L]��6 $+ȰA97'�q���0"CP�e��(��V����Sl$��vbn�0�"�u��ó�����D Q�F?������ّ���_��O�'��R�q'hZtF��\	�v>�03���?f!Hat:g�u�ɛWn&N�%f2/|��P��L��S��?�A/�����] �O�;o�c1�왍�nq�����f�N����}	<��;J$�]�5����j�_�H`*�.�>��IXa��� �Jy��4���h˂.�b�{�"��obv�SO����+f���V���|����ʭIi4��1��%�|(�[�9P�m�yD�����;���Q(:@T����]�{�s5wJ��5���X��K�Lڻy�p�!_`�qݳB�f�0���Q�#�M��s����P
_EG��"�� �ӻ��b��ٙ��R��q.k�Qp�'�a䋏&k�~P'��#\ڭ����w�����C8'}D�����?� ��2��(,��ʯ�v��u�g=����`Y��I�)|q�}���ܯ+O�DYL��k�r��,U�מ脊~�3N�L1���:E��]��i�#��]a��I5-��q�v��;� ��)���<~cn~!���'�2�3���K#P�3�����9�?���R9zp, �r�x�T���*��O9�<�����e#;��P5jp�ΜD]����{[m
N����5�z��Od3�x�T�VLpn�-wt�:�jM`Qq�8'�*o�J;J\V�U�܉���D��&Gm&��q�خ��^v�f��@�4W���7Ǔ�$����[�\��r�VmIn��]����e"���
�Ųܣ��U�\���?�Y��4�Vq�?�Z0�	m�[��Є�T�k��Vt��r +���x��Sy)�d�ő>�qY��S/=
;�׷���R�(:}����,�A*���/�ܰkv�)ˋͿ�-���j������� $�/Q��OG�br�m\�͡�v����!Wņ=0ۆQa7��͉(㢩1���&�����**��^�WS��^7|��6+(!͍�r��JE�r�Z�ɔ�el�a������X��N8l��"�lx���{��m��?B�~��S���ڪk&'���0G:G���<���f[�pS�h:B����T�Vg���Ie�����u�a��N�D�;7�m�u�;�G`ޔ0��b �o�m+��a߄j;/�mK������V F�U��/����T�⍶y�O���&G�sh����{�NYG��XNv9�\��;�����g)XVHx"W�9 .��32�̕h�<������6���=��7�96��p;(޸xY�z=�\��E����u/ �u%A�1����7�v5���_����R2r�$݈9����^�!�Pݔy�:!9R�-�/qUЍ�1��I҉Y�_�m @�G]�Yu�d�h|([~�o`�4�8.|vXpQ�����-���K�p�'�,�vyo��G��2lv:G� xg.�ݶu��)!�&�U
�6�^mĮ
���g��O�}L��ƥ���7@���<���s���]�Y�����i��&�H{b��+o�����(4!o]�Jl?n��[[���Iv˶��u��c�0I��PT�Ao'��������T9;ޥA?���^���\�T�
�ǟ�h%è+T������$'W/5�J����8��PƔ��=�����$O�}��s�G�P�`???����_�L�3/�d�]��t.�����>���e������a%}?��ʗ�~�s�����$b�v �I��� `Z��G��&.��[hT"3qbUT#*(0Ѻq]f��ؐz��N#4+���۵�C�=�>/�4 �ke�.�,u/��v3�xrM�&��-��<P���r�p:���=��{��ݢ��{��6�]�!y}���J�3��wQoT�DX_]z�@�,�����D۹@n��v�AU���@�e���u<]zE3ߙ�!0ge�`��I=%��|.��?���!x�UVlٍOa�v���y*�m�~�ҋ�KL��(=��(�0� R!�{������{��BK��&@�+��_:�I<OR}ƭE؅'i�%��)8�,��ebs�W'}@T�fe��KM�4��a��k�'ay�{t��ɂ���cng ���7��';�m��R�t�9�M�L�m�h[���a��Jl�����[̌ ��	Jq�F5^� 89��q��-9��p��4��o��"n���;�y$����Fl��@iWڝi���Ƀ����h�<]gKv�l�3�+��í(���'�*�������o�*�����h��(�$���!�`f�D�#�Q�����,L�Q�0��-"��k��%���d�_ٛG��P�6OԖ��"��2y#��J��9��!�
���A�^g1A'H��Bd�f���0%���N�1��-u+�Q0��y�z\?��~����&"D�F]oBk�h��du��n{��	km�����������vW6���E\�ȕ}�u�x��c�Ն��9w����x�"\�[]��)��	���|�qK+�<ح3�L���
o�?�0h��Z�K�/�����$v��۩���f@�})�.4�퉻�N]��)���u1��r�c)�k|�O��Ύ
���Z��f=W� �g9�bt��F�!$� �d�}k͗��KtE�����A�
�`�H���`��ˇ�՛Y\Rڒ�8)Rx�$I�<q*��($<��R9�J'g����l��@<N����zH(�ڀ�e\8�Gr���b��	}\Vu9��I�C����>�i��N4BuYŘ i�BC��92i�Q���J4k�劣-?�����l�n���<�/�ty9
� ��p!��i	:�o��ɱK��������a9F~��&C��C�}��E�^<x;%e��^�a������fk�yR/�#Ў0R�r���o���ԓ������f�[���yj�N��@�Y����>���ƈ/\�cJS��\}J72��m��@������$̵��j��/�\�i����Lڶx6�#4��A�dCRa �%�룡<���(�� Ү��t!�s1�"��f����]Yu��U�Մ!�`�&� ,�ߧ1��c����|N��_	I����盲�e�I6��T�X�!AҔ�K�+���������+N~?0�唤�Up�b���V���L��F ����Q��@� wckI� ��: \n ����,v��QW�_+�ځb?O��A̓$�L���AF�
\��ʄ��ZCĸss����<��ʅ2H��ˋi�^���e+��9▰e9�z��������#��z>:�)hy-�	f"����q�5��7��
Sk���x�?ךE7p��Y�\ҝ�ؤ�Ē@�����Z
�tJ�K��B�O��A�]�+SA�[������`���s���KovO�;P�0�u���[w�0��˶ɷ��T�i�����x�X��]��mx���~<�נTZ�o. -��
��z;�Ģ����}W�C�J��Q��̿���iǼ̪&��(rzzNN0E	�&������==��q}+"�D��@��sM���ʍ?�2��~����5�B��X�G�#Щ�fz�kY�0p_�7��Xz�Pи?�X �4qƲ�L��T��g���$������8r�ן⮞ke��_���s+H6J�wy�:��R��*�/�P�uH�g��*�}�����&]삶��Z�P�l��Jo�U�[}@ �5�{d�H�J���8� � �Q! G� �7-U}�&� ���{\K�I�-H@���2�X3:�� �XG��Ku�#���=m�}n5$�N�ux�b� 7���1�<M��h�DfӔj�UcCq�WH���:_2MQ>⸙�_,e-2�Z�sy��5�6-$����ï�`6��xqm+�����?��D�GBĻ�T�3߼�3l\��qr�և:�W�q^� k����T�1�Rl�7�\;m���òW������gE�;��|��]_�ƛ��[��B�lJ�u4��)���gET���߆k)�[{���������u��+�,"�
3�?��f��^WG-���L���/G,�<W�%���@�����t �\TxH��~��D�INŹ$�0<DBԥ���?L|J�z��!'���(M�|x�� ���� �y)YW� �Z'�$,�I�6����k�x����pY�JU�*�E�puw�CC��H�^0�/��Z�����r�gY��T�N���~�a��ow:���{N�/���}FY!�n�`�_��^��<*�9��-!�k��jwM��R�L���i_���7nt�g�#����yjP�3s� K'�5)74�jV�*��I��c��=��\Һ@�%GJ^�I��>l���bzmX�0��B8��tu2}+�M	F��^-'E�j;�v�/�:��*��ֲ�maE\�`���Y3�>���d�X/��'C�%�@��v��Pr��ݢw�z��B���Ȑe>�:���\ƕ{� *j;�'O���5I}�ӧL5�v�K��T����*�k�̚�s��2���Wڱh��j��
Ɂ,��,��dT^h�̗�lmψȬ6�ţ��Q塪!T�� ��������e�*�;q�'��LE���9�4=��u	���\�ɭg\o9�����,p���4�t��O�7��*�7R�dE	1����p���ӥ���ۙݡ"(%�L�]^k�GXv��<���h�q��U��"N���X{31`�neZŋ��}{a%$uh��;��q�l)b�2���Ғ��إ>(����^�F�^�B#ߤR��!{&D��^n����f�+�5�o���5R�nj��)v����;*�R 3-4<�G�Y�������2� ���K7:���_^89�H�V����O���?���/8��w0R�n����œ�Ki��.g��oʀƷ:Cv��w$��.�jm�a*R�u� 1�CzX�H�n�AeUX���!��4��o�r/mR�+ܛ�9"[sQρ�L&,߄��-3�7yt�Jg��P�Ɇ�ZA���t�
u�Q;�<��Ko��E��k��������V�OYN����6�'Ĕ��!�Z��5����%�����C�ϐf���N��g�ȵ&���B::������MFŧ����k��MJ[F�7����/D�������S��}���m(��1��lċ �F�� ����B���n�Z�R1Y,D)��$��=�VQ�Oj7�2��<���)�)4?a��t�
�0�f�\���|hZV�E�� @���?������M��]eP��&Y��SՔJ��bT�w�4H��w������M�!�"�bɞ�H�>��\p�ӿ��Mz�^}p�(w(�pS�|Pi���n_���]	?���CU�N�%����x�m��\�TN��6��wf++.���ia,b�w����Z�����F��g� d�5�"FN�>��@Bjre���]9�<�ST�\e�E�Qe��M�W�YuTh%!�
t�Pw��=ġ~ %y�����r��B؜g����As��z>�x*��|\;R`{��(tƍ����C��q�4�Q�����A�����X�eLB(F?vo�T>�=�xр��~R̷��*_���վ���Y;e]{��+���)ᐞ�L�1BTp"Jx�䎫�f1"���]J�9�J�MW�iz~��'�W�43۞�<<V��
ynU�*wJ���vb�g� �l��L�o�쾖�J�T:)ro�򢳗{(_��+��0B]@Du�k���>��x�H�cUo���*�-PE_E0lu-��*�q����;�N��e�KDH�'�&���`�����|Gq��W}�^
�"`l\�	v&m�P{u��e�t����@N�p�n�QO2�]����_2C�	�^pv|ʁ��G��fG 膘�d��F�P�O�s}0q(�gW�!䠥;>ҡX�f\���Gx��A_F�(��u���蜠+�'�Ѡ����Ҽ��Um;�ڞ�]7H[�$˄>��ԇ�nQMj���>�0������a�p��[�_4�)���R���b��Hd\Q��iR�:��c�y��9��M�x��)�W���"E>R� $�ey�uz񁽠үY/6P�@��ko�7"@z��F�W~g�"�#�8z�����u��>��~�v�_�ee�Lt.͉�a�}9��*�v����X?87BlxM��o��ի�Zh	�v��O�є��/��KA5�b���i=4��ħPK�3O���;C��E,'�q�'����^��옠�������\�FnG�'n�Ӌ�In���~��1!M܄{�d5�֙��m�UΛ�Z:M�7�1�B��3�u�\ ��〚���Ҭ��>��3�"���%C�a�G4s����u$nv�o����t
���ڏ:�q�ڋ�h��I��-��3��3�
��[��2:���|��b���3�W�<�s¶"%�Ft���X��L ̨A��*�;D]�+�Q6��FH$���=km�?י=�~r{�MJ�P�mO�>�qb�=Q�$�h3X�-m�*u��[���8�����KI��㩨]���(����EP�˖v���5&Z���j�����(��^郵����8���Z�������W݇C�U�iP(��B�.�ݼ�AtM�u��j��B�w�i�7��d��<
��g+W��g�"b�1��g&�S`E�Q��̛@�!�E�ý�͖��:|��!�u!�)r	1ԇf���v��*V4h����,�F��k��^1,���=�'�c����?4lO'bD��.=6�����o%�J.̤�� �ے�j:��&�I�]��C`����ra|�8uW[K��9��pw����R���J��i]ct�0��ᤛ��O��AR�9�p��c���
�_Ǡ��W�c���G��TmLH���;wR�T0����q�^m�k����~���'&W��0'x%��%8�y����'���a[1��dΓ����އs���#MX�wf��7�.�zR�����?�����0�w3,\�9�6�Ty�����Ld�rs�.Rq�B����GJ���.ݯ ��G�ׯ�F�:"I�(B�C��n���g�B��t_�Ÿ�����A��[1�v�8�j�,	�~���a�ۏf������FcP{m6�Ʈ�=X���OϪ��Y@���M���M3/���g;����߉K	�g=
���)%����n�!��$ޙ��N-��oL�I4K`*^�]h�E}rw�w�|�{ �zZ	,�墵�/���X�0jD�W#9���9G���|(�<�j��B�[�?M19��#<�7�@ �xQ�LM��8��G���4���ܝp�x�SJ_�2�,ĸM�f�z;���1B%�����yצ c��Z�|@�n�e����QƖ���5x}�"F��j�* @z\�]�4���MъCV��������k��yrz�<ݶ��n���M�l����ms]���綇��G�֐m��L�TM#\��Oi�!�Ǧ��	�_��{��Cn"Ue�1��,��d�{m9<y��\��g��۾ھBq��ڋP�pu�0]����T�")Ƅ���M���$��&J��X��Hd�`��I����Dx[��'?��S�H�����>�&d�h��0��a���x����72x�Fk:"�P�a>Z5y�-�~��CW�:=j+l�3'w\�G��2ŉ��9�2���y�0
{?��Hl�G�ʿ)͛~���l9�7�f��&}�I�՜��=�P�:ߠ��|e���D�o�*C��Aʪ��UFZ$��W�F��fz�3��`�5��=3�����3b�'��=�K<��������!�����ȯ��\�4O�R�`��F[JЦ�6H��K�|׮�a��RhI�A���1�-�&v��UYFw��'�)�p�p��B	i�Aw�@��Mtz�pf�Ķ�Yp����V�@���sg\�ǧ���i�
���c>o�d�&~����۲��̀D��W��d>�o͘W#��� ��I�K�J���5���c��)�6��r�X�d~ʽN����]f�?S�^58��R��dJ�<�EUe�qd���7h1�
�))�a�PS٪S�UR	�ZK��T�7�K���e"w���q]�Ρ�����<M��b��q&u�9��b��(\ɲ�+:%�n�_w��wn�E��5Xޟ�**#`%�=��Ѣ4Vˣ�xj�H<���uv�jd�t�Uh��Z��	n~����~h�[����E�Z]������FV_JbJ�Cs�+X�f�Le�L<�*~�����Gw���MC`��~UB��UA�6��qiv��B����J!fD��+>K�|�^,�#9羵�
�7�xѥ�	�>PE>�y*_%�&�[9]�'5�(�b�V��S�kf"�e]ox���+T=�Ct����F�j@���(�r �C��
����qvk��:5��
��j	�剿�a�K\����v=E�mXjC��V/a�B\�;L���e�0=X��!|���	6�6+|���g��1~�!W�,~�q&O�v�l�b#A�IS"�y���Yxwk�;�5q�!O1��f��dW�����̼z",f�pQ�,���qƧ��T��os��9�8��o¼?'�ޡ.*X����h?�ni5�qVR?^��z���?r�jM,.�9 ��ޓ�(��Rf����.� ���/K���5�9���K��r8�@�w�����`��$��&��HL��%����{������0O�ɪ%vnRB&X�mfz4f�	FB�f�c�����̂��M�M�b�w:�s��^؉��M�J��K���6�},_����g����X-v�u���a��gW���q�Ꮈ2ͲAA{ k0+�� �ݛ�+���|T�J�|{�2g���p��bV��U�s��/q�aI���*>�cD�~n�n=��0�NX^<F"� �ڂ��PG$P��.a��}bn\���"�x<Z��v����7!�*ȓ�_����am����!Z(?2�ڵ$[[H����CŪbꌹ��{��OIyt�N(*�ܩ7�:zROYݹ�hM�\�z�b���6�\�"1���H�2�o�h���bwv��E#泒�5[^[��ay��?J-E0�+��	�A�q �W�C�8 \��3y��ܫ�	7�i��^�>�
Ƣ�HFI׆���ZϜ:�F��r�#c����F�����^�}+��|�Y�Ͳ��4�Z0C��K~������ꉪiŴ*��{(��[�]�"�����|���|��*;<] ~�eu��Gm�@�0��M,M�0\�|R���cit����N�DR�8ԙ��r�U��
W7{����%����T�7ہ���I>�!Yy�I�	�E-�]+��wvG����=�J{bQri�ꣶ�^����\����u1O^�+ZGr�~`N;E>Wɭb���(����v*H�9�):�T�aG���wrږ�;��t�U(a}�Zc��<7b��;]��DP���ӯ���)CN ���"����/b����2�i�/A��&�����C��T�dTu�+��PC�h:9�9%,��|.���i���K���x^�I��%s��W#��K�ĉS��#�j �����P3*�:�z�f(�'�SZ 8ٗLW���y�)l�y�UP��XBI�7�J~D���7d�d�Q��	M�^���٧{g�<ɶ�lo1�X&�PǕ�A����(������W��WF���ұ���{ ���V�8qc�M�u�Y��e�U3Ǥ�H���J}�e�(`�O�b�dG ��!,�'W�do�x��>���9Aܡ��
�]��*��[I�g�Nâ�z��S���U��I��R��c�(��դf�)�Q=�g'1���͋��B:��F�y�$!4����U��}���ȟ˽Dj0�փ8�E�s�����Z+P�#����X�zoV��:Ș"�{[�-���ΰkApXض$~Ԥ��I�a\S1�������lįTv�����R�M�]r��K2�j�(X(D���_�^�tge�+���DrW�ݞ<=z2x���$��X�ｰ��׾�a>�?��=�4Rr}\�5�{! [Ͷ����f�Ϧ��v���-���G��POI�G�9X*C[)���P�W� _y�Swcn�vz�1�-����0���&�ٕN'���˾�� i2�#]�Ai