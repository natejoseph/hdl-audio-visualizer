��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��+.���1e@�5�I���� 5�,��q� �} �ς"��;�/~ղ�A.f��ߋ��4���UfGt���H����1kI��
ؿO���[�{à�Zp_oy��3:��|#�הa��.���%��
����!���\��=fb��p�AU�;k积�:NOFS)��0P�/�
 �R��X��r#�=�-I�P��v��8e*_V�3����.�t�NTK�;״X-�S�͚u� a�kmk8y�Ru�r����* 9E/��k�����d�`�3=&(p�ř�d	����b�yȊ�5��Ȩ)�_��37����-�&��pAWy�/��i=!����^�������8�b�E�	�J3bٚ�b��K�@d!B�t�� �H�G�����i�@)�>�4N�4�=�cR��_�c����n�;��D� ����-���f7Ĝ%:?������_�VUk����e G�����і�R�n�x~܅p��)�^�P�CZl���iz�IE=�k��H��6����/]Zc������y@���:� �4�:�/m��$U2�+=�a��ʼW�iAr���ŽrV&�����?���L?��kJE_K���5m�YuIQ�l.�Fn�aULI��*-�c�\3�(C�/4�c!�zI��1����>45�|�n�~�Ɨ�s�����|e0n�pj(Jz���ޢ�c7�եz�x\��3�| �����UW�������&շ���/_�0�eM�;<ɮv.P�
Y���1AU��
��~B����و�	,�ר�
�%�����NA|�[~[�nJ�'mC_�Š����ڠ�+ ��<���l�p䃲����=
M��F����m2�T��G�j���ф ���6��Ja�kNࢦ�զi �T��h�ޅ%9A3/�	�^"yN*�1�-gy�e���	<MF(KH��eC�`��,�MI��T����l_��0�6������zfT\q�������"��q��W�Q��b��O-�L���C����|~]�2���h[8gZ�!L�kU<h�dk0@=�����S��6#���\����!��QݕT�?kJqh���N�
���xSoëW:��V��X�~|Y�$��!��֠��-k"���Ӹ��
�ɏ�a���5�a�j
k0a�8�;�����e�06��m�;PD�� �o�>$RAn�(�W](+.)��DMˤ� h�����6��0�Ick�H�v�;=��x���B�^�^��iH�� ����xK�jYu���wh�p��3�������"�/ی��x��i��!���(�����	��[��^L��~D��F�r�d�=��^�I\��Mp��O$���8VL�W�h2���oZ�sd��oŬ�cH̱�O�V��9P>�����S ����F����&��'��O���3�%���8��&L>[$��rv�͞����+�V��يt�r%�Tq���9�(:#_���ݶW�|��or�RC�������Ӑ?���u�4�˙pt���x������L����u����n={����os*����Iz�ٷS��\Nu��p)7�VLa������Ђd6�ry栔@`��z:nH�9^A�*��)ґ��asj^���j����ڵcl��̔�w1T�f��7N6�S�[0�ԟ��~H�}h�Y�s0B��ϰ��'L�)!��ZYQ8�<3�zFh�ڄqZ�f�A�՜!��q��X��2.Ah���BH�^�R,��M��V�8u��l����P���s�_j�]�-�T`��r��|^�c*�)!�+kl̟˱�1���b�"�"�`�����s�d ­�Y���w ��ws՟��|�[F�?A�큈j�|*���Eη6K��-G�=0� /7t'R����4*�?GT �z�2��n��t?��G��F���Ve�ƨ��d
��1���I"��
�����(r�f�>�<�h��Af����(����vj�7���w_�G	�SP'%�*� b�d.ӵ�b$��%%��yx�X�q՝���;�!��(&�J	:�|'�	���k*(A dVl��P�R�UY�"o�i���������/����̡��8e ��6*"�xO�}����GjZڞ����Ӝ׫�ps��G2�4
$KF:��Y��{_rI��aF��D8���S��)tU����'rS.&]��I]\L#l��f�٤�6\W���Uȵ٩�EFJp����(���}k�w���5�� '�v���9�~�����?�X�۞\`�@����8��2W�4o�M%���+o�{u�LM���RԞ�2�D:P��a��}�q:P_=��TAF�6���ǜ�#k)�M�Q����qN�Q!�N^H���ϡ�_�YZbS� Z����d ���İ�o]�����q԰K>�X�ܰ��,h!2����'7�m��M�r�-*Y�:NMI��\� �/xi[�&=~�w�V����_ ���<��7��4ZH����%6&_̎I-�	�;�h���� �BD�̖ )u���t��B�+��$��jp�]�_������� C�n��:xT4UN���-�t��@�� �,m����,��0�G�f��9����6/��^5qe����-o&����H�+ݸL�7��īR���GwH���J3C���봤l,-�c�bwr�'Iq�04��J̙��_]�橭e��3��"O7NZ�udv�u�v��[�U���6:���7Cw �!&�#�g>p3���nJ�8�N֖�^�ٳ����J07k��e�Z�g�-oOz�3"��BKϻD���ҫÑ��%M[��-��2L�����7b���MM�K%���[d��~��I;%�M�e ���߃�4�Ղ�*�]_�6��	8�Tg>�LL�
�{_�ε�m���ACeK@G�c	�W��*���|�HJ�s�>~��pL@�X#������r�ZJ��J׳��a���b�m�'�[�61K�ǦX����X�j5���1��e���<tR�'Y�K O�����Lm]|b�L�.b�h]z�q2�e9���#�B/�mWn��� ӊ7�Qՙ��K��~��ںW��7;����ߎ��4��VgT��0�i��aQ?~I�(!s*�r���dvT(��&�K_[��G�-ޭۿ�h��.L՚cSo��P��C�Y���?�W-�i �J�8�@�1���z-��- �F�53G�X�t����������1�Ć��G�X;X��z��b�*Fg��:���JCt�n���>�%�2���g�۱�!N�z���G(�拢�a �C7�M���k��̌��5��uW���`J���mIXg3thz�c��p�c�"��MK�3����}^:��a6�=�	lj�g�o,�̊�b�[0��kT��a�O59�t/,��dE��Dx����暡U�t�|�'^��F	�J�����{����&H�+>|�a^��y�}�B�!�ED?$Ux�,s��X��t���CK���g��{���X���4P�C ��k�\��8 �'x�@��\�jV`ܸ	�l�����D9�t���'��ݮ�X�P*���:�Oy�H�`V���vq�@���� @�#o����~�Q��-���i��2��+���N
ӫt��G�,�|a[6�.�ᣧ)�B���������_ͬ��bRK�כXU��uh.������B��1d_�wUʏ}�9����^Lb_�dզl�����P��Hֹ����:��)����5J#���,O"iGڄ�P�b���ֆl����G#������vY�Rd���������0;9�����i�aT���ɢ��!U����w{�{v��s1�}{nubQ�l���:'l,R,<Yԙb�1'�^
7����o�T�/Ȭh�
��f�4[&�G���ezhO:a���c;]~p�#�Q&�D���ɳ��������|l�6Wr�L:R-�Ԉ
�ѡ��ȁd��dΔ�ե�z��^��I�*Ǳ�<w]��)7�Mq
8.�e��-3у'OH�5��@������mǈ�%��o\sg��������+$�^S]6q�Lkh�F�E�)�P�^�!��kKu���z��Ş��̓�E+Χ3��]%���;��/��vX=:��o�4m��rۦ�#�<�[�y�q�LG���T�o�ah�^ �o���dl��)�G޼'���g�$��[q3#���RA�KI���w�q���b��ʑ�Q>WF�b��Z;���i����D��X�Pr�ƶ�C���$�N��-s�n�tv�_%D]-U���,��r��@�3�4���tۆ��,fE��PO��D��P>C���f!��G��n�k�?��ËA��h�zG"۵��f��\Ҋ6A&ص��g�r>�!Z�g��)�~gO���M����Z(���d�c�O5@W�a�y>l,.S{&���7���D����F����Pź�m/�
�I���U�G�do�n����(�4�N��^���b:�J~(�|Q���/��gK[໸��� )s�+m�(��CL�wW4ٟ���
����U��-�j�^�.���W�4Y"=�i�u��D�����w18k,L~S�0��O�F�w��^1
�b��Ӌ�Y�+����6�oN�)��勮LK�=�k��H��{��D��p�F�D��ew'���S�L^
_�Z� ����R����\"͹経����<&���[�3	��M�x�܍���C�_������7�ߡG��h:��T)��>A�[���5Lʸ��.��"4�nԭ%L3��	�{�����0��j2��XA#��b�a��(���������
)�]p*�:����>!Y�w����â�Y��#k
��Q[������Z����юK�痄	��=n��tj���)���ǫ�Lh����G����/�G����v��?�jʟ�bĶ���%�U�#�q���E��V]eL\��d��x&Gf����;�1/���:�h^�02+.�鋬�@!��؏�r�q=\�/PXnc�s`&����|��<@y�7�V��T�Nyx��`W�X�S�H��t���׻ifMvGᚼ�|�0�e=S�9��(�����^�j)s�^k�������i =	�R����lJ'��+-GU�}��oMS�y���xN��1�և���#�XT���jd]FN����V��S�h�o�(s���� �Ѓ=������R��V���|&�����S[ٔ�9��љV>���혚M6��������;�04#i�bS�A��U����m�޺"qΌR�r§�q���'��ԡ�_��8�.�,E:�#�v�@VT���
���y���2���5qH�X�I��3�JNp�VKZa)��;�=����&�I��Ě��3����z��%>t[_!�`�G�/9x��U��R�
��<C��*:0��zJ{;p��ea\�s��g7����WI~�.�H��	o����N���#� ���K�ǟ\ ��l^'�Z}��bS�/�9 ��Yz�@k�6�r&<L�R�*�,�A�2�c�t��%E��}J���ΰ��j���\}�Q�'̠�֒ς:���[m�Tpz�:��^a2m�d�զGۻ^���#��'�g����~�]O56H���;)�CVr���$'8{��g�����7��iH!�|:DN[���5<u���'#�}��Z».�3u�PŖ�_��g�aRFw_|X �n�j��0���"�����I���)VA��}`��cF�'��K3�.T���6������Iul3:!k�a�Ԝd��PJ)kd�-����˧�n�4-�j�;�е��(	�&�l Ƕ~����/��.�\�^��15Q7SI�D�K�q�*��:Q!@�dJ��r\�Y�ïpа����Oў�G�������ʀ-�5G����)N��z�F9T"O^��)��*�s(�7h�|��̘a��b߅Z�,|��F��)h_�DzJ�n7�.3�6��3c镅�e0n�S�6�ikR��l�?�hUP��7������?&+@��������Q��$\N��'3tI��k��I0��W`�h��(䈠5�ݳq����B=�Ȅc(�Q���{�w5����e��O���t�l)�+ɺeЈ��;��Qx�s Y��T<z2��#�$��|�7�����.ǻ��t��l8�~�7+Z��1��� �o��|�3�iy�9����ur�ˊ�5�`s��H�� M�Wb��8�:�㤖)T`u���Vn���#���8�F�VȲ����Oe� ��m��k?�8`�PR^��6?�.!4��~��L��D=d�������G�E��2�#�{�������Қ��J�\mֆ{H�'C�F�H�㙦&tA�Q��T�e-�Dc�H.f�ə�l�&e2*>,
����eJSn���C��r�"D��Z}s{[τAu���d�ɩ�����S�#���*���WL�So7f�F��N*K�G#��fʯj���'��c�T
ZF�����T�N���~�i��};����m���7:��Z����O��4�nv��Nu���}B��u!#W$�ȓ�!���1�# �ڿE�1�H�YW�0�0Ӄ�􁱄�'7`��H;�ݠ�h�]�ϑش{i|�wm֚|��)^Iv>�W��lx̪qV~G�ִg�Fg��Jֱ�Ʌo�����:eM����p�}�,��;b�"u����F;y�O9�W������1�vm�p̺��)SO7(����,��d|}&$B��o�_�,�6�tb�_�Y��+�Q,h)PŤ�=�L	�s�P���Ie*p�u���ճF���؝�N���;�S�xb�g�.�x?p#2���Ս�k��۫�w�q���k�Q�q��1��"z`S�� _�<��M%iL$c�zxj ��?��Բ{���FG�8uSa���F+���a7cn5R��Ɏ������g��c�����}�[�#�xFɐ�\����W����"ԧ��L�<���L%�P���a�QH�'�}\$bc�1�j"
m����m����5��~�lq�B�<�A�"�M&�N�����b��lC �RzĘu�jT��5�ߴ�z��Lq��t>�Y�S;km���36�<A���z�)W]�y�%\�	�� ���O��j̵�7�-श�o��`@���i�S|�q�p������_�}��z'=^�X�����"b�c�
kU(��%h�٤2K�,n&�ꙃ�(�&)�ނ�֫���n�|ɢp>�Щ82�T|:�����:J����(���L+ш�.��f�範��]t>h�$;H:W��"#�yY��l�K���1i\5���j;!
�R�w�Iѡz�ۙ��D�6�sKL�_�|9	�ajXG!g�܄��������h+���N��G����P���uoI�T;�{�LH�
tao�(���(p;W���]f���yU�XP<!ݯ�6����U{2����=X�s���.�=��8C��]�|���R+
`�����6M)i�EAީ$O�#P_+=���3I�Zˍ�*���,��u�^�L\�����Mb:�� 
U%�8dGۆ�{(9�f� ����@�����(������#�6��8��aC�cDp%��+�����f�{x��]d�6<�D(�Wsh$.��V�&,�3���%��,X��V(�N��yլ�P�y=r�����r�����~��p��=�����7��H�L���̄�w@����>bE��+Bf*�}�j���[7�EMF�2�9���QN)J)PIm{�|O�p�53����F�cH��#lWbb���̣,敩����o�Y��s�>�����U��J�T�H�lr��yÖ�H�^�Vn�2���팇G"^�{Y��'�e jcn!��E)���z녒�%�g6X?8�RX8>y�7�R\��V��*cyr�D�&ɩK�S-r�J���LxP��`=����f������X҅�r�@s�.7��!X��OiМE0�n���.q��^$�q��� ԝ�.�������u7&�l2���C�s��G�T�L21���O7'8F���yL89�&�HJ������Ld&JB�i�+����i���5�S_NKJR���g��^p��_�M	T.g@��g, /5�MG���k���ځ�X�l��<[��~y�6x	s�\�
�+m{_c������|/�:�	���d��y�izq�Y1���9���~�)�^4u�~vX������X;Oe���@[�N���<�V���;r͑���B n�~{zI���� K+vz�QB�C���~��]�u*z�����4]����i�����zϔ��ˤ�<;�J�1`-Pmغ�NT��m芴Ù��A�֗����xxN0��D�o2�c-��Ix��۶^�v+�g���4r'��\� �`w�kg�n��,d�-�F$��(y����j����
����1��A�9*N�D8�`�p�塜�� 2���|��p*̜��/�~�Kem���q,�����"n��P��Њ��ބaW�]��:�?A7�;�8Jo��c���#�|���sOIT���ԢlN�b�VCM�� ��l_�L��*��<�VB����͇yxV�A�3�"d1TE�0v8�[0I����m^�"S�9�o�jl�L,�kw�6��p�:''���]3��D�P
��a�M�_#߲��e���pa��D��<�m�����	���!aN�L�[�Lj��m�X�d�H���읪̷�Oi$��"�s"�x�Zf���j�w�B����>D. �zC4��2���)~|jU]�ٶ@Q�y��5zU��u�Kd��h,r�j�0 7Tk�d�_V��+�D~��x��ɾo0��+Q�[k�`3�� �c�ƃ��\�i��.�U}n��ݗ�V�l������P'��	hWI�G���� �h�����+�3��{�n4q򒎞m'��S,�o�k�p�:O�&�?1i���1�Y�hp-�sR�}�^��x�jH�:׆o�%��Q��G�X�����#$�s�����0�+��؁.���������1d���AI0�,zbZiP���cV{�j�J|��s��*�tݾЌ���%������I���w�D��̦֎zc]������q��=�꜃`�<A?g��a�-������I�$9������`l�#C��H���}`5���)�t8rR�d����""��bu;xc���TDMG'{Q"-�������si��ٜJ5n*�B!Β�������06�L�eIXv�u�������c��b�0�w�k/d�G���C�f�`˂E��wZ8�5�L5M6)pჃp K����5�B�򉎘�nA�ȱ��-+�Z~@6QC�Li���nHD�����ic���	����(���<ߚ�)4�#��/./����(���^(�gm�ɕ��p������%����F���4̠}@���4}u�B�T{�P�u����ƺ�a���hƚ�F�a���t\�S��a� ����::��Ӳ�OR�+	}4!��ȓ��`�����d�	�p�CF����G������E�<ɥ�~�j+?<��cŸ� ��'�e��1q;?u����j�!�R���U4�qKȼ7L�#\��*�@����bs�,mǩ@ �����&#�P�Q�qFiب�Z딜|rۊ�C6�@��Hfa���Tg'k��A{!Y�u�;����h�`l�f���q�y�Mw��0a�8hdB����_P���'��VSՍ|�>5��,�3(ȹ��_7�g����)�ef0��;
����\z��a[�ꅶ�s�� �E�üX�{<Jbz���DK=���Hq�W����-(f/������R�} �jƗ���a ��c��͈�V�)L[�<i]%�*b�ȼ,C\���ҫVXS _6$u�x�y�����S+���(���/���x;�o����9�t{�2Ǚp�ee��zi�!Rb����[��C�R�����I��?6P�UW�I�JX�A���$��H�z�C4u��ۈ�!�}d� 8����l'���XM���q�Xt'��:�f�DM^uɑ����M�^���r�,S�	�(<|.A�L����_	�ç̀�p�39pI��KgGh8y����43�.ʌ��u���^%�ZD�#J_�J󉻔�����߸l#6_e��]��l�e��S!>��K�ۿ���<�J�Ul��hU�b�/�
�����f�hERM@S��k q���
��$�:g��n�ڑz�[N5FVw����(��(��D��=�|^w�L�Z�	�9�y+N��}O���1|Ĝ�z˛`���%�0�?��r*�`(���ѥ|LKw4s("w�k�Z�UﬆMʌ?�]��k�o����V���A�;h���F���`���RY:������:dnۖ���x$�[�e���i���luJ?=T}����T�q�l�� ��\�Q &a{=I�ā��wy|s�c�㶒P�4��Ljx���T��%DD�ys9g�[��CM/l��ϊ��K�_X|cA��9Q{��1=/+ǝ׊z���"'�˿�2����W\�g�G�{a�'�5����_�﬐}��=���ѷ<��ɘ��%:p��T���W!��`�^�G 	y��0F��g@��N�k^��[���ೃΨڣ��Č�%���̣��M��q�%�*5���(�)ю��D�Lװ�S:b��&ؓ�!�/#���[EqD�7�ԫS\^�+�f|ּ�K2I���#��dfc��*�6W�J�tK��д�e;�����!�����l�_QZ���#��0�]FV�Ȇ��f��o��ҫ}� �W��>9*�5!#�0�Md�ɻ1�WR�<x-��S��9[��G&�/�Þ��9�R�mc�e�=�Z�����r����K�*24t����`�M�z4 �tMkT����G��[�ύ�]��e�Q������R��K�8l}��˼H[<�����6}AxW���PJ��؏��	LS�qh�u����p3��8'�D�n[�b�쀊Q���R��]D�`�ء�j�KKVRt�q_�T>cIUE|!D||�Ͻu��sJ�b�(�G�D4s˹�g��t~oN��lw)U�7�	կ~���l{bq���D��B�� �Q,��8�R��O���u|��GZ�u&���}��-��_ӿbG�%�SdBX2�?�¿�Θ»���N�P	꭯�CY`�҅yg��X�D����i��okr>� ]'��KCW��,f�ք)��E��$q�B����Ewu�m5�.�JYmׂN�E�Y!\v�uM���i��̈l�32ˤ#C?���h�Yz
�>��I`U�e�^WtqI2EJ�J�%+��v�4�'{\�ܔ_�M�p5�>��Y�|擸k=�|��VuA��gN�5{��{����G���O����PmT�5��#K�/�&��Q YE�)#-��c�SW���d9��c������8K��e�8���֔g�Ɔ촯����*:�������c��=��rx��/K���n��C&�F<!�?A�-����.tN�?(�P!�g�a=�^��E���)b��=}���5�zRe�ZB��d������i��v;+7\_2�oSD��c*�Bi�9�7T`^or�w��S�.�A�t�i��A�*�-�����r��k�p9���3_����uJ��t�@�P¦C�-}��.bc���b��E�U�R�E��&������Vo!}�[�E�����h�%�PQwj�a+%�.��{zR#@�Q�w�z�W��Y�����������56��:Nf�=
��@�,r�u����c��>F�Tb�W�>�5�do�7ׂeC��7��y|R��]ܠ�oF%=�C G� ;d;/��߁�@|�V%���<+J��Plr?A�M*�2�/���xg��i�2B�#܌�������'�FKTܖT��H8t��Z��0�b�@��,C?���w��@M�� ֌���,̦c��G*�Vқc;eb���6N��j�R��Vq��"��j�u���d-M�fl!8��X���� c���|���?�fkW�b�#C�o��<\��5�^��>���:��U3�ޘ�ƨ\ޮ���w�!��w�ܒ�l;��
Xm��|?�����g�-��^�f:�[���K��6K#�����CQ�#�zz����Ŧ�<kd�e���x���~;�P.DM�a�a�l+��Y���
��W�xm.��`j�[JCXCha8��
M��)�ꩥ@&���Ejw}U-b��u=:��T5��\~��!P�n��NW���qα_z$��y�3���17��N�[#������r���:g����B_��f�+�I�נ|M��㰧vU�>M�'M�l!	���X�C?{$9Sb���5짉q��S�:]���8�\�|���j��ִ5˞�F��y�_
=�߻�o��Q챦k��)֕~L�U1��Z�JO�S�蓼h�y"4-?�	��a�y���b��s�X�4�n%�5�B kX��%=����Ʉt�h/�GF=�� +��K�������(��/�q	��"�b��Rsg�#�SD���=��ُ	�O�Y���%F���Y K�T���$��S��Ld�3:xUZ���V@iG�a�1�*��:ڏHq�n9�vS���jb����T�E���)�.��4��1�=��ǘsN�,����*���/��U�j��x��
<�$s?��\M��X�o�TkJ�yXcI=�Y
���$퐕űy����m!�>�5#ƃ`7�#��F�S}a�H a�1b���Ki��R��t* �2�0-���l]M���t��U�n¨̩Hi�Ӄ�(1��X���x����KY��HhG2�&x[�扈��i�-�4����;�4�b�+���b�8<�Z��έ=��|�E8�[ �N:6��4(L�S'�Rb�߆=&P���␡���l/����f�j`ˋׁ�Az�n����!s�#N�f��ˈ zǏ�J�O1����Փ�A���sk�fg�ޢʾ��Vix��������V9"��);���|X��-G?Տ�|����z���9��]A��2����ݓ	��%E�˖��|`��1��@�vk����3����C�c�[RN�К`|��na��HŘG��Nt���$�6�i(z�"��2�6h:bp4��O{b��量x7���5�yHWr������6y*cZ�2X28����x%�M�)�J�xT�,ϭGѪm�U��+�$8���E�  �.�%L끥g�*
�a$��<T;W��p��}��B �Ҿ����#Ԙm�q(�AI5�^-�/�2�=.�zC�Z�����*�<��r��������x�����"���pK��\{��a���W[�5����P���CP���c��. �p�	���Z9�W�'�-�c�&�;��}�}����U���r�.�|���W�TIW'� -��$�� ����!x�s��8�;��v-^���[ׇkJ,�G�H��D�g`E��O���u��1�0V|��`�ׇZn���N��;���;�ɔK���j�����0���<0��fsc�+�2A���Z,��N��.�K���)�!�����@����o��⑘�4��R��)1�yL����Q<���Fu�t�]�[���T���M`���f��kٷ�5��$��N��޴ʋ�7�ɦ����g���6ܼ	����~����:1�t�}���.�I�hV��8��� *��4���s���U���nP>5��$��G�Lv��k�Mk諤�_�&)��V�<�1?�.�pȎZѺ��q4%z0���=�,��dH����KcNAY䂎]>��Z��Y �	9^�>��v�2�Bp���l�\h���Z&����d�Hy�4���%��/7�jŢ�|/�'q����z��ǯ(�&m6�K������a��E�^Zq�Lqj�J�̚��:>���i�ǌ��y��no��oj�3���t�E]��!�+d��$�h� �U� ��!��|`��g�)>5����.=�������bT�n/����b�J%�蹜��6�����wYO1{�S�:C��ej���N\h�3���9�pU��q�iRJ�|�Rq�Y�xj�;��{��~׸Ie�P�%
��7������#le'��&���p�.�r�+����#�vv�U�+�3�D=G��Gn&�.RÖ�9�K*��ZF��}��B�@����u����?DҮ��w����_�!���N�uHdȇ5��V߬\���P�C~�ȶ*{x�,�rLM����t0AOb���u�1��^3��k��;�#�u�]��}<�T�[ꋤ1f��0g(0"��ԅ���S��r=�y�U �rJ	�uC]*x���Gv��:��#�� <\����8Xؔ-$��Zn����9)!��Z��y���i��]�7����c���-�.�&�
��L���ѥQF<��R���1���t�}8b8����a��3i�.�]�g�P(#k<xHC�nG��Z���#�61�wɲ����ۖ:�iWͳ��c��.�Y�F�0��E�/边�>7[#�J���륀�5��!&,K��8/���殮(V�>����ǉ�@��Z��f8-���ƺ�ս7�U)q0�EM�U�$6Iu7)�����
*��Px��?��h?%���Y��"�n������k����9�\�t�N2$�VZg)8%wΡ9vk�W��`��g�}γ1�yI���g+zIS�ƿ�j�p"���8A'VuF�=;_^"��G	9��ŏ��4Y.�����Ma��b���6�C]f�d	s��U}0���l{ is��Kc!JO�`�RϣD�?��b)kĻ��1YR���'� ͒�=�������\K1o9��sй\ė�{�e�#_c��zX����lxCc/��Dة�Fl��6���@�C��<JCȴD�J�£3��~W��
�RWh�t{A&���1)f�̥��r�����N�j���ܥi�T��u�}�#�М�(U�/ҝ7V,���x7[��T���˔?E����-�x7 �5�r�7��%!2�V1K��W��؍�Gn*ǓP%BZ��`��|H�����fl`�EW\�r_���+*�� a�8:V�f^��k��!�����i��r� ���直E>7ˇ�u���,����=�C��G@{�5���.#`��r���ilys�-q�w_r��L<R"�k�uߞwQ�FR�Q@t����M����ϙ[b��!c��5��E`��, ��t���,��D��*��|��R�w�t2�fYy���5�Be�ЯVo��[�h%i���H5�gN��/��`r%W�'����L���F���Pti��W��Y#]ߪ���k	��S@V��KBV����ed~4��5J����+�ۑ���_Ja�R�Z�3�E��v'G�;�#�z�m�a,XA�kČ���d6�O)0ިṱ�E��`�5dUx{ed-�?�Z>���5��>Fz�=�GV�7�}�γ4T�GiߥZ-v�[Ś�.|=���#Q ��»R��3��)�<A,��[�J�*<�,�ip�����؆�n�_��Q
�I�#��MmH��G
 �Ë��h}��Ceo�ߝ�+)��:I��l\`�W��΍xD���l(�k�dǐ[T�j�E�E%��J~F^ wQ;�[�Z�8�q��1r���협[<�2�OkN��'�/�i�.ک��z�v/��������!����2�O�Q�l���R���`R�|��8�,���K��຅0�����~{<�W���G��V����L�����Ws?�F�.��!�)��[3���`�wB��ӟ;��`ȐV�tnOшƨha�n����Ν�%%�Ӷ�o�+07�3�� q!Ek�8��3U&�Z�d:�4���u���]g�����G��M�BE�m-�ށ�^���>�(j�CũsD�')
�#��'ǔ�D[�}_�硇�	��>��:��!o���f6�?�#�'f�f.�/�y�˯c����r�c��Y<�Pﮜ�&��f?6���\������7����a#J(e&[�aq�N�h�D�<Ϛ��Ӥ�8�KGn��:�Ql|>�1�A��.R�Ր*����i^j�\j
�
z����9��,cr���f	Z���M� ��N4�uX�p�k樕�!�>�0m��S�W�N�O���m�T��N��,���ׄyv��ў���>�gM�D���TL���b�V{@%�ޗ�/W�e1m奴r��B-��f:�kO@T��ǲ_u��I�i��:�ᜩ��w�k��y��Si��i�=�)F&�`:�w[M��ʨ�Ӕ��u�{���I�����C��_;'��b�����T����=`%�2>�W��1>s7Vf�(:��;���#�S�-#�*v67�J+��)`9G��و��rF�>B[d�,x�>E+�ڳ�[m�����9��L��;}�?z�#����3�C{GF�J�
a�/jRLK,ry�3�nA�ĕ\@,��qL�?�E9|_*���[�Me��9d��J�3$�Z�F8G��p���1�fnKcq�tOPK�ê��R�Go��0\'�"�?k�ۋ�[;�	���"���!�,�����w �����̬�i�q.g=�N�����Y���g�˳{�}�K����8 �	��9�ƙ�4��DM�T,{�	����Wh֬=��f�k<��]Y}'��!O�C�P�}|�r%��eS&�����&�[ɒr�?�r��x�+
r����
Q
��)���#������L�%��}�����N�4L�DD6��Q�Μ<D�h������ͳ���5�@�;[X�zv`���v�����:�2���;�f��E"��V�A�"]ʮ��cݍk���.a�����mK ��_�;c���V>��Xh#��	
�%1tt��m�%~/�kW��������A��V���H�v���C��J���j%.�{�@���h�k��?�����U�MF�:O��$�����g��**I�U�D��r��D�ۼY!��vq d /��͞����$�2�.,0-�n�W�{னїtqo���/F����^EqQ�c���A����7���"<�I���o�=$�U�\��ơ{P@���!ZHs��>e��b-��A�ԃ�2YCՊ{�
����+Z[1m1�U���Lgt��;�gf����$[�����������S�g��
�-�u��H١9w<�j2V�6��?��-NC�*X��{BC��ɕr6����k��Fw!.å6 _�^�Ba\c2T�J3�S*S�ᛁ�v���u	InS4��C����l_`���$��^�a�[b��P:����Rt)h:v}L�~��Z(��b!�Q�=��� �{G7.ќv�Q99��N͓cwf�a�y���OEZw#)66:������])��U�D�=V�	�X��d�%��\������*����t:-0�>l�w���H=�1��}�US��Zu������+g�>U�Â9o��	#��
���rO�1eC����)q��U�Ҵ�ܤx� �d=*V3]$Qc���C���3������1�'86Z���;�tA*w$�<�������D�� Je��j�+��kD+�ʓ�e/�}8�z�����-�����a*x�6��I��{�|�2Β����>!r�{џ�k_��.�\� �r���F`�D=h�c%�;���,����B�䋐�"#��7���Ҳ;�DkE��N�H@�U#D�ѲuuS����ظBO�/����#���V�yut�Xs����	&,F\.a�-�&�͡�`._6�%LϺ�&��2h���$_	��!�̨D{B
]�j��9z3q#5y�ѭק"�5�8��4�˾��˦D݋�}�ow�(y)���
��� 6�G=/�����%$�d�)Ѩ~�
�D�	=V♷��-n��7i������4H�%��m>�UN�5�KC����;ڬOA�K�_�L�[��-I�ϧ.Fv"JNX����@�@���P�OJ�+�E����g	�nd9��[��)~�������v�]o���Ǐ������ݴ(���B��g�B�锜�}��稢��,z5xZQ�!좦�c��xȠ�����H���Smo���P\4@���T�DF��������3��.O�J8���i'Nó�gg#=���/�s[��RD�(�@�fZ�,5E�
K�ذߥ�݂�ꎽ�>��[P^�O3��{E0����c��%�Wo�4���I	�zs cI�3s�M:7e����#�g(�,nt+ó��qi�u{=G���UY���Xz���������o߰��cQ�{����D��e����?A���C�D�X��
C�J_O�cѣʖ�6���^;}m�g���s�}]t�~j�MIA���/�Ⱥ����P�`O㹃 ����Z�lN��w<إ`���#���-:Ķwl'�Z�NC���⪚::�x �-@�k�\IL#�v�6�i@qN�dV {��D���u�JD"{�Es�ZQ��~���A�c�'�# Ϧ۩��V��}�,��-��m�5�zۗ���p�F����bw��Z�ki�V�ؙ�sC"1�%��B�iҎOֈt/��f��Ī:���|��D���7����6�$��ˊ�i-�t�Wй1��'"�s���hRU�7��η��a��&��i�X�&����*9�_�˼����2�����"3�Qw�(����T��:s���m�i	_l z����.�!ɭ�_FweReFÊ��J��,���'Q�%���p;r���eej9b=4�4`�"��֪��@�(��5\)TΔ�yE�> PEI~������f�=A�Ef��M%�c�M�M�ii��Q�(�['HI�k�>��������
e�L��O�0R����{��x$+�>]�r0��(cp�K�|��6��¶*X��ɬ\�#�4��x�S��W"����C�Ԛ���kEAg��O�F�� ���e
^�!J��!@h�^��-����>{H>�:���Մ���\+R%�,(sJu�]��[ľ$�`�p�����M�K���y����g��A��D)V�]�y�۹7�U V��"gI|!ĝ(O��g�Ң�(l�Ò���+�|<�-^*^�b��Y�:����ⳣǧ�����#�:�1^�S��K"ٍ���B���-������造�Nj�֬.�KN������ۨN�'�n!ˑ�a$���8ÂN��O�L��zc���fc�c8b���h,~�fwl+a�`/�� @�>NBY�Ѥ"$I63koƼ�_2�\ܢ�vO׍�BGװ�U�-�4b�7�@�/���1j�k7�@n���D�Ո�"~7�B,茞��_����縼�uɼ�0�X������-��\=�m�ȉO���'MR~`-PKLR@'>��R��B�/:l���]� �b�&Pza��I� �%�F����b��9���GK�!m���g1[� }}.!W0�Z>X�6�`��Y� ����'�\i���sة]�}�1��HW��{�(M��^�w�l���Ř:d��5ʖ���6��[��̶���9&]!��%��tl�~y�49Eh���%�c�����g��ht��B�>�ff�}!�«IDG�}HnӽV��#���OMq3>�yTp?$�)�;�M�&}$j��p?�,^���IFh5�4�-\���-36E�a��a��X�b�loU�@�m��6ط����X��%�G��H�����o�~<�k~����0Vz֜�|O�{�9��R�=��\�}�X��瓃S5��U�w��GA��y|��]/-�ۀ������y�ֲ�Dqh��5ܽ�/�[O�A�/�Eir=v W�1sfE��7hD4�}�t�^�1���.���(2��*�1-=1O�AnnR�и�Q^�Uu����6������z���٠�?թ������\���>�UX���F/F�x���ٰ�F�[u��2Y���7\�}����"�C�y�;ғ
�D�)ɭ@��9)�����?�/�;�1s̡_c�1>a�L=*�+��H���`��� ,�̥�>��$�K����{Zs�����_������(B���A��|�t4m�jױYX.�G�����_�� ��BJ�(�t��<�[��H�,�j9�.D�!oI��x��@Nb��"�5�Q�G:5�I���R9��`,H�Ȩ�GD���.��T�c�w�j���;ҷ|�K\�:�\��~�2JȥMt~k���{c���L	-��_�'Ss6]�w�G��b�ƚ��x�]���m"�I8s�G�<��
8NV�ȍ���,_�B̜T����<xX����lÔp��,�G7!Q�JB^C��R9��Y�3F*q���ȝg������(ӧ���p�҂���5�qC�Bl�x-���}8����Ki���ǘJ'1-ʁPƝ�;!��HM��C�p���byѬ�q���ذ��M{�J0оt�L}
'�e��3���Y������S�;���0�9R;D�C��o�S_��{�p;a�oT1O8�ciK��
*S�c9���Sr��%<��heK�:���H��uz�k��.��W��Y��ȃ��>��A|���ʈ��9����/϶�R��6n�fv�xY"�6d�u�C���,�.�^8A8J�0��^
�R�G��SV�y�u�W�yS��X�6�E�$���`���+,�­��O_LH�ކ,)��=���0�i�h"Ӫ��n|��-2���#�*<���[�7����VZ���K��h}Ik�fy&5���G^��_7���8=����EkYA���m�PT�����{AU�{�F�.�<�|��KZxBpeq��D,Rg���Y4m�@��W���lj��U�UX��p�9���\��(�l������އ:��d��I�[v����`Sã�?�d��1���:�iԲ��rћz�Pmv/�b�G�\D5���ဪ��Y�k�s�����D*jo���~/��W�{���O��0兼qvq��0�dܮ�#���K�m���x�y�7@1�84H���m�(��;WT�n�~g��r����g��K�ם`r0��P�`.|��i,r���j�M�=�#$��
�n��+���3����8)�b�	Tb�G蝾�E�/��Q�����,|�ŕ{��^}�c����a�(�`Uɫ'\p ci��ݤn¢X��V���ֳ�m�����M���1�T���*%Eaz:��ޜ�'��Yf�XU�N��F�����B ���;�����Cv�hMsxÓ���1��>�O�'A���=J�>i��1��U�A��	��^�gQ�Q�T�{O���@E��41����|з�d�h��F�hQ/��t�G��F��~���/(2$��7�3�<�6��R.t�ڂ���;������b��j���4&¡Ҝ����U	B"�ިU;�_���X�++5�����OqX.�G�_K��օ\�H%�0IR?��m��(Iӗ��k `:�a����;s����n*d���TV�=�>��(a�E��}qѬlɮm�YE'�� ��q���b�΋m9�L­v�C�:�,�����M,��4pI��K�(U��2�t����vꥶ�)�FA��QQ�&���l����n����7'�h�͗i��"�9�)��V�0��=�55�sFS�^É�+��h��R���"���ҋc"�r޻y�)�	e�/�f���z�4�W��¸70U��ӻ�x~U���e@{�ӭ �.o#eJQ������|�;���\���|zu�M-!l�ו�a}YӠ#����.��=tȥ�[��7��]��QS�ߵ�
Y ��5�N�����o�y:\��)��d��5%�$�:�`h�,��z���<EEI�~>H�~�SHC��/��wL5�/�f>���71��n���B�E�O�4�F��#yæ��Ӳ�c��?	��|Z=��š�`W���W��n����2i,E���H)�����PY�ej)P\Vq�(c�����IS3+�`�2~d��Rz�W��E�$p�J�74�8�9G�W�G�`&�'�{��%���L�_mI̩b�C�y�d\ywx�3Vl��Ѥ���yyC�R�R�mZyk���O�rB�-���v���$E@�P��:����5q+����陉m�j��Dp¶��������Sԓm<#�: gql7�변�O��c�z֗��;���MR�;���O3���Q�K}%@������� ���h�b�Z���
�)�������rgɥ���bx��DvXy�q&}�f��/���PI[F���"K��JsMl�y���2�θ����6�|;Wm��L�cucv�{^sB��x �8�g`��r�<��-a�(ֳ�.[�##q�y�������"�g)���8��N]g���@ߩ�c���_�m�s��䬐��ϡ�ǋ���;a��ĭ~�?:r�1����[$���;�����涪�����kS�&���!�[��="EJu���hQ��PQ��b���P�j��4�/�r�n=m~�|xR�+#��rjH?�8|K��Z����ػ˯p���o-�4���0Q���/y��f����!��)DK��=����)*�}o��]Z�%�b]>s}l�`Ŭ`=2�R�Z�FMPY����X�1�.��쵇�Z�evr��|#������6���;剭D�s-����y���f{D�[ߒ0�DH�/k,�z�}���pqPi���YveP�	���P�q"A$��h�Ǝ� ������ϝ����"�*��T��R���l��]��U������u��f���1u.�g���3?�χ�t���Jz�^<Q��+�:ULܨE) �A�����j ��Sھș8Ӧ�����;y�`ZE9w0���;s�|?oߨ@vYՂ�S�/��	��V?��B5#�ҽ��9\-"�s4����W|��T�O+�?�|��k
��6�O0��N� ����ѝg!��Ѵ 4��Xm�D1WȒ��h��d�$�L��AB�M��%6,k0sX�Y.̤�_�pB�?���ܠ>��/�5j��"Oۢ����6�P�@��	V�yW�x�]\����^C�U�~v�$Q����q/5"��D�>2Y���d_IO):aU��Ud=�-��b鼵G3�>�5T`N�Ib,ˆ�P��+b�n�E�PsW��μпY�� ��=T��o�p�
Hė{O#�k���,W�L�nL6k2��l�:�}����+Đs��:[>P�e�IC4&��Py��QEw�;Y��� ��5�>L}@�mU�1����"2��Y0�i	=��@GE)!�H�� *��ۭ��:1�}D���i�#:J�&:�d� ���p!�� <�1���@E��)԰� ���=�∙������MWf���-=B���4���e�Aϝ��Q�#���!�r�QWa�����68]w����+�^��$��� �b�M_�A߳CB'��='
���u=�P��_IN1�U�ݿpK(��8��{�!�?�^���12���B��LVT��0g��6F����A� 9O�!��~��μ�m���p�)�G�,s�iR��ЇL�x.���^�`�0[�ٲǼQ�b`��$Xo�H��m_�0�����{�>��d�K��m|�Z�Nq�f���0-7�i ��;m�`G��͐����nM��m֓-��c�����	�Fk�M��\dZf�Y�9_�L%�S��dA0�Og4����^�P�����*!�^��"O ��p*�����B��m�9�w����U��ٺ/[��fǸ�6�B4��9/f8J8p���T)���]�K�$~^���{P�L����UFmc�G+z�3�%�dV{8�%<¿�<�A���������5#;CހFmwg((�b��u�FB��R����2��a0WQ�N�)���O���v��V�%�k�AtC�U�;!W���8�93_B�������Ŵ�sH�ms�im�S����t]����)���0{�ᆼL/�rA ���X`�ۀT��������,j`3��}6�
��5�����o�3}C��8RܐO�苑�������ER�!ޚǟ�����x��c��F���/�g�W�?�k��$�5����?Z�ǖ�<��Ș/���;'�H��X��qR͟T<��[��� ���]׶��`5�F�6��6Se��$�����V�p���-�g�F�o/	ջ@6��~Q�mfA!M/��ه��-�ȏ�������: �\'4�Al!L��sg��[I8\\_�k����\����Ԡ�Y�i�������1�H�$�)+�۴ݤ3�H1�9�����;�A�df�� �a�R���\'(w���K@G��a'{Z�|���
?LvC�K4���C�O��W����\���Qp�1�N�&lۨ%���d��Y1�Y���\��	������>�[��(+�e�ݤ����)�4�O ���1�Ȓ"�m��.��ҝ��6��(ds��e����H���c 	I���ګ�^Ϣ�W���w�S��Mv����R=��ܹ�P�^�����	�B�����?���\?�.��MF<�懑LcN���L��F��O�`�(���,D�m�0�u|�?�'��c� ��u�q�D�=��h�5BF�8o$�C3� �$�m��eP-f�E�׎_s��lLh�d�)�
`��b����=^;�z�_g�,��� Ԗ�w���|�7""���Ȃշ�5�&}�+�!Oe���;U��g���+��w�������T�H���񂞢�$U����ry�rwK����=W{����*=�9&��矝�0�f�]ˢ�yN���W��ȥ>��e%^*T]"r��n�cύ�#� T�<B!�|˺��/vqK3	�����N(���Z�U����Q疙�K���Z�F�(t����d�ΤgY�]�v��WyT3��o��M��F���:�`5�jt���)[MC�I~{8bϵ�T�
o���i?��N��6.Ԧ�W��"SBY��J�v�ZIvy9�W��YL��O�ىż�.u��OG��^��f��(���<;���'�BĒ�e�!�}��z(8y{�<"Ы��4(t�3�#�
L7����oAd}�]M
H�O�L�W�΅���p8�����A7bH%���UsZ��V�o�G,���[�U�7���a�����O�U=�.�����O��Ԃ�V�bd�^Re��E�;��:�9�]�V�,�C����̌�"�x>��{�G$�Y��6Ѿ7w`�W>{�ei�)��w?^(�DIj����P��῾�>qIcys��k��:���ep��Qh��T�uJ5�p�댠	摫B�A��&��K���y���Ţ^F�|MQ��FP����_�y�khBy���{ahΪP*�t�i�f�FdBC�5��6�&�-_��2F� MT�o��O{��U�I��'��h����a̬֊ׇse���	�~h����@�P�l���fw���^p�Ww����y�fĪ�g*zt8��W�T�~�6ҡ�=�H_
�x�F���gS�Ai�'�=^���v��1���W�L/ST�)6Q�/dp�:iyo��۪2[ʉ�f�U��o�
�
�M�_��׌G]{��?�;�����Y��E�@8V�5��T�<�MJ�Ù*b����Ǆ�)p(��Bc:���9�L͋ȠHz
o�K>��E!I&{�{�ֱ�njQbL�:�(�q���N���
��x<��q��H�M�%ʢfz�����4�uA)&ɍ���d��+�PǋTg�mh��G��_:�����ڥ�-a,\ �J�'�"�x��)C�����$O�ܛ�0x9������W��ʠcGL����+@!;K �ZR� ��� ��(\�<�ʊ+)!����M�2�H�L@@¤�8A���e%M�r���_}�����A�f��o�����"��y`��h���񡶮��Oc�A�F���z�V������c��9h�t+R���B�YTF&�e���H���jc{����`�T�"S�,\K��U)G�qe{����)/x� o�ao��\��2X�#�y�Ţ�y�j�~��;�S��(�k��I�����xX�M�4����"�x����vud��_��6��������/o����Թ�"�4��@�+ĉ���%��Z��?Q��L�^]o���f�� �J��l��Mdp�pj������C�@U(n��{�ۣB���z3��#&%��Ѱ��	��ly���RUZ+"+�b%23�QWds7!�)�׭G�B�O�G�?;"��{��=��������f�hWێ�S$9yn�/jZ�j���}��ƢH�w�l���?Z��e%%�3�)���P�}�0��n~�腋��
C޳%z�gA����3e8ѱ�I��Ցԇ��׹oi�ƈ	�|M�X��T���q\�$@��f����O��xDN���^7,)z��ݯ�,�������n7³Y3J��°�W�[�Ԍ�J!��48p(���M�2w���I]�b�ovy�DH���*	�}<N��H/���`�Zy�3o(��AD-1/ˑ6A���Epd��U��3յ�`W"@eDᛙ��F�^>,�}Sӯ˜w\���~^V�{>��ߴ�h��ŋ�5r��A69�1	�"x0fU,#�e������	���WI�[��$�����&�箫[�}:�{Xl�s(y���
zϤw�r�� ��oH�&�B�r���F����p�-�j8�&�n���8R��Uo�AakO�x|��ؓe؍0~$f�.U&Ҡ��Ȣ�V_G7�ug��Vm�t4jMN9uJU�ίs|m�ï��յm ��lj��t�It�,��4B�m�����G�/aN�ۚ7��_��%�D���ݧʅ9�f3�`v"��
˗��_M�$'�t���3�L[S��;_@=����9$8�_CTJ'��I3�|�]�g���,�~�����Mu�bwW�(��$S��c�A𑒠��4S���L7��P���S҉��k�XMZ�� ~(�-`��و�3Y��+��7Y��U|� ��l�F��P��_w�����r<B&c�1X,#�',#~�:��u��� ��A@�&dQ�Q&���@��}o�ɏ!#��cd%�7I�K��R~y5�)�^}���;����@Pd�E�{���������<�`7��ƺ(�U�^ܩ�}��^8<��IO���"f^��U��ű��
LX������_�jPL���y5*T��w0�3Ɍ�g��8 �CJ7��52��� ��2�r"�]k�����c��wځ��d{Qhm���P���b�u��+�G�p�4�&+(N�����#W���,$�G�L�s�c�	Q,�?ڧ������_������fȢ"���Yէ�3���  c��f���?�f5F�0���xwXV�^�W��wIXP�n� �/��9
����2�t��΁Em�� �{�QB��`_����H�XM�o�@ժ.O�3�T���E}�+�B�p Bvx�E�UR��x�4��Qm���N�㡈L	���5j�ߡ� 3�;_c�Ŋ��ķ�M3JT�КWh�ǉ�֓U�o���?���~}qW�=�\��NX��+;F����d���G1��؍M�.hbb$��g��:��H�mo�3��)V8Y~!bG��*�ó�a��l���#��iT�%ˆa�,u�I�X�X�먮����mY>�0�|u�����5#1�m2洟o�X�՛���XZ��"S�숦Y��I�D߻uX?v���/d��$�#5����K�e�4ի�94N]G�i�\IC��s8Y���zj�粌��:���GsJ��r�z�U(p
Sنn �ͥ��TM���k��T�ܸ@:��>��^�j�}�n��e�fa�Я�D��.sAL̀�e�H�C M%�}�י�K]���YJ��י�񉤟���Wy�x6i%�<�6[	����	���QZ���d�@���	{���E�J�y�����`�~��h\�H���F"9�A�p-��E�z��hø�>v���ܵȈ3��[��	��%	K]�ΕbK�cXs#�1�� Z��� ��n�}�yX�Nk��ߢ�ܣd��D۞�z.�	��4z���� ���.��-�*0R/拱SԺ��#��Lae��ʼ?�O_�t�\�Tg�
��¼�WGL���
�]�]j@ejT(���9U�#G��%��DkĒ�(��+d]����EE/S�~��̻o�'0�PK[�����(��x�;���]���駩�h�E }���~�A俪��2h��b�v���������)��������g�d�e�y �E�-���6>��&�!4�F�>�.�JG
����Ā�*���A����@ĳ����:g/�/0H�����	��śs�!RiKM���7aI��f���u������L��M�&]����/�э�J่�0*����(ӂ�4�,ܔ��f;�����o���)6=��	a~�{��������\���)<��fj�#�����	���`h�h�|���&�6Y�-�ں�Y�囊�iD�n�I��I�U?F$�ru�����ƫ4�9uR��(�ߛ8nKo9�\�c��PdQ�R�*�Fm�(�G�$� ��[�g���Yߵ^�E�,׵�1��@���
�؃����y�9czzS�O�Dt���-�~bwU�,(_<��y�՜ޤ�ZI�,�;����EK��!�X�y5��{�������<�U>�y�eZJ@��#�;P����-[euq��R���,�Wi̋��_A}TQ�L���"&��0(���Z�o�qiZ}�ID�;��;)N�J*�P��&�.*�n����ة�:��H4��l�b�Hq�ZDф�~�t�UJ��^ד�w���*M]MP��y�{�߹������N��:|zUͪ�FՉ�2��b�p �8���~LuµZt�թlrw ��]/4SL�@����f_e\M�� �r\������C�ɓ� �ڑ�b�A���JႷ�;�W�"��lf���]P�ɡ(ʹ�����=⏽ /q2��߷X
������= ���H�@�6����Z.
i`����@\j>gW���Љ�5���DMi'�[���պ8oY���j1M���K���l�m {�t�Z�rcK�����(�Z':Oe7F�\Js�)6�E5��~��d�lƾ�����3��`c������ߙE��i��A)W��N������X߄��aU�EؼM(���T���Q��&r!}T窫��ΐ��v��ϝW�\�4��RC�"�g��F�n�s1z
�q�� @g'O��<F��C��S� �š�9g��I�]D��w��~$�]Ie�+�˰J�a�=�5�$+�3�B�n�\��l8���ɼ�$��p�
���5]�^�׹����s�Ǳ�9�7!���~�LSor��G���w�Q���K�%ū���ݖ�[�2g%:�Nw��S����
TF�7�$6:T�ñq�e"�:�!}e]s��J�GM;�����JI�ȺmFJ���U`�;}��/��^�'�zoW���Lu��Y"#遘}�=к׉z����`����n*� )Ms����:�����A0j��B�o�����p=�^f��EȺa[�a�,�En�NY�8w��9��:�Í��+�	=����n���I�R�7��Q,^��J�!ϱQ*5^t��N_�6^ x�S�p�g�k��m��Gc�8����lE��E,�_6�gF	4̔�fOz�F���:�KL܁/��������p	Ը�O��&8lq���^`a��7X��n@�\<=��{v����c�
��(pW,��혚�^j��e�B"�nb4W�����r%�gP�l�5�;cP�E�"�dY���g\�Э��j�*
?κ��qִ��I}���4����Xh���+�{�@�<ݽ�4����~�<�`��%b�ܦ�[���_?�5��p����L��Q��(2e�D+hE��q�x�P4�LO�6q'j2��q�D >���<Rb2l��4�Nt)BS�拵�|��P�& X��F��#����a�����]�Ρ��� �(�z�	tl��z�ZK;x���?9�@���%)�9жb�İ�7��2�[��c���
"�>B�rT�˯q���(玩�^i���/+:�Ro����S�!���7�~�&�*{�`���7��b�C�mV�����#-`�3jvj<�	��(;W�F @̊����Rp��3��1�Mk�F�9�2y`�^*��2h,7��`�Z�4��dS�˞2`*lM.a�sPX;7+�^�(v��*���tH���0�;;!�z� [~=��J3����_�"]^�UUK�� �]S��%*�sQn��A���|@>�X���<��Y^>`H܅.�+p
�5��X$�t������+h/U�ʕN����=�#�<�ܷ�� 2�Z#�cHYe�w��\�IM�OC�eE���ի[���ˢ���d��K���!��wW�h��;�13A�/�$3���H����v�g��K��r������$�s����ms�VT��N�����@0�O��^S���ۻ&B�f�2��3'$��}�k
6Ɖ:��(̬��W4��|�1ʉrI�:��C8b���������7�� x@�ӵ@�R���ԅ�8��q{ֲ�fS���*䓄��#}x����QM�G�4���/J��j��ʱѠI���v�["���в��1����	�|�Hq�L��Ȁ�Nlg�����l 	.�Y�o.Ĉ̰3�
�nF$���*�̗�3��M��ƕ��[|=K.e�)�#�Xv��S���r~{Et:$;�$�u���apXW��[����ot�m�D:���x�Do_B_�-��I��ְ,��Ԟ�<$#�8�~c�ݏo`�$��wh����7��=c�����u�!�$���b��p�@ژ�����>�qz�v�Jj�8�c˙�B�8�����k�`� �̯��>���Ց�y�c������g��	A�c��Ԡ�J}%	m��v0�KD85�e�>I��/�Rx�E���`gײA'�+#��5�Z�G_�y�YZ���}�e�8T5϶ȧ��d��4©�\�V�������c��Ϲ'_c����Y7��{�O��s�Pj���N{����r��ii���97��@�]�i*�Y+��da.S�CM4���%x�h$�]�� �� ���|	ɿZ�%Ϙ&�b�c�h��� ��̄�����-�t�������j�v:_>'��d�<q���1����
Ja��Sz�cw-ܑ�˖�*<Q+N����TG˄�K�صX�����Ly�dȯ	�-(@z��5Y^8�����ONqE�TE�s�Cl`��;$y���[�_�(4��n����䨟�s$E]I�#� [�|^8�Z7�h]j��@(��c�B8Ӻ�_z�xq������n�1�+�8���C�J�P�����#s���R֠9��	�t@T�n�Dr=n?�:){�0.O�h2o�w���漗�\�� l���0��X�ס�%�'�4JO��пm�-jT���?�Yo��#�,d�K��1�˟]	fq6=�9j�Z%�&���{��Ƨ2{ͣD�H���ꡎsݧa�wϘ������&��Hk��=y���e�p��/�^��W��e�e��CC��y��F�tC U��/��9������x�7�n�QY|���w�����V��`�A%�_뜩
^Sg�]�ș��o�jU��,�(���]��Q�x�5�xz�,�z�{��"H�@cr[Q��{)2/v8�f,��.�L�Js8t��[槟��n���ƥ>s���H��y�?���#�x�TD�&|%���P�4E� ���~��Ć2t�j^��`c��V�+��n G�4jyc1\�e�/;����_��v�I��U���L�Բ�"5!���8�[}>��$��_Ve'q������M�u��^�׋4�X؁f���߉7�--���1�}C�,/;X�;�8x *U�����Ø_�v~_�]}me���O��`$�裝���AS�@}���L����r�N���(��Op��'�s��!X��J�ǳv����`��ˌ%�v�w)j����W�����G�	��z����s����y�!�(^ͺ�@%Q��@u�J6VىЌ1��Ӊ���TY��X� z���켺Mj^���ʋ�D~H	~��DP�0������ag��%��r�������]i�M�6��-Qܔ4x(�£��1qϐ�xK���w��LP�~�c���d^6���3~c�1O���+��(Z�>��fp��2�,�EO��G�� m)�Uѱ_	�~B	�iYπ��
`%��6���wl�4���osE]�V��(�0��)�sN�z!so��r��āz�G�3��ś�T�m�0�lӎ�9��A�����t�WM�u�ƪ�^�+����'�B�����#�W�;����e�B_���S�Ї�uj�86����-iԎi!ca5�������&3O��1�+ ��4�oo��ɡ��f`oM�T�:�Ñ��~s��[��w���֩�ߴ��h�C9�s.^���K������Y�#�2�r���pZ�ϝ
B�ė��8!h����##i�s�ަ9�<��H��V�n`�C��=,G�?'��	��L�0l.%[�=.J+v<+�Q{���[��O.��6k�)�;z��i����K�� �ڹZ����h\Rx�,!����f��|��F�E��j�YM��ydW�I�Dك�1y�t��<�*�kA�9��C��8����Ź~$ݗg#ܡ��yfI����{�P� �����?F���Z�o�8y�]����J���V�ǖͭ���W�W\^1�^w��^���8�tۑ���BY*w�QI)��U ��U��\�-5��17)��|�r[��!�G9|�V�v�]i3G�m�8",³~ċ��2�ȱ)K�t �m�@��v������=�H���u��?��oE��=�
DRQ�6�U�AÚr{���i�����#�~���� �/^3����H�"�Z�#m��4�
�֧>E����oT����g�i�9��Oe��m�Q7���7U���a�$ǃ����wL�IN"dV��9�Iϝ�����=�ݺ��A�=��7u7��\�qۥ9<\r#����ᢥgc_}�-������7�-�ל��.{vr%����H�x[}���QE↋�����;�|���Ҟɨ��27�PR$����^�,��u����%)�$|�~͘�ù�����}�L�Μ`�BD�o�@Gb��Ŗ. o0(��1X����wt
��Twa�h��|��٘h���%��U�,�TO<�v�(��4nXM��I\�շ����E�t��m�4����Z�����N����O�h�t�Ϛ�dH���,�j��T���+�� �`F���`k�Fy�hU��MH�k!�n�H�j�q�3L�b�ȕ�%5���U�yec�ϘGW�	v���4��RU�VN)���:NWqس���u�!\��"5�f�q�v.)X�i�Q_������|݀{���� ��>JZ�1�GQu����~�g� AV�Η
#����b9s�?n�涫�p�b�gY�����㶃����ߢ��!��1��jgڈ����끰4xR�0��pu� ��:�|�me�>VH��|�m��1�׹xa������ەu9��ooq����������1]�03ij�֥��I�tM+l��r� �$v��f9^Qo0��\���JN��K�zB�5�ʸRT�����=q���I��3GA7�c���J'���
YD���D)�'���U��ey���^ћc�����I���/��sw���N�0�	�]�K� #�w��z���0H���
:O���*K�(�Y���y���Wc�IIvO���3o��{7�Vs��
��lʕ�X
���l��W���Z���+}���?7������,�B����\`�$�/���Ϭ2H�� ��5FQݪ�F���Y�L.\e�e�>��(x���˚y_*�]�J`�46g7���U�ZB������G��%&Pt;o^�-1Nx��H�	~M=�9��
k��6�����ŷ%���+9���b	�I�ز|���媞�(�R<�Hg�B�mx������m���m7i5���=n嘕?����.���tmi���:�-����j�M9�|@<�MԕM1^�����B���t�Ն�6B�vK�qĵ��m	a*%F��f�Zs�_r�R��B�j��R��a��2ev<Du$;~ �I�����;�����8h�璿g4i�F��q�.�)�5��$̢P����Bl 뿢ضk��ķ�=�u���a�CV����M��X�g1&�B�2�=�>��[5:�l�55R����Q��y�y�qh���MuB��f���'�9��r
RD߁�Yx���4�g��W;{vlp�<ɈZ~�h�����8������C;�^��YN���y%B�X�nؔ���mwj�u�|�8Q����*���C��!d�����4��z-`��BVur����%n�Q��0u}f)ub���^�ܸ?o1�Z��,I�mJ���/%'�ǾV��M�K�<>��m�I�nay'l�'ߪ���t�&�Yt-<�9��|��}e�]���+p���&n����`&��j�L�A;+,��A�+���m���%�+jD�.Y�����&[��rcƒ<����aڀ4K���6m�0(��_���X��H����4{6�E�c�#X�
�c�Φwy@���h��P&�/%��ȗ)Nհ�#��M���Bjl�ɸ%|\�v��W���iꨲ�n�r��]M����U=��GF���t���P��	�1lB�J-� �*4��0Ax��V�
�f�{�饋�%0��c���~̬r�iAS|�	�����`�lس�=+p������8�I�,S��%�bp��$������~q1�ҿ&H9jE�8Jg����Ug�4��<�����)�
���(�!�$��P[Ǻ)#P����
b���m�#7�z9*��p�O���>���Yh~BX��CQV�6����7��gfg��Pn�ԫ��}|֤��}��(v��`Ps��N%�`�rś+T+6�iБH���S���ȯP`'�������W�����Xo�eyZ�����4�'mv)��]�S_⨄�N��V�F��C��([8�r0����Q��
aUy��&�{�a��/��9ir/�w��Z�A���n�9�#�E|ujg�8�B�n�:r���N�9ՏT�nn~�.������j�/�x$ߍJ��^+�M��7�#&��2B��ux�9,�g�\D�ڔC��OH�9���tU����vH�kd�d_͡�>�l���Cd%�U���C8��������E_8�kMA״locC�eZ���I�Y�`���&��έ�ĔaW���t*y--�O����G��<W����2k�̏��h�������6���"�E���S�p
L�
�G���u��y6�af�(�j(�@�f�- H�p�-��1�{�G�f���s��s��V��z<1���$���NI��������U?,��0��0���Ճ��zj�Cl�<k�m����z�hU�Z�c���'^��}6F:�Hx$E�3����pp0���0���AE�+�lD2c��Qmݳ6�K������e�0,rq\B�t`��,s���C�l~�2�7-OuÂ7Yܶr�a^_��m"#��_���zd�����E)ЅGjx@,F��	s�	�"���H0�h�X"Kk�����'X̃~��G���A�����s���BI�R޻�p���"6Ĭ�~,U�h��H�>q(��(S`A��G�����f�E�k�#S�����S���n�Ǳ�M��6F�Ɖ�s������JՐ�(��,a`䈢%�m�Z�)�IJ�Ґ�y��sL��ڴo���t&Եo�υ��3:�
NJ�k�\C+9�H P{=�;�;V�Z�;�#�E�l��"}44���{0�N:b��i����J(O�@*�_l��0g�f���efM6~x	!:��˕�n���s�@.�j�'��,�z���� �L����9Zⱅ��b�Bw2�)N���(��M�<~d�ExL��p��]#�;0�Y�ۖG'OG7~�A���3�+}"����xu�r�	�>�C�I�3��Q��!��h�0�y��nFA�Y�����_֡MF#=�ߪ(�sX}�-P����읽&��H߈ÅהwjΗ3�pk�ڿ�*G"n�#͝S�(�^5��J{)�~�:��A�v��U�""l��}Xݔ���уg/�@�UԸ�.�z��J���T}�(Y��G�[f��U�5;hʰ�(ܡR�N�M6��$;Q�8M�Q`/�Sk<�����������0H��q,V����'�B�m{���mC�k��&��CǢ`�f�DԵaS�u��v��6I�jfG��]+hW��&�
0�÷	Ҽ��vCY��^�4s� b!y�/}�''�q�P?Z��U0m��׍����8��u��Cv��{��.���:���Q-]��^.>ݙ�r')K��Z�eV��j�[��j3��W�["8H�>���N.���rZ����#�w3.�P��Z6�����;��X�up��'vYҥV`�~�L.e�cm=2!,5��MuY.`���x�R��M�^gL4� O6�7�������f|s<���1j�����xX���?����QI;��9�,�֗R�K��uF���ģ
'���{#�s�țk3h�����A�bP�k��d�kJe�R_ྐͤ,Uq�h�6��^[��˻$9&B0,ωU�V��-�e�|�[�gi�ۋ�B,T.�З}��t�&vس���1���k��lԼ�9���cc���Fx"lm�cC_��j [A�d��/�}��tz����R�0�Lу1��8�i�j��0H�O%s�=����Z�Q̩�%�yٖ�銍�CT��RSPjJ#�A2%����\<��c"�%w9�8�X42����o����֨�V�`���V�I��=Ï+�.��܏��/qӈ��G�hm�G�'�cgk����+^�F��ZM�@,S�vd�kGfe���2Ws�������������M��D��7��yQ4�N�%ۜ+��c�~3�,������Y0#Sւ)���@���G/�����I��$~�#���4m��m,y.���-(3%US�#;�1x&Fɯ��sE�Fq��o��|�@��
%����ўJ,�2�	%�i�5�Ջ�!�g��#$e���g�I���l9\��救���4�r����e@��֓^&�;��y���]J�Z�Œ��f	9=�a�$���I�w�����B�m�Z&w�qI�^���3,�no��Y�}fd�f�:& ^�&Me�T��f�ٕD��2l2��b1�rع��Z+��;�Dt�X��@��l�$�ۏq@!�����.�%� 9DT9���8���7AS�S��2,����˸�U)ɜ���A���]�Щ��*� �bg�C��A����T.['�yZ@x�l�o��A<=�6��i��6I]YB˨?3��bҌZG�K���`�J�c�Ul��vyL�.���q�W��Ֆl���f�9F�f�����MQM�E�]� �������f�K�6��n"�3�y��S��Y��u�+��,����g`vu�18�Wo#�|����$�� ��1�G�ލ��w��jrS7����25J����t�;BaC,��_kqCz��@�;�(�>�����Åڡ{�Z��$LW}LG#]����G��Ȕc�7:�F����頞5����|�ܔ�.Ci�r�Og=.["�9C~V�F�&0�i�1 �0 �Mm�>4��4������˧�.���(0i�Ϭ�L �D<��~>B�g]�t�85����.$����'��F*D��]G�du�[��3�Y����9<�����T9�p"�+�r�5_�; �%_�œ��,~5=�i�y�G�/���v��+�)��`��}�SZa6x��{���*iaƐ�DH��*��y�`�>�0;��kjR�a��:�<���g�D?���W}����*F!?_QJ=ӳ��'��V��IW�p�ݾP�(
0��@#�O�ꋧŠ���1��ݱ&y��Kq�� �L�ۺ���H��Z+k���Bw�sX�q��g6 q���זvlP�$�m�q1�I(pj-�:��:�壦�
�߅��o�^lp��
m�=i7�s3e�'�%v>�v�q���h	I�	S�R V��V�_d��4 �vyf���" ��0݈�Q��֘Xg��觶ê��,j ��aj\h�kV�%��)�s�B��ݬ�L���xÑ��(8�-�Pk
�>|��E~��)�k�ֵ��׷w-�YՊטl)�ˢc��q�R1����cu�?@N���y_�s�fYOC�Q'~ͻ)���;��k�f+Z���B�j�%=��4N�UH����s�(6���<���b�":��ïhk���%!�#����y���#{��N���I��(e�B��t�74�	�iq��؛׉Kl�T�w���/[�ء���L��\�6&���D_V�q���+n��rK�~_�[ܕ�Gߘ!O�LGv�ٛ$@��`�v�L�u���2n��yw��z�h<�M\�XS�� 6���v����m�y��N��=$g짥'.�N�E1���fE�a��a��*�H�oK�h�+> <mO+��0�'��b�{b�R��a���ŉ�D�%�̈ D��q!�4���K}{�ܴ_5ԯ�z�r��G�UU��+B��o"�\&e��u�ǚH��`��6��1;ˣa:V�c�wZ�7�����Q�!��N�~,%�������T������)��c�\�e�ޤ<K�ky�(n���? �t��#
Đ*�)$17X*P���I�Sĩ��uAZ��UFX��/�G��������z�5	˘�n>L�噶A���.�:�A����s� m�,�� ���l1��R�t��Xhe<~���[-r���<�vgJ6B����$���[̃n�֘I���j�_�"}��^ګ�J�Ƴ���_d͏�����t���! ���S��|)1��.�\b$-�K��#�/Y쮻ӀE:��4��j*,�b����7_O�й���uKذ�f����=3F�P��'F��!Ѹ�Lg��ԴA�K|*���V'��Fa~��t1�\ͦ����n|"��<��`�ľkzGD3/0,�:s�|t�n]�J���y��\����ۇ�{�K��-Ԁ�g0|�IE�Y7��t��Gj�R>c~�� �g|9��g:�U�l�ٜ��5�O���_�B�?̙͐^d��g;�O9�G�s]Ǭ��a$��ޟ��5�	�q�v�L	q��J�����׷c�#%�?�����X�J�C���,�QE�XL���bUZ�������U�1T���y@���3-�����4��_a(o�w�r�O�??���'*4c��j*[A}����a<�׭����B��eC�!w����GZ�u)7�p�4�h�q��	�,نi*QU�?��,�.SQ0S:�+�������u���CF/��眰 |̿��$d��]�(�!$�?t�"��%�ߝ�.WLc��U�Eg ��|���|���l3���Г2��z���<�mv�_�?7du�c�c)Y��� 4W&ěaV^�A*zCL˰ҏ���n�Z1��;�󩎆���_)ݢc-@��P���zY`>Lk��(�,��w���ҿ|�Ԣ�	��R461%���j���f@�C�bVc�Q�'8���k��!�g��2g��G�<Gʊ.�Ƞ��&E6n�v�k�us	�!��"eK�+)p�ɘ^"|Bh���pSvٝw��e����>۝��<i��u����Gޜ���j��聬�V�0Ԛ�j�4�{��w��wuh!�=3C���β�ٕqd��0�Ë��<_�������r���2��J�5������&��R�o���N�w��5�/�ۯ�U����|,��P��	��n�p(�+w��ӱ����
�v�.��e&��6-ƌd�������4X��X� ޥGU�D�|��FT�Y�¾��+b �!���t�/&*�<Q����%v��V��E�����8�G����j:��J�t��>2`����)�]��6gF�84QY�1�KbI�$���yM�E���v��2��MAY� �j�l�m�J��@�Fk@
���qVO��������������d�u[��t�6�d�������5#��0�F�5o*�|�|�P�����ԗ���sNb�Β���0��>j�޿cW?:�]0/tK۩/0�**V��S��h͉�)���*Q7�ӑs6 �I�mlncri�\}N���m��X)un� ��z��_\B�rk���Y����-�'*�+��p!��u��/�����q��&���Ke�97�V`��d���9!���V8|�/��$z�9�b��z]����9S="��d/z���>|�AG�ٰ��Z������SjpA�}��Q�e�ث+e�_���]��&���Jr��%��_��!p�I4�����A���ѭ�j��Y����I]����:�qQ�2ٲ����6VL��F[3j���4٥I���q���b0�.�3�;B�f�m�����D��GF\���%�/xw��.�������V�!j	�Vɧ8J@p'��]-���Ӛخ���D��߹�\��F��ǔ�B�ۥ��#�[�6�2b��&xq���z%�ų\�pd�%tYs�T�`�G��!���,����fgd���i���;>ڠ��V
����˨��T�Dnlm�����I�g�,j�3/��H֎�`=�{svVY"{x{���v�R�X���E|��C��)`~U-D&ߊ�9��y�� �Svhƥ��μ~���7ǔ��]�IR@�WC��'\Jҵ�"�$���(f�ɧh�))���.~�&v����^c&���G(H��J|��J
��_P΀�n�w넇	�7@��9;�w���}�V����W6�p��ﳖ��*���h�L8���sMRJ�;g�}�ę�t#$S`M8�q�n��? �|7U�ЮRu9���T�.�Ѷr��-C#�K���6�	N1��Z���A�G>��P&���cS�p\�4�������,��$���W�lE(��T�Y�J���h��?/5�X���;:74_�̜������ɺp�����#@�syjd.�)C�X~���6���vty����d�D�x��/T�zw�Į��cK�~�l�y��?��&'��U[��H�%r��� �"HӁ��ǆ���-��4�[Y��+-�/���iX���84�3QL�˒�h��a�IϞ��n��C�Ԏ�6�q*���v��%$�"�4���$�[nѬ&�Z���ѿ2�������Αq��\+8>�A�����@��+��I�:SH̒7�dq��U7��{�C��+��b��<!�	Y�c���0xS�3�����ˌm	���K���K��1�Nz8�h1(!7���}eY,F+w�9ˋvH��.@�]�]IS���$x8���LRԃ�$n#�2�ZF%���t�_��(�=0"���`�cV�zn`�e��0a��%t(BYKs�������Mb0渘�yV;A��qg�=�]����:Tg��xc�ܓ��~u���)�fj�h�(��؝�g��/R�XH���>�qOwh߱J�F�@|J4l��3^�����b�^�,� ��O��$�=Ⱦ��Z���결=w`��ۙm�.Ofc��l1ADݖ�\n�d�-=� ��Ǉ�.R~�,�;G@Ux�2St���#��ͨA�\«@7���D��.�����,E�R�8���)xs�EJo�"��۶�3���n�}4�0k��#�꿾��]Hh��yI�ȋI��J�����ҹw���(c@ʎ\�$���;�ޞ�c��4pm1=A�o�,G�CX�x�&ړn|-i�����Џ�烦�E �����h��X[7�����ÝC��O��ԙ4�fU��(�W��<�pP̤�.�	]�h�HR�Kt��=G�c5�Z#WTo�&�Џu?S,�����߼�|���^6���������ܛ "�Y�j*H;�޷�Ȱ���<h&�3�Ir�S��Ƣ��_2�
k�i[���S#���ͣg�L*�M���_�7Q���vz']wZUF��
^�EQPa�Զ��4�b�w�	9MP>�+`:L�q�M ���}�њe��GU��U��Q]Q��6�sp]=FJ�IօU<6<�/�#���Ο�������Iĕ��fK�.B�>���p76���.%�AX�|��n� ,;�g�()���/��,t/�X�ېմz<w����A�u�9� �1=x�H��A��6�b�� 	�~�Ibݙ�G��Xc�o/�'Yn0
�P�ǂV%nڠ��QNڽ-�r9_˫�j�h}�Ez�����]���B��!�~p�<���4^��Q����� �~j�{�P������B�����r����So�]2�3��Y�p���,��7Ŧ����ن�b_S����1Ζ��s��RgtL�+�m��\{']3"�׭!K�&H��&���<CJ�^	2'��L���R�T`agmjDvc���v��Ʀ�O�O���0sa�oj��.�Nw��$6�	��('	8M��8#�7�������5y��7��0)T��C��+Ą��C8�f�w��iw�݋�����E�Z@J�'�L�'�9��R�{f�I�'XI<�z�:���)�}��j��}�y��:�u�<�[Fp�����Q�t�R�qʱ:�A��IkV�H諩lp�-|^�ӛ���%wE��~
�O@g$���Vw�����M��H���+'��b�g4u̴����'�k�=jJ�
쒧**c���t)K�=
���%Ҫ;�� q����OIN��%�9nq蜰�90����!��pk�b�rw�H��pA����vi"��HЖ�_ � ����Z .���(��:zmCV6]�q��	D�z�D��3��!�F��zS�-Yc����|ȗ L���jV����~[��S�<�h�<�XK���!6�ƴ��B�a��<�Qا0"��?�= ��V��wV�zf��gy�|��=���0�|��4A��>�)�_�&Q�*q��#:�n�M#A���I� H�wLzX��6Q~I^��Ԟ��>$�جʹ�Kv����шT+�9�=�BD�7YM��;�=�44[�L��:�N��J*L��'[�����#}��::�ֺm��R�G�����!́;{R�0�p��9b^L��c�nn��v����o��%�usٯ�1���VE��`B$�5S/�\�_�+���y[����p����%���紞�*�rM�G���.`Z`5�H�̕ǔC(��U�v>��B#�0�`˒k-���ms��o�Y*�=�_�Dij�Q�4�h:	���9���-ƺT,P�5�o�꿟�'m��OwA��bsSC��K�d�lj_r�������*5Khm*`w����&}����	�/��o�x���'!J {�m�+�����*��M�^��zm�_�q�-;
�v]���jh↩���3�PZ�\����Mm;	0/��Ru��Ȗ�i��.�H�Y�R���H������k6In�7N`��^?p������r1[֗���M�{o%�E�����)���[�!v����`��[�Z.����?cXY��!֧A�N9����10~�1���,��� �����_�9R;@��T;~��S�ύS�a���^
�G��D�}z�%O�A'6A��[/���Ez�Vl-X8���q���ɿ��؃���<(ɕ���/c9�"vP��I�z�[2}!w�&�He��;X����^�­f>�c��ey�ǉ�[iu����_h$
�kp]�'���dU��n��1Ea�Ġ�g�id�(�g?q�U�*w���4Nh��"K�������aX��P�Q̿2�]��{��960���!
E������l����� �Wt�~��èn��X*�PRB!���_k=�N�)�몁dɯ�[�t [GE/���8��l"�ׯ��^l@7fH���ӫS��/�d�<�]��b�%w�i/w���ƌ�c��E
���:@���<V���2녿5�[#ok�/,�����P�H��G��^�H`h�D ՟B*T,AJ�g��=��m�~};�]Я,�+�^�(�&�25�c[=�Mo�̒�i���c|̼�EL��s�!r({L�5�C*G��������&�wDn�[,
�#^�^aM$�I��;�/��.T=���/1��j�����O���[��r?2�T�'e��VS�ni�[j2��}$)��"�\A
�a�`��-�������ұ��_,9�S����(�s�Bp��@���	�H��.��$ə hy�%������o�X��y�g �.dc���3�hG7��E���Z���Y�W�F�Nׅw���;P}@�����W��^����տ���u,ai{q6��-�w[���e���1L�f�j�2�/�� ��Ю����6�Yܞ�ɟ"8���[�GC�K��sEPTgz:;���ܳ��C"{fn �=�Y�t��D�|`e�	�i���Z��`2��	WH<�f�ꡯ#y&���b��\�r �Ui��Ѳ��4��%���W"Tr�o�9QPMb��B�eqܖ8W�N��G���]�ު����`�o^`�R�[�P��\_\�[����o���k!�?�4m�3��gYD0%�/T����N
X�Z�4.Y.53��	��)F��a�#�� �ˉ�D�є�O��^��,�m�����7er ��)�ѭ���_~��lD�Mj�\�8����;W�@�@: F� ��'ݾFh�ɾ�Ẏ�3�oS�N���̗���3��.V��u����[���}Дwy�u�D���}&b]ؕ᝺3Dm;����fޘ����_�!���1���+�t W4�5���Iv�Y.\�u�ٍ>�GCVP;.�}'>.Lk��x!�||�z��q�j����\�U�T�Ds�e�b�|���Evo�Z�*���?T�DN����a཈�T�
��MtYٴ"�$��	f��Ǡ�L��(Q�����	C�'� �������� VK��J���9l��;����N�"��L���jUK"	�A?�P�q��A�NG1���j8	�wZ-��+(1�T�e �NI� �hh��� ܙ���B
A�]T�򍾞g2$gG�ad�X8b}A��]�f?䄙΂3�1<����u�b]�ߙ�'��^���8-0N�&�F�j�S7,��L�7@��=�[��TWU��i���P��|�j�q��L�1X9�_m>��7�&�S���^�2#s��{)�Z���)�C�B�+�=wx����3(Fr�Xn��D�N#�c�
 L�ǪS�O�f/��`9�;dC}ߖFh�/��Q���N��Z{W�n�ͳ��̗�����)�eVp���X�T��'�n��Wf�'O�e82u�*&��?��3P���qt�����yBzU� v��B�$]�`p����,���M�&��u�O�TI�Fl�+;��6{M��w��l�t� J��X���
R#sU�f����Lz��h�z�i��Q�i�O�8�p4�TfV8�=�bU�;�g���%Z���'%$�S��^M���cR�$�����ƍ(9 �j��9�-F�>�3�jp�"m�$�Qv
�$��j�r�_�����X�O�r$��Bl���I��1���B�?�r���)�b���|-���Ce�4bJudޏ;k�D�H��	���X�u.^�e�Z5��P�Q'�Uc���5�S8�˒ZfPG7�^�]�Z�'�	�hڣP�����9AU 3���(�t�S]�'��if�9
�� �K��0HnHS��̻{(��'��T���?�eO�C���I}����
�*j~� s�e�)�$��%�����	��_�(�͌�����Qn�(�ԗ�xpa�32e籘����=��vU�YU�1���G�Y|�_q+�E�$�h��o�<�P��cVcB�y��T���W.���v�<l�����I|3:�US����� T�7�'�<��CqG�"������T���3S�9�G	�W-���(?P�e�2���r�#�
T��$���~�����ea�%�BWN��FE\x����JѨ�:<r���e?e�Q���yj<x��y'�B��B��cX�J����(�w���6����i*���B�;�6'���זNOg{,�E-�.q���g���.[٢dB�@-�bc-6'>�^V�5���9Ɠ�+K18U��ޓE`)��/������T�E��u���R��I����fsܵԛ�9�P���6������~�ì��5"��<�إ��f�Z��!��l'X���*�n��&�~@�a@�km�����3���w�8g�{�ԚU��o�=���Vǁ@��_Na��Q������O�Q�t��F ƌ:�$DoJ�z����L�Z%���B�������j���3,V�[rw�V� ٜV_z*��z�«�R���玉B�j��s6�F����N���dwV�1���>��gW^'vu����_�|}�y��[~.����\۝#�)�d��^T����P|ta�3��?�.Q��ܽ�l��l��wrsQ_��`��M�	���ݷ�.��ns'����h[w����6_.@�%/!�N)E|�D��zcR�.ѩ2���v5u��9��z����!�><��ť"�Nh\9^]�#�W����'��qs��Ӌ�֮f��[��Q+bth�Wg��"�J��Ln� �O�`�ϦJ.��E� �k���I�J
����PKa۠�.*���L�Er,�B��ߓ��R��3rM."���6�o3+�ȩ���GJ�Wc�����*ll�m��z�%��� ��G��/�`"LD��Weõ�nm;�O�(��Gw��|�nH�< ��=�J�4���0Ya5Ȩ��V)�7����ByŢi5�b���cZ���z)7&;Q��C1/�ȧ����ƽ�'��aa!]v�o�F�AjL������y������M"��(w����a�$����5�V�.�����]H�i����#N�b����ѿ��n�r{�R��U!��}�_+c�՛V�+,�vh�\gn�;�f�5��"K����y 4,����P�@��ˑ]����jf*S����Zt�ߚ�#�eS�@����m�)�X`<vn\ҿ�*q0UpX|�)�08ի��Pw��@F<]��'cU�*ܤh؟��..PXiůN]�D�z;?/�H����ڳ���]�G�c�F����<��+�����d�h�I`<YU�Y�"�>�!T%Y�!�n,�p�H]�ć8�)��0����>�s�K��v�4f,i�uį(]��k]:=���@*�I��/"�o�l\�����b7Og"n��@��EinWW�yA�2l}�|�UR_�p��Ϯ\�"�{���LJ��*d`�m��ݜ@��/��T��F�aR-��|�=���C]�9P5ǖʞF'��r�K�hIO��R�-��B�N�2�W7��X
��8�������W�bh�� ��gZLEv"�4I�ܺQ�W�ak��Q�5��[O�4��PN0�3w�h���/������r��**�$��Tfo��Vd�p��ހH�a�/��z�*�./R�fљ��4	�D(�H��a*���e�k*�W�;�aj��{��G��Q�9�|�&��T��<��C���m l��@8�F�����u�h�F�
ފ��y�����}��Y��.��;�$�.8��FP��r}g}�"z�y�ș��%�xs�b\IO��l>Zs��l�d�7��tF�1��&o�x�.�@��f`'7;��;�`C������'��u�n{��)/`�Q>i�u�1�b*�7�k��i���g3)��	,�ɓ8z\�i�C�AD�o�M��_U��]��7T�Q�Ee�B��&���&�S4�����M�`�:��v.��iy��:IB���zo8F��S8/jT���07��+SeC�A]m	'r~/qv���a��*�#ڹ�$���3ٹ>2I)�@pv�ʣf�Wo��S�+���^'���{߈���}T�ec�&�.���\�Hs`C�k�췲z���z�e?���|6s_�Mt a�z��<�{a��#��$77N�q�k�����¿C�2�4CD���Z��V�)1�b���ּ6Ʒ%��w��{�N�`���Or������	�^R�q`	�()��Ud�������q�jsA�O�{q�9C3V����-U>�G4���(��x��s��q1u��Y���{�	6�-Sn�<w�T�b�V@�3�к���1�����\=1:Dx��K�î {r�?�K'��w��gBm�9��}���B����O��(BA���C�N%���@0�}w�#Қ�q��7@�������}g�UuHge/�l����Gs�gs��	�����y9�}Hr���,����ӶI���\�|ғ".���F�S���ɖ8�;tv�&�c�br�FB�]��ݻy�c�Q|���o��y����5�m�g� ���g~� �����w��$��NN
����ց^�̟V�s�9.1i9A�����ȁ5Ɏʟ��d�cN���ܦ�:���	R�y�f�����6Px�"��B�S'ؓ�@�8��9��v;Cu�8�zZ��g��F�oE��%������TM�Y�Tz�(ϻ�K�k}�u�7�Ϲ��O�#\P�e�bC$މX��Jw-�Mhؑk�U��T�g� n�,��%�/K9���OR��c6�B8��b��?�w��s�e���>+9�=�>�jܛpCc.�m'k8�G-F@�Ȱ�V$a7f�!�]�t%�׃�	�h�s�4;�Zi�\J���$K��lt6���K��LF���#8h�������`3O�@	O��A�� ��m�[�g� ������6@_NA���C7',���O�ߠ�ﺛuU ��6O�k�t��F//�������0�7����韎>���D��vb��&�����Uȩ<i�
:�W�.�Y���L8x����m��Ͱ1 �����KJ/H-gC�r����e^dR���|)����^$�o��r�ʇ��:�[ ݢ���� R��9�V�A�s'��>V��47{�g�]�x(�����X^f���G����Kl�(����2�O��c�S���A\�ހ��2�!�?{���׼��s*Y&����޴-�FTNb}h�;��Uܮ��ܣ��)� xXN��Z�oU�0���n�+����ޢqu8�x4��A���r�nB{,��uG%�.���}j3Y�2�ݽ���mvΊ�F�r�v�L_z'g���~�z��:�eb��M���< �5��%�!�9Ũ�3�p+�9������&���d�S޾�D���\˙0t
@����^R	��̅�X
$�����S����=��w^�K�o���p���~��s�mQ�`L�M9��f6�K�mF��!&�됺��Lb�R?!�8����2���dp�Bv��0��|��&o"�n�8���Z(���P{_ɤ�����n�Zl�M���έ�Pvw/$v������|-����A��\jNr�"hQ��0�Ɠ�����z{ު5��A;U��*0��F�A���6�*q�6?�L�?�>4.zNX���Ʈ�]�e�0�Yv��5�~
=S��d���A9�n������`xMv�9uC��<��_�(U_1�WB��fQ�r#��\���6d�������A�FH��H	�!�.�״�-��.IN��K��5ehc��#�7��44����9»�%��IȂMX�.8z���Ť!�o��n�2F%�c�����J�g�B森����8��`��%)�ﱢ�~S���DX�T\�؄w���_a�&����?�p��cz��j�i�Ҧ����?�&�n7[)�?�l�]��t)R�\f�U�16F?pN��#��k2m���w/�����i�p���^�&!<��@�6�&_�z��C�0bT�A�޶	?���%~˰Z�z����.)K]��H�k��X�������ڳ[O��^]N�7rRw/�$�����q�<	�<2.q�{j{ÿ0a|��?[���4B�-{��J����::b����@v��筦��*�_��2����n+�/��mE��M��J�٥��N�����6���A����ξ���t���0��l�����R$��]�K�:�H��V7�@�GlI'�Q�x�=��3)8�蛒��[�k�4�����ޱH4Exi!`U8"�6��(sJċ'G�󫶋�4�3�v6�����_��Mw������Cxg9?�BS�XW�M	��mrK̜�,�t�+5:��Q%~���6�,��uN���-"(���3<�2��@�y������ WL�0����gXƒ*��TI`q�P�/�(yA�Ld��(>�L�&b���0�m ����X�7�=$����_{*:L�)���(��4!`�bd|N�ـ�1�L s2�N���H�6w+O�(��<��@���/
�+�M�$}�� E{�Դ��
���՝rl��W�:���.�N�W���n��-6�����A�[?�:s���kYÛo$�ҍ6?[�n�y������Qd�
����n%5��qZ�y�_\�;�J�jl�3s@����
�i�0$n��\&��Ɓ�\���yW����*q�,>[A���e��G������[v��29�n�eQkg���&ػ ���~J뙭e��mw'(�M��H�qx�3�UTP���DZ�r��ĶB�[W!��Uh�/S�"���O&w4���4����?�ˡ��.��o0'}<�K�.Gܴ|~o�yd<3����+���s/��y��C���?*�0�#w�?Q��s�i�$i��b#8쐎�_���;�v��֣��>y�����U@�w�pTb���?��D�z`p�`�b�L�:��Rga���`t����Ԋ�8��
#(M�����㘏�_���4�ܣ����-��[������'F�yxM�&�E���\+y������yPy���s�G���'F��f���7�Šs8 ��E�y�
蠫6Y���Y��0g��c�#LfS��%U�S���N>&CϮ�Q�I%mR*��?\�@��]�*+�ZQ`��	� ��~�2��� �]��AiO�S�>���xR9i����tW�51+�beT�,6�=4O+�\_��=Qe�(*E��+�3�jP�Nȗ�P�@�TU��zղθz�G0�j{~�����'��t�ŷJ�жe�Ŭ�hz��Lv����TJ�!�W�4j�_�ij]�n�<,0��;SQ9��3�\'?�?���ܪ�ԮZz/v]���j��в�ݲ%��)��v.k9`��F�!2n���Ϛ�,~�|�.=p�1�8�|�t_:�=�M�Y�$��!F>���X/�c+n3�G��2��$W��N��wW�����*��?&>�I}'�0zZw�k��<FG�@�m%�?�
�Hw��&z�C/�
�U��_�4�$pB!Ճ��x�+ϯ�գo���ƙh�`//Yxh����;�*��=%T�	;�Z~���w��(�}�ދWڢqnO�DڗLH�����;_;��2 �|����Nό~�m/����-39�Y�&l;�+���A*����n�ܝ�=X��(N��|�'��l���xu)�c]X���������Ҽa�=�l+	�(�ζ<9�2GC=��j}�Y��������VE1�e�j��R��������e�v��ό��]"Zk����ݏ1r�����s�h��������6WV3W�����(|3Շ�V�H��,�kcKk���=K�]!�AC[��3Fb����DTL����^)���f9ri=����
���:4Q%Tݍ�����$��ܱ��>^�����{�!!�8̾����񞽈��,o��t&}�a�o���Kj[E5@��z~w�E�o�O�8�ǫ��
`���={ٔB���H�}M��~ m�C���FY�
���ֹ�!��cS(g)I��`/�&_����$������Θ`�t���ll����u��Wk��Z>���˪� n�L�Oũ����`�a�;���1@�J_���sz5^����0������;e��`=�F>��_�q�	��y?�<��Ub�c𜨁�B�la�yy�����fl�k�oL�f:I�o�Nt�m:��@��&w=����5o=�SƘs��n�%�O��%?�M�[�8�~��I7�r�x��:z��I�Ȓ�駚+!:So��'��X/(Ev�d���tj[��x܃�6^�K�.��i�2�9 ���}g%T-�"�Z$T@�09X�P���
����4N�:~Tf�t��d��p�ؽ���Ex|̧�Z(����)<\{5a����:�G,�m��^�j"�k%�����2�Z�Y�����'>pg�o.d/o�n��ԒǗ=*V���2�r����i��*U.// �_�yҹX�y��� ��d[�kEy(���}�I��#c���A����0=�8�\���=A<=k�{�������� ������Skɿ=� ������}��}�Q�ុ覹G�7P��w��_��h@&A���)V{?�U.�(��ڡ��������*;K/��d�֔��n�K�5�MM��'�ȩ ]�����;�s���j��\��8ʘ�k�G6Jg���\ ~��Y�x��ݴyw�暓��8Q�>�k�d݁ 7H��KoS����1��U����D3��<!Q�ŕ��	�V�O�7�vⲷk���00mnw��{`��������Oj0(\����j�^�ҝ��ľB���('�:v�-ȹ��0$a��RZ9g��/��+�nfw�m�〒'i��L�����˷SBx�_��S��Nx2�<m�#ls�1�(�����@�z�I���L��xy��E�cb ��o���y�kFs���y!�c���+=?P7(���ƏL��� ){\��M��)�Q8�K�'�E��^=����* wz�iwh�^�GMI����CqD��-ԝ{-���L@����g'uH(��A�=�I�p�w�օ�g��=d8��p�$s�@p� 1<��kx��NI:a�Dp&9�d\�L�K�P�r�?�X��ꄯ�-��<e+�,�*�T�oK��$}Dabջ�^��H��g��O/5��O��O�W� ��!}�"�+���Ӯ%O	��m)���J����L��_r ��R��%xΓ{	��P}N�0��\���5Ή�Ry�������
�-ܵTlP{�%<�8�8��bJ��oƊ�7�����'K�q���x�,a��.J"�_5ʠ=s�t�^_��P�q�V���\ � si�sԉ,]ue�{���aVB������6���H��Ĭ��@���ވȔ�Ą8�ۑ����^(&(���c�����Z�$�ON���K�V==	�/��&qW��\]'�tz���Z>	26���&�͐��K孓�WmD��y��i3ia�Qu��ml�T���ɛmK��O���p>�[��"{��F�`H�F���ee�c�6�%d$�>qr9xe6���!.�[��r��?���A�`�C�	)��lf�����暣-�-�BޙN�s��F8�G��L@e�����]V�Ĭ(����H�}�j�(�Eas�t3�Z�!�yx]�Mp �.pЭ��{ԍQ�>٬h/�w�L���Y�7e�y�0�K�;��e�;&���F� ~8*ikL�$l�{����ߩ_e5G�/b�w-���X�E�E�-�!�.n^x�R�&\�u�U��N�8v�jN�5�WR�@G���sb���u��U^wa7�ӓ���!�f�ol����:�#�s���eiۦ]�[	�ht�u��d�}�l9Va>��L�y1"�ߠ��B!�3���R.��x?�5tX�5�h�۲*�	��EHR��]j�{����"�?���Z:|rW� ��Spy�Ο�C����k׃Ǎ��C8w2i�$L9���N�A�&�w@�C#��bu��MGP�U�e�q�DE�����Ƒ��H{�1B1HP�)Z������J�雯�WEHl�m�0d�ش���]#�U��ݘs\	��çwq��������[���ֿp�ԏ�I �n���1���Z<���&v�@|�ߦ\uV��+��8�еvjػ`�����p�A���-~���.��B�)�KA��0�4b4,�Yc�!�����
��u(���6���ق�e*��6aG����.���κL�%��� Ǣ��g_
_x����
��4P��V���1+�u����{m��|�٤?�\p|��\�Ȍ&��c��a}x�\���Ԡ����ɇ��p��x�rC�:t���p�b�+����\G_���߿�"�$���^�j��c,��v�j*:��^�Z�l����*�w���X��4%��9��{�1��M1�6�����J���Abk��E��$�S
WT��w����M�3I�"�@�7暞��kZ���d��*��P��S0�s����|N�'�K��ju1��X�Q��c�{}�XA�O��ͮ/r?��Qs�����M�"�:�sɳʑ��`��Oӛ���kZ�����l�y���T��Xcq-k丘o�E>0~�&�]�� )-�\��h�i� �ׅ��{����Ω|e�I���@z�1���o(��������,�n��Z^W����h���$��D��_�O�L{���mj1s/�Oh�Q��׷C&rap0��P�-n˴\�̬&��:�4:��{�C�E�	�+�m�E�&E�����i�D1�����%�K�9'�tS���َ#�כ3CC�͊"�m��X���󻩙V��4�ĸ��D��c�:��0؃��!��1��"�m]v35��7�ǾJ�W�@{ܪ��R�����bП��Ћ�چ�n�Y2-Q�~��-���5��7��a�gL�e����4k0K�������Z���R̊���l���PTZ�oF��������;���:T]^��eՋ�d��D.�l!����^��!��lҽ??� c���e�ui��̛���g�^�h�N[���i�3v�C`�H�,�#�ko�"�\0�-<�)Ar�o���<]#��\^����{�|�_�@p���24�xx7����uA�A�P��AX������j(�&� ���;�4���|�@@�B��G��]%b2D%P�����Jv��g�8��,>ڣ�X�[���XL)���φ=�K���G`�c��YN����k۸*ɲ�Tb�s�%��.湥oS
��P�(��Ӽ�2�-Q����h|��3f��Y#�n�oN�we�/f�3�wXx���.�+��\Jl��aA��� ����X�'�<y�[Y���Q+|���z �ˑ2i�!� �Q�0Kf�����ܶ���qE���:�3���7���'O4�y�m,|3b�գWk�:�讽E'/��	��OvSܕۘ��2��\~is~�%�W���s*�TU:��Z�L���m}���J���b֗����O5�T$�Irc�AYP���F!�z�iWz����!"TmU}C/�KR,Mu9��Dٔ�p�	�e?�K���T�\�A�����j�C,�ձ�%z,!ZY��d?�D/�>[�豐,yfM1{�����FN�
�yt3�Α=׿�g����O�����8�wg�؈fɰ#mO��nԡ���N3��~���j$��#��k_�A�]�����H��SP��͞3��:]�F:������M��ңJ��DB�;�!#*d5 Yb2V|�N��qR�ĩ�w�p�i��"Ӗ���n�9���.�o�<J6WVH*_�x2�n��~'���#�+oX+���4l�m�;�aa�Ƌ#��?���>�p���dt�'���r��G��z3�/�Z�>�P��M�qHYtW�fc+���i��T�t�a�R!�h�?��nm�)�n�`�@R1�����KM�=ˉs#�����~��K
{!'H�>Hjx�����K<*k�N�X��zL��ԁh=^���-�͛�x�$,�����(���"0!���r��I	K���G��Ҿ��,�&��-�y��;e���,}T��W�.Nx�x��:� DX�J�T��o���[�=�2�����y]�5�(#��Ɖ-ժ���]�X(g�R���3���ʸ�Ի�*��x=� ;��"��7�C���y���=�P���2����*�)IO��0o���������L�(3�P՛Eۙ���,=d���MgZ�`�*����W������F'�$\��S���yd�w�0������J��Q���ۜ��A�Z���}�
(5�W.��7�m8p�%���\���͌�&8��{���M��,E���9��-��]��J"�����v
�3��U�v��9�ʼ�hV���n��j����2s�  L'M�K܄9���:f"!++�6D�^H_}^��}�ݶr�P�v#�h�7����d��'Ȧt�g�c/����x�tR���>�QPk	J`��S��Yj�>'��&U���W���\$~l�,ګ�#&
���D�Σ�,*�[�ك(��#�6.,��Kt8�7�ēUdS hx[���'���q�sض��'��7��D"	N���A���65P��#��x��o%2��<��+�S.����jQz[	%L�k�̈�+�'M�2� }�\̙
�N�L1fh���ʂ���w�k�$��1��*�&7ֆ�rZ�\�!�W��o�Ei�0�/��_�o��^n'֒�hl��D� �x�m�l%�gz5�V���j׼R1���j�E�����%�=-Y�}�xa�վ/��.zG���>��.�����Ň�r{�~E@G�S[�	@;�7}�Z���Q�?GK=/#K v���J#{�Ľ����pz��ע�1��hq���N�jK9Ի�#��?*!�)yX�����S�A�������Y�?jۜ\G�J��	,��Ս���>@��;Jԯ��j0d��y[��������F�~7��w���Ü����Q�+m�
�ظ���A�pn��z�	/nKSI�1�����s^��p����e܈`*b,�6���:B��a��0��� H��@��S=�k�\v�qTHp;�,���b�����r��yD:o]E`�Vc�W� ��&��5�g|�xc�K�N���[_�U�7�-oݞ��6�p]$��܀3c|��b�C��'%�b�zb���D��CWI}&˭�ݓ�,[_?	F���؟
��7!�I�iRU�%��Ne�m8T�p��!�n�x�Y7��'�Qx˗yc0^V�V�[ՙF`�EO�GC^�^�ʑf��ҙ���s.bez�_S������Z��3�NsS�M���P7es�ҡ�)%_k���R�o>�Ԋ��|(���<	�
]�怓�k-���Z�{"ؗ�=��>�������P5^dś,u�Z�	2�/����'�{C�6��\֤��\�bm3�t��)�qL|K���}�352y4���{���+Dn�i�d��y�s�
�k�逩z�����S}f:������]m���%�����ԩC����^Ν�EаhAFX��L�6��x1�=S��Fu➺��0�5":"�m� �_F<�i�B����`SZ��๧-�7��^�|�͓b����:�fy3�QV*j�A�R7B��8��:IY�I��%d���|��BN ��iLT63�W����2�y
�mo����U���ޣ3���$0�o���	��&u��G��G��U`� �B���u��fr��֚޹��d��G��Bd��i�Te@�2D�n ���/�^�"S6������۽�dL�}{����j:I�=�b�M�Us��bT���{�M̬���@d����j�r	9WD9Τ*j�XZ<� �!���5M�<�$
��g7IG��y��-,4�e�7[k��=>��� ��_Ah���jj#���~^|�i7�Į�%bAg	dwf��.��f���ҞfRum-R�5��'w8�Jk2�����5W���X"+�b9��n��S�d���#�Xr�y�<�L���Y�E��F��l�!V���Y�A��;y��m���"
 ��b].��C�S���$��$d�E�Я���2�yE�|cЪ}���Fv��|q�jp [i�l�eC
`�rý:v�\x�R$Yc)���:�Y`(�����p'P-�B_��CY��ޫ��p�԰\db����O�]�V�E6�<o�o�x,݄z��l��	q�_�;4�z���ȕ�J��i̖T���_�s��C�E��h��O 񶓜�G��Y�"0��z�mҢ���|�,�٬�}7��B��_e��s�^IۈX/��}&0f�4�������3�Őd�>/�O9���K���OL�40	�4�^\[��5@�@�F^$�V�M}�j�F��qDV� �rH����6\�~�R/Eؖ��~kǇ�G9��п;�\�a�2�s[�蹦.I;�kU���K��S'�NS�e&q\�Uʹ��IN�!1"{|����(���;���o)��[%-���������7R~8��u7�>>�*����}��S��3y�gO٭=��N���j�yy�a�D��ݗ������f���oO�cM�<��]��� f�]��-~��U|uk��K���5s��;��%�C�����mjL�N�{�]Tp��`8��rp�r��JVl�B�-4�p&��1��~P(������}���ޟ{��:C�y��T��n0��@����f�����2>
�-�}(���>\T�+��
�)s!���7�LQ~�������6M���9�����#P�o��=��<m�l�֟�qu�u�Ŧ_,"�-�=T�l��J6-�	�N�Y9�?�&��f��i���ΙҐM�L^(e����ɜ�Xr�lF�@8����O��Ӣ3Ae�=s�S�b/�)�����J]l�K��IT7�1nb�A���jƣh�P�C!��t/Q�j�n�-p��nB9���tDG�~�����U�j1�8-	h2�j�R�t&��9���/}K� �lR6��l�ޥ�Wv�E�I�'�G���]�EN� 6��dI{��	�*^
3ov�A�D��1�=|����'~_	�_iY�;�h��
lN&Ӯ��$D�*_��?���k�N� �˫�|��BF:8c{�Q��S0z�,�1ضLc�s�Xj>�Kk�E�O9�mպ,��IXD���;w��EY��{��{�I�l�j+U��$]`Î}/�r��7��+'sQ���t�tU9��2
��4(@�������um�������+i8<n�nh�l+C\�4��̋jH@�ـ-j���~V!��9+� ��F��FWF���;��#��%H�:C�*[/!W_��&��oT�h⠳>e�q����3�7����T^aO��5
���lں��0�a+�4�T������!:m�+�x~1;K�m������`��H��^ER7�o��)�-��T?__��s=��δr*�b�J��_�����U�2����g4-������S�����Ŏ�l4~dd{��r�ٝ�Oy�b>Uo�]��w<�PtӤ��԰����d��QVIOsA����_k�u�w�؊��l���X�&%Ɠ������6O�:4	sdS�?�;�gXs�\��W��t|�n����\�H�Lۺ���f��֐��a��6���eoV�~�Q��H�#����$�O�����lQ��x/[$�u�g�YS�R�J��1��|��	�l��Ɣ|�;6�bp���s	r��& ��G=Js[�Q&�/���7~�:�JG�x�����é�ǡ�░�@���~Y������0H*�`���*�Z��T�r;��4�]F�m��#�m.Ү�lK�w�N����s��opDᒋܑ2��%���B|Q��ޏ��)��LB�`k��$��Z�B�9�q�*��z�󚗎Ͳв�ZS���#���ɉ�_4�lhRw]E-(qj���-���.OE��g.z��_an�EF
w�d����K?����df�^�G��`�V���"�si�n���L�Y~������!דgb� �I�����q��a�#����8p���-�5N
��K����q��!�J1�n��d>N�Aw���|_?����%@�w|Q����ެ�@U���W�E�-R���r�e�L�p���I|�H,i@2̿��c���ve��H�6�K^X�z�1Qg��9��E۹�	�?[���?-����'J�i2?�]�ˋP���M������F�Eꃾ���J����R��g�Ύ�$ �E��d<?�ż .�>�f}�1в_.̙����7�X��ų�����FHG�.�5O�K0p+�T�˲���)[}�vjz����'�oG�U;��	��(���Q�`4���uU׉�"W'�<��;T��&8�*p
�љf[Z]Dn����n�P��
2!�@u����;���&��]O��@��lu�Hg�N��vXW�-f��[(1��o1<�B�]�?��-��3t<l��ֆ��d����q���f�<�o�s�ꩰ|>�wԻ�Տ�B���縵&m�e]ͩ�W=�6-�`(U���D���׌��o�� c{�d�9m�f�L��⤧��v���6���5!��qZ���*:�N:�ʀ}� 졇ƨ+�.\hS�)����q�=?�A�M���@��@�MVYe�e7�B+f7�����|���\y���D�:ɿ�D��_��_���j�����%��Oxk��[����k����h`Vހ�����T�&�t/;Q��Y@�s$���X*ޤ.�1�J_���H|v��;�@����>�50h	e�3�"���a2W�� 5�BW����w'@'/�A)�f�Ь�`�TݖեݻV5�͝�q�0��K}�>vvT�@=)�Y��o*�N��]{O���?����&��`��,@Ď��@��c [
�E�bR7����k�>s��F�V�T0�w�`P�Ld���~�)�&�)�٣8X-�i A�
\�y�O6h�d��y��Ԑ�U�V0��c�]h}8UrҪ�Ol���5���W>V��` 5���3�SisJw��9��\��\��j��|"P����s���k���$)�IO��X=�g.��5tc��J��fn�v�筠*�ލ���c%C<�o�SL�ayu� �q��o!㌳�d*čŢ���@�~Z��k�� !�ɞ���(��k�aSZ_�����34��|����o]�h�z]$��)Jzm�W�${�Ncq���V>�ĝT ݹ��!�jj�#�p�0+�8��6q�o&����n�%^�[oO����RN��p��)x�0���C�B���i	5�v��ګD�+z�M�2���`�d���wlm�0�a_�G�_dQM۾P�������`g�	@ z&ԺŵԞ����,�<��"/X�j�<z��P��^��2?������i��E崸����y}��>��'�h��z�)n��O���/
|���NZDG�,b�lw��z52il�S�*������ƜeTY�0�Ht�V�a���n�xEe]qg#Ʉ~��� {Rl�c|����M
$;�.�9	�4����0��2 ����(AN��f�R?q���9��O�W�;���@�&����r�L�i,X�J!��	�V(r~8m����v��ai`=�,�qw�r=*GX��R)���9�a6D��ڕ�叅�0�������å�%���%!�o���t�w2A�|'U� V��p����E�Sf����9,$���Q*�²�"��B)�ae_駱����),���yɺ#/����"f��x�X#��&\��b��M�nݖO+8�_�o�
u�4�ws`n "���ٱ��F(V��Y4d{�B8}�1�DX1"�ߪF9���!'ֿ̉<���K�L�Es�K�U��"���m����o�B�RU����/B�n,��Ґ�Tԛ�n��ryC��>͑Tua_}����K�خ�Qࣾ�8o3?��#����=�O�ؾ��Q����Ս�XL���[)�b�c����UVo���@���'w1��r��<�A����px�I�9W,��8<Q�!g��o��_���!�#�lv��=Ke���h�՞����١�T�f��P�`:�@K��<���M�-�jQ�Dc��J=n���^S��5^8�	�܅��s�W)iA5� 9q�� ��.��/��E�8�)���DzѰ�*�r�ҿ7���bP��=�8;,�u�tVt����ΚE�
���MFP(4�q�<'�I���p�8D�l�z�Oz��jVi���n�F%�:#�b^":f(-FC�:��n��&��O� n����MD�����(o�q;=�*�(��R�š���M�?��Y;��8,(��P1���� �XW����P�_:���-[�7�^�a���K긩��tve j��Je"�E��뾱��rO���<�6tc��1�x!b#�qk�/�����`ȫ��G�����[8���|5�N�l�Jج�̕W�NͶ=�}��o@�F/>�%�z�����}�}�;�t����Q�B!��P� B�v��X��yf�~��݌A�*�:M̸3^����Y�(�Vl�I	'��LT�u�N߆����0�&}��b�����(��2��<&��e�b뷤^��Չl�	��
i�N�sт1[b�,OV-`�U�}�a� �Wa�(

#3?��	��q��MM����(��GW������o}"H<C�iшS3��ܪ(b��q{�h�J��庇W��t
�F�(������e�.��F)��i@/p�a�񮰻�������M��J1�V���I��E�Е��[Ƹ�`�e���o3m�|�4�-0n��ip��Z!��y�X�J�����LČ�j�7�ێ^�3m�m��G���3�A\�u���D�������~�929�����W���0�_MBBV�hc0 �_B�==�M;R��@��k�*P0��-n��`�0g����gY{�'vw��rM�X8�	�E�m/L�	�15FE9!@B�[���0"�!R�(#_�9���?�
|���PET"�R��L�����M���S�]|J�6��Κ	��ۇDmo_��z
(�?պ�jL�=��S�.
�sA�o���4_PdBlQ!����+�1�P\����sWi������F�{�9qB��%D�����wRsD$a6)�6ܗO#��!Q�3�|OH��-d�n���ĳ�"u�`����`�(�qA$����|�ٜ)]�Cf�%��E�:q�=�+ -Nֱ�~>{����b�8M�VC����+	����(�R��	���;������jDm�����ɭ/�|��u�Λפߣ4��*�2���J�����19u^;3�_��A���e5C	ʌB�n��B0ɿo )>��ӯĵ	z=A�H��J
1JD��`!��#�n�2��龸�e�e�N�i��LA�7���2�@,���"� �[��Ͻ�^~�r�r궞>���U�����>b�_�c�54U�%D�ϒ	�U�L4�E4�
���M=Ƚ��{Ag<m��۶yᓖ+֦^cƌ[-2c�M��o��>�|�'x�(�)>�t�y�
��j�6��]�c�@�;�(�EA
l��jT�%�Q;S�0P���������/ 戏 ���+�\Cb��� ����7��/G~1��L��`Cm-��=�\�2wR��1%N��F�Zm
3˧Iw�}��%
�i;٢���]��8������z�\<ps�I�l��)��n��7��Ѧ���,�y$�g?\�b�6m��ʢ?��o�0D����,�G0�p�?��@��0���U]��_��B�`���;	iK$s����������d�X�k�.db��N-E�=��Y�"��.�6��N�Y������gT(��椓^Ŋ��B��r�1��pr�K�t�9�v:��Q�Y���^�/+ʰ&�iǭ�p�b�j�C�'�x�h44=�.o�E��B��b~b
r���C���͝��p�oc�~u��$U���,�ɉ�|t�a�}��K�Ƌ��mm�SN:�@�B��1Q=#f�h��a���'	{��?�H27�7��ߊ�O 54�`�M�ꤟ�>�Og��vl�9��Ev�� AZUy�@-H�T�����(b˫Ul�l���k���
݈3��M��4���� �7��n�\�y÷L�-��#�x�%ě��NRbD'�ƀx{�ID��_�9�����'�l��\j�\��?�*?������_�D������M��J)�t�PsaB�A���d��F/�~�'�@3�@gR�d����<䆺��N����l�a��iF�Q/ʥ��d��ѩ��rɈiM��X��|W�'~)^Ei$:�!V�!Loc2t2��	���N����b��[�{�r	����P m�����N~B"��1��д��$\_kĊ���,W޹�х v��S.�rY����9=�Si���q��N�Ư��!�n,��HN�޼*�|�/7�ɆB�����z�����EOB$ڏ%��/���b������d2��+ٝ�8���x��)y:��n�#�|���B�ޱ@El���G�|��ޚ�Ո J�p·���[$9�G)ޠW���~T7?�[���<�Ӏ�l�ܾ�(�]}�ѵ�Z��^U��!D3�����Ȧ|'��"� I/뙢�󜼠o��C�#�w�:���3��ʋ�.l��V���6M��,FH��
��P�/�ǵ�bH�^���3��ٙ��3�K�%}{S��H�xe�8���F_D��elԍ��?��Ɍ���0 ��n}>'J�1��.���M�x�~/��#����8g�z%��gL;
�|:�wF ��0��e2��#Φ��Z����aU׀�xw^�

}��;e-�Wc:
������&���]��m>2Q;�<������P3�~) ������~7��ʹ�������X�{�4l�ݝ�0?]]*_�'��KmrC���?��y��C������̇�9Ȳs���cc���
f=9��������u�,^n8�FP�s@ �t�Lp���/��Op��zt)��f��Qh[���65�`�.��ې����@	�ә*��9p`�A��9#/<����s�9�!rԒVn���G>��V���v�E��S]��.����� diʽ�=��$�ٟ��ֶ�T�~���uR�ܨ���8�˼t!�v|��OI�&)�?�Tw
����0�mDa�,c���J�dk�T a	s5W���ɢ�ȥ���0՛>�]Ht*�5��5�)�/�Y�"|�t�s L������*�Jަ"P�.fBZR��<����"�0�>����,n3#%�~����DI/o�}C���Y825�n(�F/���x�{	�e�	��18N[s�FDa%������,��1�r9�������F���
_�_�V����e�S�%�{��+�F�"u%�A������,���b�1Jw^=H]��?�n����ĦB8�Ԇ#@�l@]~�Q ��kh>~ӛ���|��]���(c(���.��Ą�==�,��Tur+a��|mNV��~�ӡm�N�O�l�sF��Ĺ����:v��֫�C_���wJe�i��o{^[��p�w�F9u�m�����ȷe��*U �g^��DD̆��C�,=�(<o� �ri��g$'�3�3Be��!	���s������ȫ��.�=�7���4i�[F�F�9\����Y&<���#�1�M�5k�܄סV�1�����\[���;�"���eX�����S�Q���74�Ñx�u]vK��r��n�R����?��iJ%ݗ�ޞ�,g�2��apno�tV�_ʐA���9������W�]�0��>�ҡ�®n\(?`��me~l �@i��j8��E�*�5֏ũA~O���w�Pܮ���F��q�3�j8O�������h�:�R�6n���V��$׻Ki��}���W���U��t�Z�?�^�Vʆ��/��v�;F{��a� yRpՉ���\/�h�m�CnhS3�܇���{���r���|t�f�!�jhVl	q���g���h��@fh?����CN*�]��i�I����*� ��].w�J�>�A�� �����t��?����|��8�Fw*;���f�V�h��{x�n�s2�M�<c�ao�3�����/�HW _=0Կ���Y���I�20� ���	��I6��}�����޶�|��=U[$GN �HU�olg�,Y�dt��;c�N����j�JL�y��r8��I����_:r'!H���|~x4.a��,^��γ���s�P�3��<%?�z.��ĩ�(8~��kcA���~ߌ��9j��n�T�8WY��(l9O���'n⫖8������c2l.} �	w��74��Y��3���%�?�g��w�<9���'����5&�W��6�)��kd�n]g���[IC���)�UU�Q��HR�A-~�K�v�@��l�7@�lv^�0���~�@{�N��hY1~K��J�'�&Q1(zk{%�J�t�D~@7�%k��C�:l{�cSXM�����fR�xSPc�d���H�6��������=�u�!s���_��ҧ�p2V�E�V��Z^2��������IX��)+��]��
�d�Q<SH��?�O�}��lYU�����'�g+v  ������4��������J��E��3�ċ'���:��p|�8����TІ�}�n`�-#ņ9�/��� m��χ��ZJpˊA�.���S���J�2[Ī�c��O�����J�ݩ$�*k��%1��,%
�#� ��cd�|qww���t�!m��bϮx+���^0[	�>{���fR}�(���*�+��2�&�e�QJ�E>g2�ٟ�#��g���q-�H�pQ�C8נ��G�=����.�=��i5�t���Я�nM�Ge`�k_�������W��\�	�U��E;����}m�ώP�MK�Rй����
�;�$Tw�$6,��.2G˘-o]�.���Yj���S��h�9��)����x�y)���ż|H��z����>���eT=&�R�H�����R� C�G#,�t�%N+�y��cP��^	�6�s�<20�M6�g��������GS������`������9[��z�FK�gzHs�x� �5|/@k�%�a�m~
-�	)�z45sx����ȼ�S�w�P�#z�]?���p��Ģ�y-�*�ᢳGE�׳��K����`^Y3%����9/�R�qMZ��(b�>�p�o�1*�R���#�������ׇN!c� '��z~QJ����G�nd�`�����"�-y���B9U�y�gI#j�x�{	�ybp4��������=gfz��.JW9Ys�����M9�P;l��4Ap���?����
�qx=j�K��[l��Q�,��v�s�f�F{�5�EW��5̬H�֎���^o\�^jG�B�(YWACԖh�tٿ�T�*(���,���G��+��l1(V����Z�WM�&/�12QZm�R�˓qu\��(w֟�9�u|F�˝���Ҷ��/c&*������E��g�����zࢍ��vp��a�3 %�w��HF��%TĄ����_F"}���'�I��7Z5I���ԯY�j��X��:8vܪ^�³)_��t��������\>��J���ZZg?�c� .�V���]>�c�[�G��d�dvDbj`�z��[@�IT�'<�^U]�xz�������l]��=>��/I}�)[}f# tt