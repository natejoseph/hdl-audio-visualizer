��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�YO{��|+T����� ��9�jk>Q�5������3�+���Wv�X��u.�������|�[�}�QMvTB�űB�t+�%�B�����$�;�-Wŭ�L�R/�c��cu���jh�����Ѭ���_�<�@H{0��]iG,X����4S���$!�b1���B�ZE�i�\N�;6>@����j��L%�O����XVN ;���u�e{�P� R>�hi	��"��(cR�����R:�2-����4>A�8�(��g4w�� X�m�.C�_F��'��r�tu����F~�q���Pc|y��8�N�sȸ3%~7Υ�OwQQ&7_H�ĺn��ϩ�i�y˱<h�!��#/��;{{�pп�E�'���T#&��[(r@��.���I�az�L�a6�� �l�)�@ݥ=	k�F3!
`LD�S��aܷ�r�K��^�l%�J�����XE��G>��
�,LF�ִ~�>�p'����x�/��-���7���~?B��l^^��l���$�\B������P'6*l��:��JL�3�W����wa�I��w��0k�+�dp+���1i���3GK�{X�V�;s;�@�Xry^Z�P���;`5M;���h��+G^ᜦ���G(�H���Í�n�0�:5|��7��M?\�w(okd��݌E���i:���n������e7��$r]��Yui?��lC�`�Ys<�+D�?�&6�X@��N�Ϥ[<�ӛ��F��љ����E����a���ܛ�0�ڿCߍ���O�%I���c=����*yL$ţ4d~7�.w������x
n~0t�<B;� f����r3d�qy]����TT���3�H�j����J>��ӹu��t:���ۤ�M�)M�n�3�E�$�u��M?ʸ���C���D�-�����/W�b��U����/�`y�S�&�/o��t�o(��1QHC��}�̭��pNHr2��*��5&�
�ぞƬ	i�����;��`j�w�ko�s��bH2�2��'dS��C�0�E���,��@����������<�X��?
���m%�Ϫq��44TF����o_�t\�J�Ԃ�iܯ��VK�N�KE�	�-�+e]�䡅ڽ�k
V޸�nNg��¬:���f��d�{�|b��A+�"�4�dzJe�S�H�a�7�O^���E�5u%�=�Aqk��A�(k�)ʸa]�-sa{��k�vQ1�4R;#��5��	"اrJ�X�kl�z�/"?ǳ-p���*�(>�K� ��P ���]Ls��ӯ���I�ϋc�ޒy�.:�
rҥ��˚9���IQ2� �۬<S� G�I��x7�ql.����!Wݟ���[O�+e�g��������~D�I�n����n{}��O��-�ە���N�B����"9�9�;���(�ܘX�@n�ٷ~P��0M碢<�2ֺ}�]x�A���C@`��8�"�a!��K3<hr�T�f�y��h|T���2���N�W^p�Ǉ��
��T����x�q:��d@Q"�˫�?�ZE�4�?���ٌZ�ݴs�\�p�6(�5�uJ4gX%V�(�+���2ű&��j	��o#rX�FZU���]!�����BTSF�sD"��Տ����fqds����1��U�C�oS��D���s�JL��;IР������u��GYk��
���9g����⚡Z8�l��c�o��ƙ$�U,#�5��p����dU;�Ҩ�ؚ�~������A`Õ�2��-�QL�l�,�B�Ta�@���.[�� @�������w��$z���\Ě�iKn��+�r편~9ī�}�ݮ��u&�ꠣd�pSP[�4�KS��t؝i��2�L�6�LV|~����!�G�Q�3a,9VJ����9�!�d��)�Ru~͈�y�ϒ+��v6��4��f��&��	���z��/����N���o�]��I�F���H/�#�"��J��� ɻM63{o���R��A��$0I�'Cӭ�!�����r ����o����9�Sv��5��	D��3r��r��v�� H���\S@�u���L�L�^�\qD]��EܻbB@8Zxi7	]C���,�����F�Td(�ݾ^��Xv�A#ȵ�3k$���_*0�b�
 ���o�.�`�k��H�^�t�#	Q)��N�(�u�o�Q�0.Ɏ3On��C�V~�0������;�Em�e�.*����{�Ś�l�/C%����2�FY�i�N�����7q�q�"�܉�-�j98�q*TFS�1\��$�@I�3�k���t���7��xn�����"�Ø�A ,o`4�Лܒ�P��Y��T]_q��㮶�k�@�C}�|������t���e)}����k�鈚$�%�X��l�`�Y�!&��j�`�1ɪ��j`:-aݕSԺqB<%nw|��]\�b����/�=�`�Ld
i�.��.i��S��IFRи�������GL��Q��+�>��2��F
����<�~�x"�E��b��J7��J��]�Q��A�W�����}���)4f��>S>/R��$�a=P�����ڎ���f�MCz�a{��.�U�Zz��a��A%�U'M�'��,��h�n�ԯ6�H)���!Y����R܊М}ߗ�De�����=��Dм���b�T�י��/F���ǒ���<�[�ޭ��a�.FH�R$���Ԡ��B���(3����p+Kf�w����O&*�TD�����i��ŀ���]�����;W�Vـ���	:�¼��D�W G��q�`i��|(I�P$�Kf�=c�)}<��K�XX���n��G����T9�z�շ�����pɆ���šB�|��s��c%�o}Q�S,fMb�����Q���j�!xb�,�1�������o���;~�'F�x/�:ȷ�K��K[�s�k��<��n�����q���a
q
rla�h�9������Q�lN�R}�*w��_H�(�VjL༙�W|[1��n���1�d�� �d�_��򺦥h�_�#�������צ�aV�R_D���7[�̌��qS��5J��͂<�iEɪiP��&��ҏy�,��D7g�Qj(�U�tZ}iC��ɝdE��U�ݝ�h��(��]��n���q� A���̗�(����1n��Fk��Jet��)�5R�C��]���An�S����e��02�at�Olw� ���A��+ƺgP����$��)b�Ԛ>*���8�9�dg�mC@f��z�ҘgX���Uv��f�@z(�tӃ��wM�_��0�b�����+��P���2u9��D�| 
��D�G�C������O�+�R^�S2-�{���$)�ʙ�Uy��>FƲ��֛?��	��ā�� d�>=R�O�B��;��~����]�����8��3�"�����|�}��׼1y�Y�x#��k�����f=8�ݩl#�Q�}�^1�hN���᧤Z�O�Ƞ����P�g��ףp=����Ûi�1]�jk�IGv!Ў9S{�9A��>y:�o��Z����$̟���2)T�	����%䵑7��!5��ϟ�?��HO�K[�'��8)vw��a�X��N;ߡ'iE-�{�"�4���ۗ�LTeY�*�Z�'�Cj1�R�����|r;�D����b�|?������SnH~�_�����g�C�r[>M)���ZV�F6�J�#��J�6#�����.���O�(��,9���b�<�j�)�܎H��Z1�Ur���qy���Z?-#���_:��O^}����"�$�z�r9���w��3m����\M����TH:\o�m�x�|���՗�:Ɍd��'��ia<@�PGøfL��ec(֙���Yy�~
���i��/����/��^f.ӆHF(�h>�ؓ�:���v9� ߉Bws��ߣ!�r��9�P|!�Jn�9ov�$��J��.� tw�(��..l��'����V���a��'�='hP�?�p%l�O(���P!I|ݿ�U!�#�cT���"q̉6n3{��lvmܘ��9�+��2�����"Θ�=q�2�"���crM�>�:��>��P�)����u^�=W%iI�"�>@SwK�{�Ԟ�)��[!_��i��-�Mr����>l$