��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O��"涏K}�?u��+q�<�j̫2�A͢l�Bt|���~�0�:d��L�0	�I��w���u.���M�jh�$�`�lՒ|A�Y����<���=odI{�^#�F+��H�[Ku�4�L;[������	��V��#_�����a&��'���-�+�%��~/_��@��)��L��'SG:Ҹ{8�"ݟ��u�]��4iB��8����X�S�{��-�ɔV����\���E�4/�n�{��v^2=H;���F�����B,- �۰i�Ѣ�-�"��Y���(?��㘾�5���l8�%h����v³��J[Л�E�2����UFDC1~�rO���n'��f�VyP!}m���BݑtV/P�e�uz��s�xm�&��aaPBb淃w97C�D�H�i��D�n��֢�d5��t�����=��'���W�=��x��5�����(��Cza��*4��y��K܆��� ?BpG,�]�@\*��~��{�Q'�#�PVE��c��k�v�"�[l` t��fU{J�����SUi�&�t���b���,��ZTzx?�5��,��\0�KR@�'|�/zptd[�����~7��|�~�K�i�W�ƥ�&�8#�o<�����R�&�p�(�\��xp�t�钴+s���5K���}�Kq��Q%�[�$�^���k|Mg�*\s�����4��qoM{|����u@v���P�fg]|�cuSj�;ی�Z<qe�`�nCn�?��bU,�HM%b�
,���|d�F�N�e�rAu��T���5�Fa�n��^�rY�%d�˲@UO�KÂ�/�W3���.�Y��������#�м���lS�%��$֛ z�7�Ua�6.�~�J=�ݣ��m	��6Fܢ�/33��<�Nm�E_*���s�
�6�J�������lc�Qk )_�L[:������Q�Zb"�vy�孑(���L��=��e�̎��j��?���|���ư���"b�7��}�t�ۖQߧD���ΰ�n��yYax*��`4�L�t��/�'��F~:Hv9XӉn���a�1�Ɇ�e��t�9Qq�T�T#�}Lqh���d��ğm��ϩ*� AU!U�@<����K�M�F�j�>�abnYҗiV���AR�$�u�d���Bb� V����ض}d���`lږ[�6(�w�N8���KK��),2��a�A3����k.U��J��+h�W�{����;[��;���l���Y�{�|L�6�4����[C�܊x�?�
�k^�\���ku-h	'Tոn�APbH)"D����Y�5��ܩ��ݭ��5�+�ҷ�ӣ����m���O�[��ڔEx�ZF�Q�·�~;z�άpw"�_�v��-�Xf$;*�Z�bA&����^$�;!���I�<AO�I��|����t}ې�9,޿�4&�tq��ⲋ�rrH���ջx��2�=W)�Fa���ܭ*��V2>�z�8��!{�j\��v���v��7���qB^^���$iݳ>wl�.U,��u�W�=rԒZx�	� ����d��,'�`��s���,��m��Mݗ�{�/+�>�Ւk*Tr���ׅ�8�$x�S��>�4;�oM���ך*����I����2��/9���F���H�8���U߫Hh�P����C6�!�=���߽E�����b�H�u�n���?�zs�&��\���U�b%V�.�W~r��mm{6u\��k��^Rq2\8n�R�{�3�V/	 ��C�"C	c~=�m�׉w����8���/��-������i\�ҿ� �[)��R/;dI%j�!yG�l��Q\���GF�"<ì[���uZYY)�-�v��7�?F�1�n<�x�	*B�$�CD��4�F?7�8�C���
�u�%Pv���������
��m,*d��e�	�ǩZE�dl�0騇
�X� �V6��SmA��QtA�g�e9�T�U]�L`�I �������|���BS!~�dO `[������ �E�*�=y�dC�m}��(�w)(��$"T��Ge�	��M�v�!J/q�ik�s�O��Ť �ݔ�U�3��da����y�>uZ �1��NP�~�����Z����2+l�S����j��⩁Y��2
lLM�5ϥ-�%!���$e/B)���X��{!%\Y��0����k�qZ�n�ɇJl�2�ަ�N�{�{��|v�O�&���=��Q������H�I�CL�7|�F��5��hJ-l���[��^¶K��\��7�e�1Y�#<��%�>|��d�V#�9����tS��'�u2
,�ykia:���b��E徲x�L�[7<�� �B�k�s=���N��PD�`@'5�<V�cĂy�������d׺f+[������A_ׇ�E�a��iۃ����'������K����C�� �}Q���ޕ�ܶ`�]�m������,�������)���oU��60\�'y���A��TI���No.@Cf{�J2�U����`�q��CH��$��,�򳯯x�M$a��K�Qw��V�K3^XM��Ľ��,������@�}�8�Li~�p�xl~PM�^[��H�<N~��'��e#w�^}��I~��p�����-9��Ef�z�����w�>�l:_�k����O�������B��h T[�I�!�I�٪�Չz�%�+<��x�c`
o���8>;�+}4
.�:r�c�}��m�&��:�xK��B�Ĵߨ}����+
���I�GZ`���9"Rإ��Y��'���$���6�~�X��fp�ަ��.��;K$s�a�C��WX�)���.���	���TB)83�G^����]f���"��`b�k�)�%Ă �ݍ����0q�+��|�����ay/��	���̨0Daݐ�����L^�utUX@D�|�V�/�p@��� ƾ��G��z�/�0C2����?�ͼrn;����'�3�4l��׏v�	bϹ�n{�{|"ZGRW���i�x��Se�5B�'�WD��>U	$�j� ^��K�����[,!�tLr���K[JĘ���C���/�4V�M�<��4������Ƥh�]@�$�l�j�I�*n�1�V�B'm�{��X�ic��;��0 1U�q�Ax͑�8�cbi������J��0���`��<Ւ�7�	����;+'�9��������B��V�Y�'��t�Vul���ߠZ��q�$�����j�{��l�M�,B\�6G^0�'�gd}#x��M�7�Rh9�����v[����o�Q�C7��πlU��z�U�F�o[i��V1QC�ɔ�� �a�؏-�9|A[\�*Y���&�����O	�
�m��e���a\b.�9G���J]�n�"�g�Ue�"��'���f�(��0���>.2
�A�m�H��6��C~n����C�1��S��A����.PW�9��=Ԡ�#z��x+`G)V��|V��
v�pV졶���^{&-o ��糍�O��p�E㌆�1Ï`1�u�~_���{2=&���;��U7|�}�M���p������X��V�����_�D�V��"!�a?�(��<�e��z���^c#1Iq�zV�J��].�x���D휷�M�yPu��ԡ�&F&�6�`�=�2:����@켻��[!	&� �z����!�s����]�˞�  / WXP,6
�A,��!�K�r�lF����+���u��|�Wg�5�_��jz��R�s�:��	/������10��n\D{��m�f?���y6<ĊtL��]:�C�/n����R��Vb(D~����*�J�㰑�<I�4L�NJȣ>6|I:A!��h��qV9K������_�CZ8�>lACcS����C ��r����o����X��>~ٴ�<7Z��搤�c����|jn
�i�J*�$���q�`x�{�u�����/�a���P#Bi�Jz�	�X��I�	�1�6H-÷@�_�pxFD�,jj��H|�E{ʔ6��:��e�#�.O��Rӈ��������1eZ�Ut�^y9!��(�ɜ�HzHQ����0뛐���������^�����9�	о6�j.�&��U�yD4����͗I��s�_w;����Lmz����_�<�>w-�DC5^=38?��vF��x��t�S��٣����Z,�Y���k�B��6X��~��0�7���({=����14y�2V/vzpɹ�� ��;\�i�[侺q�����^+��q��2d�B�� �G�g����1/^�I̹&7`9�&_��l����`o�"�{�������1 ��Iic��qi�jX�7�n��'���/6��W#Z�wB3�r6.)���g��[m��I��K�'	 ���~?�Qt����`.�ל���i`[ɢ����TW�� ���K�y)�6Ț�z塩e���|��f-�AjT���jC�sZ0����9�p�Ma�rl�r �����e��V���}��G:�T�� �.|��͵�zy��(¿W�Nt
���~v6<v�Tj��3���a@!�Ԃ�$�g<�{~i'�g�b�
�>1Efx���.1�6�9�V#�c�
�4�"��e5I������K������E��HːQ�����8���A.p��W�W~�ɠ�P�r5L�`�|¥�L�S�p�@�ߺB�{��\Tkni�S0Y��a��e�R���&7����Z��/B�wp��o��j�줌�,��l�_��ۣn���m��hoҁ��l�*}����3�q����ew.=�	�ӏޖ"��)ȏ��(P=�/�jc`�{	�K���-GH�z�F��⩶2*	c�/WQ�` 0�,Wo���x>G�4�¬�B�+<���
ҝ
���܈�ݵ;&l�c=��6�/�t��f^+%_��FW)��&bO.hӰƧ@q��|q@:u�����m&e �����˲�ۖ-�d��,�^'{�~}Ȕ~�ue7@e�^sc��c0й>�6I�J���=ּ4X��?��{�_ѹ��3�e#�������v^ Z�.oJ�D'�W����XוyԸ]S���L_��]�逆�Q,%�
���-Z"�#�k����l�i���*�'��11y�i��T�p���$\� ��*��4fҔdD��3����ݎ��C0���sg��}�"�����ޠ������I�	,q!����pP��/(�#�~��{�j��;s@=5�
`^kd��[p��7�p�r�JӺ�U|Eb����bV��d�1�`	�'��Z\����1���A�}��ә{��i����0�f�D��,&XS_\�U��Ȏ����/��g�����\�u�U��V�cݛ}��S-��N���8�/R�e΍\%E�
�Y� sM�z�Cf��t��^�Qhʋ�R`���'vůǗ���JN�2�4��cl�Un8������> ,t_Blc]T,�K��
n�R�����W���S[�:�� v�1�*����R�[�5I��-��ty3-�{�0~N�ݜ$4�y=�Oi��V���J�?9[��Q5����.�̳0`Vl��
^:�	�@�~����^���;\�Z������/�p}y���[�޾'��)L2�&5�%鐓3SS!R����O����F�[�!~EHJ�[z�P����H��nݬ��z�@�$a��2rw����a��2��l8tOs�7Ka���li$�YԿ/�4�Դt�\�^@�a�y�Ʀ��Zbm�,{��B��6� ���:2���,#t��;�{iPM7�j��T�L;.�ح����!M�ɦ:��Lj4h�Y�PjE��ʏUd��jq5:��h����O'e�L' Jh\F%�����,���O5�r� ��ŵs�5�L�Q^2�#�t+�2�.pD�2�ar�8l�e�� �z�5�i#���J�Y��BFj��?�c�jx�Kr�I��x�#��V�"M,�d@�o���}�#��%�ب�&�IB�^a������v!������%����"]��������N�.c��&���kl�k��lx���Jg"���Ɲن��l 2�~�6�*H��¶+�Q/I��.���
:�dw1e�[�7I�$sg^�g,����Xn#I��q�?OE:���Hi�E�����>���x_Z�jʾE��s:�KۇW�n������Ł>=ݰ ���*@��x��&�����'�:�7��a^$�9�O950����M�j+CS ���:�"��!�E0m�)-�����j�)�b=Nv�!�lm����qp��IkU��6)D���� �PA�[D�cS!��`�M��g��v�N�}�G��YD�]bHȜ�~��� ���=;mr��.� Υߟ��fq�S�ay2z3�Gn}¤sjY��S}8'��ˎ-�_��&A=1�M"P�7LK���NN���@���X
ҹ�F������q5�l�������Ș1�&���eQ�����x��sdq�.��ˠ��}5N�Bő��B��k.�x�����E�ͭh/���	�Q�B��gyى�1�z�ķ��ш�)�X�f:�N�C����O�q0��K@��fYBu�OĽx�
	�VX��3Ǟ\���l%��w��B��b
�g�f�,�f��[?|��]T���5ج[�c�g6y?"���Ƣ�VKg�a��lk^p���\�gֶG#���]����ADm�K����rh��&<=1�Բ_/�.)��u<�.�����4�{�󐷝9��Kt�Ⴠ����ږB�>`����/����u���$z�I!��뾯�i��6VH�b,%��L���j%5��X�;����g�0kȽ�o
��Q��#e�4+���\<P۬K߅p�IY�