
module pqs (
	pll_0_refclk_clk,
	pll_0_reset_reset,
	pll_0_outclk0_clk);	

	input		pll_0_refclk_clk;
	input		pll_0_reset_reset;
	output		pll_0_outclk0_clk;
endmodule
