��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g���`�SF�Z�6v����(E�ݻ��<���� �1��4Ee4>
*9�g�Y�� ��3�I���mw`��ڸc~;V�!<���F|�Q�o�;�1�Ϝ��'۰�8n^aU��q�� K�y��l��㱫ry�B��x�!v�h�;��&!%�x�b&����_��P�,����A_2�	\W墺&�+�Z�t&q�T����!��a4|_	']^"�d�ys�d��[�k����ڦfwG�Pւ�$��%tCc�� VSq��g�����c�� k��y>�D|�#/�L+E%�*x���������B��H̼ú���Q
HO[����z������`��K�O8˖���3�ش6��Y��6>_�e�U$�0Im�4�����Ц��!۟Ed��,�V�`�"��R����I��	������\�~�o�Z
,����V���&�l^v+���DO�1G4cO��(���x����$?i�|2,a�[�a��L�
J�]��ݼ0�J��t)���GG��j;3�(�?��
'�P�i�Iɤ�S�����&����J;)k�DF�FQ/���,�6��[�����U]��`g4��1����L)�\�cػj�ARP�y����W��������AJ�>H��عϻ�Z�,Ӑ�M>�\,���O�7�>>�JM/SV�~�>�s��q��P����FV�J�cv��Y����iȲ�Ĉ��{he����t�N���k�����fȸ��c�
F����4��j�E����t�k,ۉ`]�&+4$��|���~ƖG�����G�Er	YT�*�|E��c�2ԁ޵��c�S��	 BI��ߞ]��O�:�S�̊�řA/($*^���n;z&�K���e:�d�M�]p��t-�ui��ĉn47P��=���8=�v��a�* ���Y�Y���1G�(���+���$cT{H@���%.)� 38vc�(��/�Jh�b�I�0͊k���&>��o���D��ȉ����syY���|i�AHm6}��Fð�^\�0��&��`�KRܫyՁa��~�\��S"�y�$a�a���8\���NAۼ��b�6�⻛���%�p��P�m��m5����G� �&1��D� �j��X�g��� �S�I������W9���:a�Nň���omU��K�(��A&�wjg$!,�כ[[�J��"�른ҁT}n$J�e��N�$~'Z���64=3L$��#���#
	�M����5X�d�=�3��'b���b��t�D�{��oͰQ�?��7��Dp��n�(-|�?c(�}���
�Al�p��#a��Y�-�U�O@VC��T�7���G����f�"/"�G<�m���@Gb�&��v�k��`�x.�$%%M-F��!h�.��{������<������ 纣���>O�����Z�yk���W���a[k�x����[�@�!�Mڌ��[Io����H�rm��c�kN9i9�hA�Ą�fu�c��H:1���.��o�܂��y-��?��N���\
�9�����pQ�ɠ �����oPh_U�/�@_]�Z���Έu173L�H�p�cb�k�`���ho����7���3VG��: cs��?Ӡ�2&l��r��Y"}+9�W���L����BOަ�6���G��
$C:s�"A�^V�~GU�(KV�4ʟF�����|"��N�R}5M���׉�6SG> Ɨju�ņ���y�*Bc��Y�90�+�3��J����0�-�C1��ǪX7w`hT�!����'ޓ�!�O�\_���[q���mP0e?AI�Y�F$#kH�irL�zqZ�����s�v��Հ����>4�tStN�gq�W��4�s��y���=�u�
�ܞv�Z��54��{FP��_@p�(C$�2BdD�I����E�o��.�Y�ch/��ݞjxa�~۽s҃D�g��gZ�R�g>�Dj��)_<����:�4ա=��:��#����r�MQ�O����f�h�/����S��-7��H�ƍr�@=��?E�p	������;/���Jh,��\Kp�q��\���0��Hsq� �幻��	;��8V9��5�S�����YzxN�T-"�����6�������7����lY�mN���`��R�����p�����m��.�y��*���Y:#\� �*�ߟ�x��n�S3���)�W�:����#�%fo�ZT!�� ���1�X�����8��Tc� D�9�:_�4Ɠ�-��	v���{��y���f-�b�gO�2�5�3���|�� P�2�.րdJ\��@%ċ���a��7�/x��N��a/��o�"�4�.Z?�}�f���d0X[�.%���<�%�2��&���x��Rc� "�n�ǱQ�T��.�T7�Z��3\C=g�X���.�����C��!������Yf;�U���F��Q' ιa#Wѵ�Mr7�����ܣ&DO[�2؍^��k�V
W_�	��'7c"bݎ�� �9J=t�#Zb�妹��V�\�
7HS	.+���u�B";�5C���Ee{��g���_�l�Y�a�UU5!�c&:98�m�g]����s���D��m��(�<��)֮���58��2�3��NΈq����w7C`{E?����;.F�G%N���t�;��
�aEܸƆ�$�N�L���E���敷�����è �ā�,܂�Ꮅ`;ܒ�6k��WJ������e� I�j�	X�+=>�
�w��M"�^CQ�3�{���E���y��J5����g{���i�쇧�?#D�G.��'���^x�"�nߤ�v�������W��Q\�pX�rt��aS}�Ja�#���X(k����L�P%���{%'�a��}mg]A�m�h]3�>�!���#��O�q��|M���a��=$�����,I¨d�J��ы9"=�0��/u���oV8=#"�o�@���b�_N�u%�x1_1�e}�xm�zD����u,zR�6�N���#�i�b��'�5�� 
��YU�5Uv�_��86�N�(7�K:@ƁL,�޽sL*�����>�d%�g0���{/�JC)�9��3��O!%.��7ԙ�v�v*�k��=lV�$�Z(�6S��N1��ug�r��:sօ*"�:�]h��6�O�2�rF ��l{������)T���T�����]�N�E܆A���|?����֒}?�"��	G��8pX��ll$�&kf��i툩>�H��oI����Kv�0B?+�OX�u:ĩ;�������/�<�����SW!갋�0A��pp�to��ˍ:f�|}��4e�)
'fY�9u���x\A��T �魤d.�,��j"��ozx>�]��}�UD-Ca�Dכ��ݴ�_�JG���t�� ڦ<�nbt�z`�υږ�v`��*v����Q�;��d�ޗ�g�}K�q�A�-\DQnOi����\�qN��U	�Z	���]���rGu��^PF=a'�e��S�G�r>�t���X���4�!\�cđ���a9dsցα �?o.i¯�T�}�a6Y�O���_��������^�'��J����!`�Wk���ѝ�$���j�3�iT���ל��"%̸t��ǥ¸F� N�5���=!���P��VR��CQ�]o���/�*˷�C �WM�k:�o�2�m����2���J:lf��=ͷ�o/Mc,{�9*���?�ض���h��w�h.5���q6��a*(5���t;�;�[���Q&�m�o� >m9���H�Y˴��)��J�^[��2Ôl�H�0��F��m���&���k�����D�l6�1V�`|�tؐ�Ir�\�l7�H�G�)��S#(��X#��T��8�}�N	ҥ�x:6�6�N�}ZK!.>׽حA+��R�z�x���`N�qVV"��MՎ�E��q���niܻ��T��x]��_$���ѦvH�]XKM۾M��Y%GD�U�議Zf�����F��e�*�t@fWTY)�'*^�� ?�CU�����v�l��Rmic!�6��&U�wn:<��߾c��"Q�ሩRb��ma��x�6.𚇿=�ˣq.Z��T�����ݫ]sy�����G^E�S@�Ρ+*Hr��&O������p^;�헓fd��8�W��Q�S$�*��b+J�g�~:tJ����|.|FSH�?��׬��)�U �����ܢcM����U��Y �Lъ=ޞ�/�$�+mx./Y�&/M=��C϶���gV�LQtO:�S.��$W���v���7��s��:����m����%�7�J�d���+B�mjW�;���:n��.U�����[�p����6<���揱�G�wC�)��`x���!�o���N��I�D��پ塒ُC��F���ОWc�_����I�,�ŵ�fW�@�yf�K�0x#�q��
����i�X/f;�,	g���iչ~Ǚ�s+��{�v�z�v�9"!�>���q��:�D[�Yv����CB(�LU���OC\}�H��2��5�ݻ��1K�=6��%)Mn�Ͽ@��0{*Ǽ%�t�7JFU��oc	5"d��Ǯn#�2Da���r�G#E��_p���.�v�C��J9���d7r3/�sY�U�V8T&i��A������_^�7N�Yந�OU��kh����;����ߗ,�/E�M�F�|s�o����kF�|K��6s���;��y�۱:�3���G^6��Y����ØEٔ��@eɖ����1,��[�X��m�VƋ&7�/Z�ɧߖ	igz6Y�^�����,�������� ���KT�J0פ���j݅뺜�@#}�r� ��:Z�-o*p���_�����Ma��A1�@K@,��	>�c�T�̯1�� Ȓ̂lW�b���:�G��w�E���p��� j���@�:�
��{�B����������t��1/���$f&*������v��#���Nfq(e,��`���s����5�	0�.�o�D��1I$ܝgX�ʑ��z��Զ���Y]4'��buv�X�f�-#tL`~�v
# ��2;����^�	?�O��%���{�����N� ���W��$�FMv�c���g{Q�5��Ϯ�����:$��	�b� �d�R
�J�[a��v�H�z�ڤbA* J<��f�h�I�I�1�(ͧG;�i��`��#ӊ�5T�{P�Zq"��n�w��|�"؇�d9/�k$fEh qcq��-h��W�+�]-�)G���*�<,^�$U�g��[����.�HᥚX�ƍ�=9����}��y�	1H7�*�mm�-�+���Y5����H�+�F�CE0�A� ~VA���<
Y��e
bN`O5=���j����;�(
�q��\m�mk�Ҟ�×d4��g�nIC@}���6^+���ԋ)@%���`�C^Ex*aP�Pge�e�#H4�:
B����+q��q�i��A�R�=�lBߊ��+ґ3 P��'2���x�(`��p�MXy?.���V�G}φ�o�G�>i���$'�A�F�3��#�*��1w_�}oS���+crΡ�e����K��((sPB!`��U�e��z���li{�N�n��@�N=tE�"�O�'�3M��MFx�������R^���u�����-"Ń��C�g��}L�����ȉ�,��J��2B��x�h�.]�����%<G�A��$:,l5��K}pt�n��!������YX3�a'HP�5f:���*�vw�������x����TgP�|��� �kK�9O<��`'O$�M�Sc`KU�_� ;��� �4�(
�<����S�Q҆e,�f���U`uX�����d��j$��׮#[Q!�e����X��7�Zp+�
��.�NxS�&�k�{�u��#44���?J�_�6���{��H������N������:��G��T���$����I�9��J��|>�f�/g�W�;ç/ID��ǽ搷Ĩ�a�g��h
��4�㉯����H,�,� ø��f��u�R
T��\�i�鱎����nP&��]v��x�M��!�
�/봄����b�h���46Y0?2��5�7ۡN�$�H=RM�1㕟��j���#J��7j{��v�%��r���DV���|�)���x�A
8Hw;^�)+�����!ܟoN���W
�&�ሚt�_��E��Ow8�g뗷Cʊ��V;J����=zvNd�/,꙽A%JT H$�`��r �﫦�����؟��h2$ޕ�Y�!|nί%9���~*6�T�=36��s��sPD��Cs(h��##b�h��N��(_+�'L�^.""3�?%f
,n9rdT��x�i�e4�x�L�t�����ë����!`�����gz���I#KT�=ݪq\�N_XDH�6�����D��SM��ً#gv�s7m-pu�v�D�(9���K� �����C�p1L�'R�I����&���>�6qY�^`B99:�,ǅv�g��V��/B'Hs[�ћ�}�r��nE��L��[�QS3�Z(�l�F��|����HR��E�� �=����S����:(%���Iȶ�4u3�yv����xr$�d	k\֢��xnh�I���9��Õ�`�;ӯ��ڲ��T8W�VN]��y�zD?�ɩ�KBy�\`q�
�(*�����'�:ٴ�cqL�����^,2(�4��%���bFh'�F��mq�S$q��D�\[�4+�ʣ,��t�����"j���)#M����:��Y�1K+�w�4iq�%��������h?eW����F8"��[S(:���[�����VB����B��������_,J"rBɈ��%l5�=�Z���T���<�+
�ho��=W[_%��M��E���e����bT���E�~iwL|��v�
�D�a�O4�"!���Jb�S���1j�^�#tQPD��	IK@�"��$m��3���x�n��)���լ�Z�l�c0�Y�*4YZ8���n\>�&nf�_�Ҭ5�i�?,H��-����AS��h�{l�����&w&Qg�y�G;Z^R�vA��\��%��P���)}����9DQ���?&�� �!P#9,��9_���Ʉ�H�n�{�?�����ݧ�4�S�"�h.�7 JoO��g���>�ĵ=��E��_ߺ`/8���?����;doI_��	�� {��zxZ�Y�r��h��74ｻ_����R�xN&R�_=">b�Χ���w��+�w E��T�֙�!���B�"^������o�YZ��r���lpZ�����y��;�TE��I	9���޵��$����Jx�! ���R/N����ŅF��w��*�l|�$������֓�v���hu$6�;x�%v��5;��� �TW�'gSC�K�a�<f�	�q$�Q�	;Cp y�b����H����3�6���� \%u�eYꩩ$ao�P�����3c�����wd���ԩ}?��Sa�xq�Fu�K�:=YsEK|G0.G:���^W�,)��XS#��̇��o�ޮc%��XP�WG��V0��# ���e�U�����6�����"�L�?�>a~)E>u�y���a�c��4Gu#[��r�:�Ax�<�t�TH�����g@�\w�+�FL��U�O��Uɟ��M��["~
)���'��T=��<����d�f�(1�b���QX$�!�~��o�Aθ��嵛>0j���9E���64DO�2E[�dEgt����h�#%� L]�5�zs0
P���:�2���}�X4�l���%����2KE�٣��p���`��t��E�� ���F/���ia�x�����?�4�o�:O��@x�5"��\cR������g3zl�aY���ӁP-�i���`�tD�����@GZ���a�翸L�~n�X����Ɠ�U�9�izW`q�Nŝ����0jo�,\��=�(ER-
k�SBFh�(l��9ۿ*�^h�Ji��&�ǧ�t�.4�Yf��9�]�1z�
ѴJ���L�t��t4\k��Z�a
�.i��B�1Ĵ�S�r�����xt#�g���.#Kd*c�`'�@����.[�A-���vg��}�CS]Ns[g��6š7�1uAt���s1��z���޿ZΝ2�)�c�b h �F�S�[�����-f�8�^ٰ^�!�̱a��J�W���&w'#1`K����Y�i�.`8#I�ߢ����]��\<�� b� Wa���-���MDN0���r�ٟd���M��t7iqjChN��	����7p�p��M �"`K�J7�y�'��K�����9���Bk��ZP[z�#Sz|��S0�:�I�9�PB�ǝ���v̖��=o��Q�� ǘ��>�Y��++@�ˣt��ȑ��N=�1����3T�ʛb�v	����Ӎ?"���f����T�E��e.MU�R�%�lI�y_-4�PC�d���Vn��r1�1�EIH��GN���Ldj�X���<1G��߳?�i�
9tﾥ4�@�.�A�s%�o�������w�c�L��r��LIG쟈a��#�U~�I������C���p0Ƨ -l��b��1t#�k�sj��t��u�m����FK�.��]!<fi���}�䶇2k����#�{s;���Y�x[�&���� 7q�+8%�3�P��;Ϥ]�:X�����<����p����aeCY��.��q� �g���v�������_�8��ܾ��9y· ��u1���Hn�5B�GQ;���s�W$���Z�� 0�X�Q�ډ��q�..��M胘 9��#�����Blh^I8d��q�@��M�i�G�:�"��o2��ޟ��s��]�h}37���������#_؀;g~ʟ�"
�A?>`<\(y�[
�=�v؝�Z�џ�����"&���$"3֣s����ӣq���"i���~�U��12��[AX�O���	�Ǐ�J���$~�B���V���0�
)z��}62h��1�C�		Ah��/�(��U8�[=��W�҇B���©z������h�2����E��֚\�Q���p{J��ݏui�+�_t�J��UZA*�R��lG�.k����]���}h_�T����|���$P��G�(��p�O�ЄO���*f`����*@�a+��C�����`�^"0�~^��;i��J�w�|��S]��: �g���t���̚�W��Lhė�%}�^YPA �|�`1q�j��
.I��U�mUm�3�~����m-�bӖjm2�R���c)�{�%U	����Y���j�]���]yW�Lц$� �2Ӧ��m)5k*Лp��b�ob�����l�F��5""�[��oᳳ��D�q�ƅ�|�J�*�^�7�>���|��#��0������-��?���%��B�ӷ�s��S���]�V!��w�0��۩i��hpH�˭�B]*���|ƀ��h��]�|Z��#[uV�wy��Է�# ���N��Kg��@�;KHM��BP���*>�Wd�)��D��<��T�IqKD����'"I�
�O���W��uu��_d�Z�w�T-�7�3�DjH+vڢ�b|������t�@�`�Uy.M��S�~������	ĳ|�+.(��߈�ta��+�Ķ')r���b �#~����fX�$���j+������h��r�F��$&P���l�=�֣�������%m�6�A��������h��^��e��=?��� w���;�ݪ{V����AR��Iκklh��>�*����_�O��c��HR��{�k�>�-rnl׽�f~�ƨ�Q�i_��pJ,%� v5HӰ&�t=Ślqo8�C?����{�%�$8�F����b��J`?��.@�#���8 �0-�ř���)y�_��{���I@=_پW};v��ۃ��}~������BJ��()��[wo��Cߖ�i��X�A�~-�^�o�Q�ά������X���6��K�����K䂎��Q�>�#���@��$P���a�Nf7�?����s��~:rm��zms�pxl�}f�o߇��y��c����:�I�zW�0�mіt
�=H}��Z�
K<q*�F_��}��3�(ưn?�	> e�;q��i�}�Љ7hc�T�[��6�p/L�L�?����+�4u�D)��9����D�ƞ��Ì���)?�0&G�h՝軷d�i|�a}V�:3����yL��׻�.NhQs�G�rY��ZW���Y������1 +}-�x?����w�/F�Jlm�~�
H���4�y+)�hR�S�xs�)U_cάf��m�5 �jUL����C��TP��8$���	oi]��g U�%��� ��*ᡖd�k^���tc6k^@�O��}����O�	п3�M*� ��o{JD�{a|����;��R��GX�x	87P9�w"h/+˙7��Y�v�_F�P�!l�dQ��U��XC�������@6��l�Ӱ���2�
>݀��Y{�ۀT]���%��HW�v�v��X�KP��w6�T�#���eiN}��~�:k�C@TW��>Q`G����]��xF��Y[0��a� HL?�!�i���׮�"GF��AHhqVS�-:���?K�0��]ᘨ!Lm�`k<�[�C�
�u���*n�no�it����:-��,�z��q�X>�*�P�c��?�*l����d�%u����F���@ �ֲ���9gϢ�`�z|*�J%g�o�3�����:�%V%�n�" {������gͨ��&�����C��������OD�������#��6;��e�S��F��6v%���޿أS���Y���bmy�܏}"�SS� ����JTg7�q�D�}�/�� 9���|����D�i�	��tS��,�	T_��-`�^?(��5 ���>���$�;�gH�����5����Ճjm�������7W��3�H_�!���1|�����g�(=Av�a�MVO,������&P¤��6���o,�ܸ��?��`��O��#59�� A)=E	�Z�I���CX5. \Ѐ.�ÝĶY�o����Wx&U��E^��\9��pbP�{
z�<��--�$|;�p���}��N�ut�[���rO��?�dIJ�[L�"��^G��)c�Ф�����v��\א>v���ط��M=�.IB-�����D�^/�',N����4���V>�������Ӑ���v�ԧ��^J�W��Jj�h��v-4jm5���xC���՟&<�����榻q����)\;�2;�l	�AbVo�����!<(�O_]	-W����aGDJ���S��T]I��H�.���F�pr���B`���"*�KU$<uc��ܧ�;ԉ��pQ=`�2��U�0,l;.X��{ =��^Ϧ�_G���Υ>���4�� ���i:�"Ċ\|�T����O�(�(��;�5#-L ΍�?O�'	g`��;A�sJ��h�Ϥ�}������7]DA�,�~��z���Hׅd�YO�Ku��X�D�*�W++����ߧ�&�Bԓ��:�Ԃ@��V�G�0���a����B�%�2�r�\������U7`I�+C���r�7L��1p���%�z%~I�ʨ�����.�H #Z�՘��^t�8����Һ(��j^�)�y����T������J�5>ыK��T�K�u0"p�hs��_��� :�?Җ��(��aO��S'�Z"b*O:�6����A�����l�H�p�>uP:�+���7:IW�+i���F��e����r隇%�H��P�TP<V