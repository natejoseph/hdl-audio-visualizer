��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CB��na����`�5��S<��8�M2ͫ��� ���r�/�jY�Cb'������غJ�ތ\�t��Ώ;��/Ӭ߼�W���ul���o�����)����%�Wθ>y��My��1�� � ���[���($�0��z�ɚز���ӕopah��{[���~�I��VEB'Mb�����
��`�\_�����s�;��	R#�v�10yn
������vD�O��l&��.Wѷ�̲��������:�%�86���&G��06�3��5^zÛﾎ	�{�e�N �� �]�\2h�n�	M���́�+G�����j���;�.�m���Io�U��K4s�A>�Y���5��-��{�f��R��놉&Q�N�K�e�O�'���o�L���QI�L���H�ri&T�>��]���3��m����n8�9_��5[��!����vo-Slަd������m6��z`��E�?��ˣy{U��0�ܼ2���"�%X]7�� r>��L�;�{{6�e6�9l>�FQ��\*m?��/��fpS�<���o��_q�_,+ˋ+�q4�
R�����^OѝT������?=�3 �P���{*#X�x�XD���(��_jT�#b�z1yKY�M���lJ����)��d��D�H&��Տ�k�_;���!�?�����Gbb�b���S1�P:�i�3Rd.&�:)xwC����,�V{{;��!�Vrby��T�m�#�$��0��j�M�'.��b��{���4�Ol�J�B�ﮂ��SnC֬�U�ŻH��x?�Kb��[R6c{N�{?{KoY(�)�o�|I<����D1/X*۪د�e��t{��̲�D�`��	��O� ,��R8'ջst���z��h)y����h����j��\���6�ls�F4v��N<����i�lT+J�ո�Zu�u��P9]�����Y5b���?r�؇���2�WZ�����17��ů"�m�1��>��8���Ч$��+t�#��1z<P?��?c�Ӱ���E�\��[�3v����R�G-ٵ���z�Gbw����R��1����D|�6%��xV��e�'��UL��ߐ����}���Y�E�)���5�JI���&�ɒ�/L/�xmH�{�afKce!5@\���e+�]Ȏ�AN���Q~�:��kLKF�zQ����o@D0%ã���uJ���9����t�{��+K�>,S0�*�Pp�1s-�ڣ[��ߨ��X�>��^�����0T�N���K�J�fS} ���N�ѡ������7���ϸ|�T�]����I�1��^b�J����[Σ���,�"5\�]���󜽗�:�����0�h���Xݤ���.׳�{���
�����N~�Lu��k���ǳPd��o�(M��ٽ��u��C�_���;�k��On��}��ж2��ٛ�gE����J��OJ�o�-���̓�tv*)}����+J�qDx��-��5��OQ1joϘ��CN�b7�4U=����Kshq$��C�A����5�i~Pi��w�������m���'����<
ب�o�������4xO�� ~w�Rn��JVkC��{1n�K{��d�Bˤ�nR8�X�=0�f���iU��Ϲ38���β�����Y`@���-�e.z�rh임�AS�����Y�L�VI8�����f��LI�q����	M���i(@j7̠�kX�	��4��0�F!X�'��P�x͉�O��ɥ_@��DB1����w�s��ǳB�=�$%������2��bg -K!�F���$vB8U�a�ࣤ�9���gg��K'�LtJv�����/��|�]|�C�"�L���@��r�8��,D[�.6*y���O`���h=�}'J �q��	�#`���G��s/o� ~�C��~T�����Un���a�5�����.�ʃ.�'�����I�B�
����ԭب��ʱ}6��\����h����S|ON�#�^�ZU�o�M40k}��o����ny����VJ<m�(�#4���3��G3�1eOJ�=��[�%puW�D&<��N��+��;���XBM�0�4ڵ��֠���S�ǏH���1:�7�L���=%�M70S%n,�J���n��붎���O%��ש�G$5n^�ho�r�����Z�|�b���y�$}�qd �wR�������}�nhd�9sV��Q�x'H��۫zW2� ��~�����|i���Qi.JZ/"��-"�si�R=1����%�Fh�q�7����.��W�:V)�Ex�x���k-��;{5)`z��3�"���aٜbe@��@�nϗ���"���捭���J{�oHp3�s+�[��u��p���c�0�DZ��;���Շ�grJ�Sկ��l��F�Bt��� hK�o*_帓�M��52���Gܛ3
���\Tn$s����X�먇Y?{����ޓ�#���C5���CК�i���G��~k2g��� �$�8�R�e��LZ����p�C>�-��5Ź5�mچ��`�06>��Vљ	��'C�
���e�XX�^���(G����-F��vU��f�L���DU�%��&�+i��4��,y�k�����	nT�aJޜ?�J`�������y|y��z)bn!=y�Yk��E>
t�Ͼ��c5V�gdI�@��P��ڄ�C9�9����a�ᢇCujC|�Sv��f��靍�]�`�L0����c��C%WdX�#K�_�^
�:���-�S��nx�I�������=�
��a���z���ڇ��k�u�Uڠ`�I ��X�eCDl�s���tr��}�I��Y���3,�{��尳 ���)�O�ೌu� �K@�T_՟FJ?X�:U޷���>6_v��:L�5�
�{��b�NrW��<§�MԮ!	9�fY?	1B��n'�q�3l[��������ܩ\��a腿���34{�T��6���8��!��\����m�1�N����8l��s.¡�0��.����`����S������J�S<��X!Yɧ_����R�1�;_�v9pI�c8YK�a�� �/	�7�Z��u������?� f�W}�@�HX�2+��z0Ǘ[��7�*K�[���V��qC[�v�4��9fP�uW��N��R��CZ$�}J��M�D����:�G`��rd��w��p��]ڎ��\�rk?�EW�h.*�5ژ@{���;)�_�׺£!��e�RU�yo�4Y{1��7`A���ڥ���"�o�u,�q�Rf��8>�(�Qu��+:h�Wwk��ZV��OH��YrJ�7	 [�f��K����D���u$G���"���i�j�V��-"�A���؋s[?~�O�[?2'��v(oЉ~R�X�/3��&T�l雹Ȗ� ~
�qd��&������=u����!�`�1)�H�W�q��'U�U��,�⹎��ͦ�>����8&RJ��S�t�E�T6o'��tȤ�Z.�d��]�T���bj��^ѷL�,].`|��1=�t����s�hc�
	?�;��4s�������E3�2���q�:eo�q���ao���cjG.���xQ4g�h���@@,:yEy�	ӥ���N|��H�Ke�n����`��
��ffG"EՐ�=�,D,��+F���u��\�u�l�}�:��p����*zu��P;%����Z��3����]�^���*V]��ڬ�_%�K������8��@���4��/�Wa�$����B+����P��*�!�*qWC�X�w������Kd��RIڊ���먐8����\�%>e�j�?�_ZD�����j��,�y�CCGЇ�ϡ��96����\Hݻ&Ϛ�NʑI��`����N�n�c]%�e
��f2wf�&�W>ia7��f��$:[oV���U�̊ʅ#�J"g�溺8�q�Xd��.�bהZ\6��"�e�:��xh�;�2[�8��uT狆���uܮ��hi^~r4b��>�g�G�p�����o�m~|�/��f��wW��%63L�-��]�f\���/�S���P�=���k��D��1k�` ȣt����i��>�
'8�<n�;j�`�Y��Z�*�zO�q�:�%7��3mq��}���C��� o�Wɼ��y礑@~��ɺ�v?��U:){"
%
�������}͵�V�cDmũ�ƿz�`s)��u�.�xw�ֱ�kw'����\�d���s� �'�a�H�����&9�X��񦲺.���$�N�������:gm��W4���$���>�kx�j&@���qѭ�5�n���KC����ɦ��<[���3���eH��汄�d��_�_��KG�}]~��xgU�i���ak�=��-Q<`@�&`�h!H(b�yM:���7��.����{����ԧ�pS���m���e^��(��e��%��U��U+`p��)�wd�j1�1�.Ā�b��x���EZ�;���F�^7����)Ci�>�5:1>�t }�;��3�]�# �5��H��H׈���3�A��{�a0����P'���=J��[�d�#���M'E�����;�(+���\��������r�M/R0<�,��L [��p�d��&T�8�0o�������͸��@ S~;R^7��د؊��N�Qe�R����/3�s����� k���
;��9t[a����/{�K���P}����^zQ�R+�F��s��z��Q&��&�2�k 1�� *��#���k��ۥK��m�[�X���j���f��vx`�`��[�Tm�^� c��t� �`�~��"�.��[>P�A��s��v �?�\�N=hC|_b'��۸ª�k�k4��^�{@<�Fn&�_R�v�-��Bu�[�<��j��b�mO���� )^\<����>�b�v�����谖1l��e��\I����u��t�*!���;���{)�\�m�j�OW󻡳���3�Gi#4�c8��k0@+yKaZՕj��O<s|�y�+y��>��3V`�Re]w�?}�����������ޟ�p� )�F,H ���ϬI[J)|IՖ�\�66����s�G���y���<��Tģ��zk,L�ϷY�/s���i�r �r��:,���RVF����@+CM6]@aX\Z���_02Y�0�� �o�vp�\����jx�<���zA���	CO�7nY1p��bP�v�Y"� �xq��e�V��蕝�y1Y`OD~�>�X�e�>W��4ߚC�IVu:"�-�b��5�@�P���e1�A $ ?b��Ea���x���%�	�E���ԩ����	���,Q*U@��:�l�S9�ҿʺ�g@w�ѯ�:�	��ԧ |@��*+��o!��e�H�r����Ʌa���:ڢ�YF��\e����m�L�:t�1��-Cg�x���Z�����or
�Z��F�m�+��q����L��@��"5��Wy��A6*]`
�j�H�+��%x_R�_�,x-���k�fbB�w!�=���/�f��0P��&�
>cő��=`C���K=�9H����2��`����x��Gܔɭ�{b��zͱ`�X�9�eB��`n���S�4�>����S�b�c�|�=�^�3���@�y1V�,6��#�'�|THĝ>O7/`���v/� �~��ъ���&�R�͖X�#�K��l����#�IҏS��uh�;
Xv�$on1}�W��ַd7š@
\:s���ffn\!&*��J5�0!^����	㲇^�"'�T�r�%n�V�]5�p���Q�$8T��#ݓ��됪�c����[c�3�X%>�=*�<����Z[�;ǡ>u��ЍW�Sf R_dT�`��� �#~����猓��Z��?�YSt����*jP(bĩ1c�Y؊�lt��,���E�x�~��0}�Y,{m�Wv[�d�v�P��w�����2v����F�3��ZU��,����g����v��z��n�������f��D���a.0���=m��-ޏ���Ez@G#�L�.e��G���sR\ǅ��L�3>l������[�S��乄�a�ɥ��ʩ;�?� p�P����8_7�
5k<����.��ͅG�ǝ�K:d�1��{������(�"�����Ξ��P=�f_k����%������w��H�;Qp]f�0C�s���G��
��'�İf���tƩU
8fJ)���=tc�S�x*e>̰m!�ח(X~���tn��2-�b�`���[>���@�(��_���#�
��ڼ�,.x�wKx#['@"�Z����#����$Sn+a�����}��2͉�e���٬�R㟡�nh|wV4�x}pW�v��ª+*r �Jk��kmE'����XV�Vf�Ͷ�A'd���cS�Z0}ԩ
����m	�S��|:H�-ۧڧj7��z���>�и2.�s�Ga����m��Jǎ��:��!��~~�7��?�Em�/��𙋜 ?g�@�|WrH�DO)#O�O�����Y,��cj^�a5b����t��(�x61H=�j���?�)/g����6'Q�i�;���b�Ҕ����O&�.�n�"��^λ��0�������<�W�8BjF����a�uw�,�<6W���u#�p�4j��4%�ʀ�p�=0S]�%�F�t���̿q�ә�ZI2O�b>ϓ���N� C&D���w�l�g�p��3�*G��Z�;���lT�O�� W��`�g�˾#�T��	#'��`����\�e&Ѯu��C���S��'BOW��"">�*��~��5z��'�9�r��%�N���8����%��n��P���#��ɭS��y����̹����<�7��J�d��0e0��B`H�� :���΁�&X�ӥM�ϖYAo�}��#Z��q�@&�q"3A-F�d��`EOqY��.$�W��؜F
������� y��K���^���|�C�2��т�O�V�t�9ѯ�w�;w����V��~�}�a�:�gd������'��`��˚1)���we�=�Y��~�5��}��R	˧�}U,n H>K[�Fq�Ķ�R��.��������q�?f(b[ᎫAja!P�l��g�IEI�B4���F`�%���ԷQ�D�A]�6jO��o��O�
-R��������Rd�4mi��h�_��+�0g���DL�+��%O�a����j��-e����]�[5��3��]=,�Ж����p���^��o���u	���K��N�ːU��
�AD,/{V���ȣ�BC"uv��=i�`πx�ǹ�����*�Nuص(���J�����r6C 3�PW���H�N�'o���B��HX	�(W��DXF�Q��A �+�y�+P �E�B���Ў�X��ep��CfI��d��Q���s��]��k��vT�P��6�����߻EF��f\��[s��I4�Idp!Ui�.��r�p`d�b;*���P�ȶ�`����c"��Uk�Q�w�9Wz���1=�y��r�wW�VE�)G[�<��7e���e�W*wɝTKߍ#�h��Q���Բ�Ot+�׎�:$��{f1���lZ C-������?�8��}���.��$����R�U�ʛ�:su��zz��S~�1�o��A9Y������:�S�y���%�,�>U9:��1��(9m��;��t��x
?'d�f<Y)�s��:�ϙ�C,��mxu����V�<�AKzq��t�i��{� ^Ev�G��%=��׻I>�x�Z`�zy+O�A%�0���Ӯ'�!�����S���k�h3	��o���0�#��W;0�����T�{�uA�
l"�����ͳL�m���榕���	�`t��xt��U�?X`vT2�Z7��A���@u���^K^�'���82{���\\��W��!�յN7t��$,
���'��y�����%�r�:�/�Y�Au��q�m��9\v����Q�u#�U���XS����Jy�v�9rK"��f�ӑ���s��	�1�Ɵ��v0���~Z�9��ۭ���v�~��k� �S��ѯsx�J^���@
GX�[���+�Zڲ3��`�����u��F����-��y�?
���<�hx�c~��۩2��e���g�g���yJ�ů5x�"Cb��2��|��Y��h�%_�3{���A�����/�辘�
"� ���'�u��i_�˗�a)9���-_���h4�aa�I`�K���s��w!M�J�4	�L��L��ޯ�M��r���@<H������E�t`'l��d-�u&��a΅�ӹA͛�M	b���y������^&�Ǎ'��}�W�khKl��1]wI1uu.Ǉ;|I==����{�3����W
�9Dw���s"�t�E&�G�R���n3�m7!�A2 60�_���j�4��Bz�|�ϴ(U�y\̮B޶�V$SdWy�П�$+���!w�LS��iܱ�]QYx�u:�P�ῤ��<(��%��۰N廞��vfq�H�Xv�-^7C�J$�;^�|w1 �Љ{h
�NG��f��߮̏ëO��S�K�Qc(;�s.��Y���T%P�ܫO��?�<�1/ô��o�ƺh����GŬ!��?{����ǽ�x����K�4mJ�����W.eN�;�~��Io.��Ɉ$�Ӆj�j��6��PN�8~Ay�؀�\܄�_p*?�0Zú_�%�8��z"�4?qh~�H�G�Y�8��Y�^�c��?�W����w|�&��-	S0�e*� �W�]Ãe`U� G����&ߌ�Д6�I�ӆ~�%���^�N��,V���*q�C��?Is8�t�X+q��n)8�x�-��0X����c5l�)�^���J����˂5:�̶�qxl�g�֧�u���ǀ˥��
��X�y+��y^n�w�q�f�鄅� )��P��O�~Z>�$�����?�
p=����Đ2e`�_?L"�8��U����iONS�ckA�b\"=~=QwR�:is$�8js��a�M�"�����6��U�=�j�@�єZ�U�(x͕�P!�(�y��k�y���@��pj�2+�P�4��������Ro�tu��]� ���~B]~�kx�p�Y����ǝ��r��0�W�sV��2���њr�XJ(z��E! ��Z������`og����?ʸ���l�._�/�p!6B��x(�v#��P+��4x߄ר�PU���l��IoIUDzu�v���� ��������p^Dו���SF-�PO5��s�z�>���ɒ�	/w��W���CI��1���H�*����-H���5��6^��"������z#��E#9�i=�He��l8�0�L������pY��j�������a�M����g�E����Q�И4K(�����~��~n�H�)�������7�^ ȗ�]��ݟ���:B����GSٙ�����-�"
5�1p�*�
O9��A*�T2���D�G3���A�MC��SH.�3̭c��3Ђ�ܙqz��QW6���>�����=~���ҋ�<��!0��͊T�����T)7���Gh/��S���{�/8�7�����4���҆��xG�:f�ل�̼ewL�J}��{�a��z&!�.� �+0C[ö)����R��������+9�#+��W�1�v��f��Y�.+�N4��(%/�}`a����9��(���	�z�v��C��8��ʭ�r��w#z���L�phZ&��&?����GM�P��Jk���׽PSqܯ��j����^����P��D��>Э�ߐ�0l���	�R��tW��"�B���"��΄מ�X3��b9�pq[�h�����\�~_�_0O_�.5_��c�2x�V"��ץ|�_M����p��ѣ��x�J3����$��FlV�Jw'��Mg4hhCK���ً�tw�~|�И���>d��}�P�Tvm�U��[郋
�2�����C�����0�?��/�lp���)���Vq6�	�����pS��>�7��f({Y��J; ����3<�	��g�&(;=�K<� ��$CW)��89le��+(w�o�_W탘<�Ao�	VȖ���1:�!��p�I:�Bs[�|�Z�\Wj�U������� ��6d�p��M���WG��@5f�݅�+��:6O�W~^�5�#�#���r��Ov���{��(���`)�4�֞5'�g�4��0����	ތs��iʻ7����������S<cJ�ƚ(�d�����T�f��^$M�[��&s=��0�9�
��֏�p�Fv	K4�L�EcD	�yA��I`N&�M�9���gs!��M�؁%�1�
dp�j�@GW/U� أE�b����+����3� 9�U���<��#�6��k���HR6tf�m�v��߈����J�Y�9+ԛ��W�p�yN�.2��jŎ&S>�y��:B��͌�T##b�؟�U��U�B�r����18Ěf��m ��wtZ�=�U��^�PB�N&��3�4��'c/(�"=�	ok�N�eֶ��~�����n�����J��Y��m�6��ij�����r5�h��G�a�	���R`-�!�,��5��t"|�k-Ǉ��D�9��t_*�	^�*����7uuj���I�\b3�,�:`,�L/\[�n���":��Ȣ�9����sB�'e�A��[u�.}��@���*�%��q+�?����X4y�2�J~RC�f��w��|�,������"��%
&Q!bQUʖ�D6��B�C7��N,�f�ŔʧqE뿜�W�3d�iܸI�����%�u�]a�[��Ů�QP�67��L"�#��ΓN��W��:fw�L�~��X����DO�����	?�\;�6M�^@�f��Z��-��)0�ɧ��J�͌Z��r� >���<��K�������ab~�(+hO��6l�y��<My�ψl"�)i��Pde�T>�]mb�:���bD�:���!N���������X�,C�#��N9�ͨ'��S�6`L`�3r�/�(J0t��FK����ib&\:�q�cf>a@�k�����X�\a�0[K�:$���<�4D��f��7�+��3��ba���[�����|�k�ӍS9.y�`�'�>��v��4�m`�Ơ�ۈ5���;�t $�/�C�|����w�����5O�4��h�H����\���~Rμ�Fs�#�)��^RNji���;�T� ���NS�w�N(;�T��d.�0�Ɂ�b/j��ZOѤgo�Ǉ�&�Df���t���5֨����6?U8 N�7!�����֛�Iy�&����X�7�qj����S�jm�h�0�S�|�����@��md��d6nS-�{M�r��bD�l��y`��x�22 n9��
R*����tcT���E�:��?���oe����S*��Ʀu��@L���ov���|2"�T5
P��ٰ�9g"~!�Ǧ x�m�ӮI��*��W[a;�ow��TT;��*�)t7g���gS��Å )����u 8y���apAJ�*����ء1�~BTOX��V�����Y�M]�ȍ��K��>^��8l��P ɣ�'~5��R�;Ih/�.qo6��ٟ�t���m��W�))�9:���3�M �|ʂ��T�׋�Ex;�)K��1�6���-&�����p�&ħ�,�@��%{v�p,ߙ�����|����G U�S-��9b��Ơ��|g_1�_-{pN����
<2r�"�!݃��f�la@�ћ�Sh��A%��N���-g�[3U�q�,���]@�{��#��?�#��5Inm����<��U}�C��k�߾�-L��{c9"2��;y4ݱ˅���I�)2��UD-=��a&.��S�W�]��l<?�Φ�H�M)�2��곞E�p�R�H�E��V����Az�Z�i+��C�Ҋ=˴�?��oI��*^<&\�1u�(*K5D@$/��AAT�
�y0���P{5�jDn~`s2��3�0���{hӍ[�V�EA�l��ZY��b��g�Ww�L�YU���S��ɇ=���OYQ̗�>)y�U�^��/��l�+~jKYL�2O�1�ʏ��l����W2V��>�v��G9��] �/�4���L�*H"/kP6����~��(B�u��✤V�0����O@g�����P_b`0R��\R� �c��ӣ#o�]��aU[7��+[e]���:�uQ�)E��c��ꖳg�/����S�i	芗�
�����̎�LT�`)�z,L��������Kܱ�HQ�ĭ[|��`��'���Î$�J�� x�pq�k�Q�4���-����Xa���H�B���|ۡx�T5ʴ�u�)��{����g�,VQ�A�b�<�nȄ�s4۫�FN�������'��S̀>���pZi���EFԖ�DS����4�+�ߵ�H���ڥj[L	�P])3�c���E���b ���Ώ1,�#�'_x����cʃ��}��R��l~L&F���n�H���֓m�a�J��z���e0�ɸ�/�2���ǯ��t�q�0��}ˇ��s�p�b����.^����$Ѫ�ԐF��Ea K��1g�[A�'fYq�/����ƪm܇H���I��s&�bh��w�6�p {�ۦ�f��7�ez_��(��
J�uv_c�+�]���F���s�
�\~VfW����z�8�����S9R(�u5��J?�1�!����M$��5�:ڧ������e@����\�J<j��!\N�W؈�A���ט�OY C�#iJ����VR���?@�"�'?��d�9�S�믢�.��bXX�����C�dzҍ��(����-r4k�}�Gm�	�Mx�f(�Q]>{CEW�4�ě�p��ւ܋�+��t��x��8^�F_�)�$s2����w��s��Q9�9��n���v��e�U:[a�~'{K���ه���s�UA��,�J�U��#�1Ƞx���YnQTy�ő�b��%�KS��mQ�%�����즎����~�bK@^` ����sQ���"&��é;*W����ݯ��rV�D<ǆ��h��s7��m���0���-	^�Y��&)55ٖ�gPXbl�3�u����K�D�
U�֎H���i��y���=p��c�t���(.��t����xn��!����D�
{�Ɠ7<K��6�c����G�*:GC��
�q��2���^�Va�~R9��R}��P��b�5����r4Qe���q+Z�-�"�����d0Esй��w�vO5l��ٌ+�f��p��+��C.�@�Ij�p(;�l�֖�M@E�r8��@�v7>��K��eHy���Z��EM��P��u��5�d�X�4��TeY俛��F�Q>�������f��8�H/�%!��C�U�d��z87&�th0����S/�ӫ3+u4x/�����R�/+�;++���T���ˑg�j�ʹ}��v�����2�wO��"��\\k����*�]E�2ܧھ$S��a��r?Uev@b�K�����-õm��-�ưH�͎_n��]��-���R��Q��p*�p^��|^MkT"ANy��J���B���X���Y�s;�0Β�yj*���B�Q���_I������~[E��� hK�>1"�@v3s���O�T���W�L�l�ESͪȹQ[�K6��nx��1����C��_����@������v�/R�oɐ��T�0�������T!�@�4�i��lg���(}���8���c�]g�8�V�U�W��*���h��H�"��T����>��%=�x?�������.B4r�3E0ߒ��%��\����z�&ɿ���a+�f�䎜���$M���@�򴠴���Xzߦ�K3Ϟ�#2��XA�0 ��iF��`����0�(nﲁ�$Ь�.����9T�R������9�5mݚܖإ�y��&����P�lslg�L�o$��H�j��qC���y�>YgǾ�cdv�z��$�L�Z��湍����N7v���1���O V̉�(����݊��e���eY!�j/��T=y�/1�냚�O%U�xl2p�I��kI�]����I���B~�n���j~�έ��{DO��f�e��6\TW̍uV�p;fX���(S���X"|�Y}��%P^�v������bI��_����㾤Ht�$Ny�T��ės�&���A��E��¶
��v�R��lq�}tQ�8�Ȗ���Z��P���l˂O�L��zU�	��jU��'KVL��oд+�ci�^�_�	֞��B��#�4��'�r�6Ri�����wӢ��+?���g�Ͽw`?��E�t�>m`0�k�ĂW��4������9x�h
�~j���>[��u�.��B=����=����,�1v����������a?̅����TU��\�O��t�̌��z�MN-�L���б���
�:��Y
�H~L!�֐��!�D�>H��/��ˉR_r�ϭ*>�:���f��K:��ʱ�@�nmrc����A��������\���v���X��sr������pE���YB�.��$<�S�
x[d#_	M�";-g�h�r���z�Y%���EšsD�x��V��]�+�,˲8����qJH�ziZ��Y��s3������3v&���iIL�� �߁M����u�������s��G4&��k��X�Z��8�@svG�ݼ�Tڡi�|�'^rz2j� ��l���(w��q�����7�`�<��������tC{bk}�~g5�Y��޼�|BABPV��3=���`�T͋Q9�����g�����q[h�J��u˄��Ԧd8n@��X,�n@J�X�)�B�����6�ᐰa���K�c�]5h���|E2T"i}��Ȉ� ��߾�kj�<���_M��� m�hj��v���� ��]�F��Y�\���+�<�>
u�y�5a��]�gz�3�����"C���]�F���u���ל�����8-Z��ٟJ+u��N[J}dX���F�3�쾳�&���a����6�مi��?�|Y��4��g�̴Ȣ�i;ۑ"t�i��q��n�����t�f*���5���3�u;:��7Q�3�)!H���zN�(n����Dd�kB�_��-x&3�SJ���ȱ��Fb�Uo1�cA��Ù�7�H����nU�U�j=wKdo�tZ���&#B"��Z����yG⢮�/��*���{!Eأ@�ɛ��mw��j���eP�X+�r��4�/S�e��H�������NH���G�Sy�3��+��K9����ea�K�Q��n__ɹ&�؝i�t��k��T��dp�C�>-ɬMP�f�pc�N�����
7�	��f�9��.)Ѐ�K[���ms�\�\5È�!��A����F�;���6�zB�'��vƧ�a�i 
�9*�޺��)�B��+1 ����Ԟ1W�H�d" ���*ӝ ��^3M��U|�EuԜ�P0�^���RI��)���h��b���W����o�t����� }jt�X_��~;���IX	A�+��嵐7R���wZj^%�ar�����°;e�8	�+gy�b����Ƅ�B�Ȑ޺�n�c��bn��� � @J:ڢ��yO��V�<��*D8��U@|7��$JN|Z�ß�nF#�N(��s4�<�zJ����=�I�L|A��K��N��M.�:��Wߨb���զ9ă��[5qw����E%�����_�*%:���'��
+�����! ^��9S�]�=�YÚޚN;L�b�b�'F/�e
���ni�_"����X̀��$�6!� d(����s$�61 ���3�p�����)�{���X���<Oc��m�>o��:�GɄ)�?Ra�6u��)5�L2y�y4�]aDw���_��ؘh��J���v�VE����f��|y|v ����D)T��3��a|S2�W\<�Ռ��s]�՛���� �#�{����H:Kg���5|���*�Kv*�&J����.���f0�2�=�����_���X�T	}�_hl�O[�	�U
W�X�V�ťN �d;�?��P��t�����A5wW��6H�mpxx�C�|?��>a�&�#�
7��O�����rf�w�rJz^�2/���EC��v=�y� �w��,����o�!W��V@iU��(gH�uW�h\�M��:��
.]�+o
�Q��〡Y�,>[F�D���[��)�| �X�#dt4�e��qD�E���R��LP�c�k�a=�@��a!�S��I�d�^�e��Kzr����Ԕ5\
�>��Ys4���N��խ��	jl�l�-=����HPDvʌXq�+��a��=��h����_���2�F��P8o5L����[�Ao9�c�m�G��Q�`�('�^����9F�K�GׄҬ\�H���f{Г��O�*�6/syw����]�b�h��߸4�i�l��g��Q�O�9�����Ͱ��ӻA��_��m|����3��u��~
g�w�ȵ�R�@�����e~Q1ߊ�3�r��)�����|>���q��)#�,�=.������r�k��j�W���Fi����	�~�|��`D��F9�o���\�gU�K]I8��>,�:�E��Q�N,��>D�E�J�x���4�E�!��t���7+��	�O"������e�bQG�vLzׇ��)Q�c��qe<�7u�Y#m<�s{�Rh�O��<��z�P-�N�7N����~)��*�g�S��3��F�T}G�������Ŋoċ+�Mଧ��5��DϨw�la�'���@ݭ���oM��0d3L}�2��ٱ�Λ�[��$KԌ�CڷT^�J˦�A�l*��JX���gݼ0��:\%*�p6�H��F�(�䕻~����;��'��jC��fj��C��k�^{��)p9��嘣� bN�ըȊ�#us*"��������R�MT��ra�q�1"�PR���f �
�f'�%��Yf��Ѹ��T�m��r�$m[��zܺv7wH�U�٠�d��\���Ui����Z{�G�1�<BH��s��d/��?J�顮��I�K���d���=8�6ϯ[�y4�țxg��̭����ŀ��L.���d�Qr@��L�Ҁ^>@�WsRI��~Yw�0��Ü2h����B���ڋ3ݮ/�`ȣ��Tdئ?��Z�d7C=|��(������٪�c;m5�c�7��fK�?�?�[�����N�"v�^�ͬ��3&"+囧�Z�6����'_��~QHqx4�y�-#�ɡ�8`�"O�Ip_6a��z��qWo5_c����U�|�$S/Rq�iQi�r�7�����NdA�F=1&u��K�s�Bv���ŹK7ש,�b�:i��k�g��������4I�`��/]|0ubF��܃m�LO�^�� ��`��U$�a� g9RL����J�9!�X.s�i�8ؠv�x�V�g�)�䧧F3w9�s�m ����ar�����+_�ȉ[�:�f�����$�����`G
"~�B��X@Y���y���G	�f��*(�l�+�b$�e��*�fm;.���*{�{�{� �2���w�kY�X.�K�>9F���G����{%A�+�,Bp�;u ,@R(F��SI�h�T}UVr��
�8�g�Ȓ�ӯU����i�7l����<�?[ݱcR�=��w��}��Y�-8�ċʖ�����hN�Т��Xi����#��_�S�8F��*����c�^_��8�/�����/
�7���o����I�F���y��9�h���Z\|�埐�%��*4;Wn�k��Z3�~3^����F��QE��V�t��7�Ī�V+��%��c�~Q�I'F�Lo,�/���+svr���M��"�U$��~>�}>4/�k��gQ�t{<����h�9�保�y�{�.���l��r���I{�Ct�ZK���ش����.�C{�㘎YF�9�l�<�8�ȵ�:Ri�JbC�A��Չ���r#jZQT�m�|�g�l�
��e�
޲�BNq
�X���*���a�,�����`�Os��279�&��Gpd��8�O��a29a��&�0�PU�#��k����A���i�ge����ׅ���s�5�OY�lvs�����,5�@��8�ў��ܩ�ޔ����1�8$l�@޷�GC�#��S	�Ѯ���}��"� ]�G��.Fj��{�-�!������{7%�C%K�g����f�r�����Y�~��a�8hj��!7ܥ<��;`~����Elb��9�&��ݙZe�<#��k\[{�-	l��T��$���',<.2Q��R�l��n�3��>�qL�tYnt��~42�rڰ�����%B���-0�E4S"�`�IW�q��v�/�S�.l\�j��ڸ�2նhf�a�V>�3��6>
�t���b�5c�������|����u���W7��-ҙ{;�4MWG�Ιѥ l���vB�ڝ���K U/�cn��)BFm`��nD�0q��m�'h<����T�������0������D����P���	���@\�GI#X��]��_����W�#k�	�B?#�R����p�A�0a!�m�_l��lkʌm>��0�T �]�gg`�������F�;m��2R9�$7��v!��(H�2�� �@9�I�S�<|�t� +����[~�0a�U^=ûR�S[4��v�����O��*�13�������!�+��_�,>Z��a��a���񆩑�X�f�0T��u�(�yG�?f.�z��V�\�����ʏP�VS���9�:r��O!���u�Y��M�<��c3� �����L6�s"x2}��b|虠�4�<�m��m�V=�~��}�s�̌{o[��ٰNe�=N�7@�䛊�,�	1c�3$׬��d-Q3
�>�Kr�꽈�St�/��9�Ǐ�#1�t��;��+o5��c*^�tt��B�ih�k5#׏���4;���YI�w�y�+m�5��5 ��!*����� ��������'��[:�t�؛aھ}���T"��g "Zݙ��Pϔ����_��F{!y�K�S ����GJ�FJ
u{� �������(wm�E���Nt#���1�i���?H�=sΫ����><�o����)�|�'����iUp�PY
T��z��_�k6��]� �l��������iY[��J߲ɪp��	� �V�,PN�6��_�[b^�:j��cS���#OڭL���/���r�ʕ5o/��@�di>�羯WL�ha�Jt���(��J�үL�T�n7��'��x�,N���@6?/#���/�D�v���t�u2UB�r�9^�;{yJ�����S%錪>�N
hCyR���X�vwy��E�������������8w���3�S���#���T�r�l��P�������E2x5��K��,�=,�wOH���:�^>c�I��Ug�F���'Q�mr�����%.�/�ч������b�*a{Vwa�T����'� P5�!���9�ay{r
�����O�4�$�C��ǻ:_L!���3JPj�zTn]U��{�FV��o�ǘ-�ʷ3D�t�{|�m_.��pa��P��֓���\����a0�2������y������\Z��5�5�M�M�j��	��`gҍ�|Kw��v���������o�z4�|
��(��G������5�~������P,M'�DxNq�Ԭޯ�uT�m$�U���aϾ�A�3�[�Wɛ����3܎iJK9�<�v�f���V�!dv5����^(&Pֿއ!��t�|��=�V��#TQ�ݥ��50�@�g��ʄ��=�?�?��r/q����MG��?�=��t$W���[>�0q�Ww�̧�w���<Ο�_:W��q)�`Z�{��)/�fB[#�������1��J�1)��حj�wKR��[���$�L�dӒM���0���Һ�Oť�q*����e���3�����v	A��i?��ޥ�Ա[�W�,={��n��8��hVLl�����:�J��Ö��kԌ�.�:�I��DϨxʥ@Z�&��4�p�m8�:�<����P c/�	�x,�1!�6��e}ۛ��N��Ў(�`Z�� O�^&�l@:����j�5%�i���k]�>x�`
���s����,�Y��Ia�]�Z<��{�dC�ع���&P�-�I��2�� �[h��g��s�$]������f�b��Y��R7��� w�E��9	���F�0ܕX? �bv�aا}���ZQt��Q��e�Yj̅���	���'����?�)������Z��8�f��H���&���'�vM ���}#	ݝQJ�%��~y��C1��K@�"����G(��߀��|�ƤY;1���HV	�:��ơ"���1k�£�����5iW�XPy�8��3����Y1�C�&��bt�{�M���/�ª�f[TBx�Rb��S�-�W����o�iw�c��UC����3d�_�Lގ�-}毺}�e�������%�EԬ�-�X�<~.��5g�h�E�����S������W�������
���w�7��:9y�6��r8��1��ڎ�1��fc�i[`:�O&���Cu��C2W-ܩ����\U+zӥi�V'�j��_�����dx�����st'Yrҝ�I�;ǎD7!�>Ý�s�n(.��$?۰!`�v��|�#?��\%1P�?5��u1�ÂR�!����H?��$��A� jhf�Cum�^�k 9��7��7M�#�Av"�%��੢���5�?x���[�X�������	h��}���-�ًEy�����DV�s�F���#la�_T��;���N�7%�SP0������4eObܸ��� �ȥُ}��tQ2�ut�IN�4D����ClO������3�2z��I�����G�����V�Z�+&�J���@�5���.
Yh�@����T^�� B|#*>E��
JN쨐M\N�g4�[��Cn#�}�3�Zܫ�F�챥sH��+4�xf��-���s���q�oq�zM�d�{*�J`8(��Y�)R����Z�X�/bjzC�/ẘEf��¤��>$�d�0�o
�`7�	�$�K�(�뉂2��%QwJ_�4W�5����&�Ap毙�S�+��G�:�S$J�X�c6�#�n�-*��g��K�Ν�7�@����į��.�m?/{�		��0yH�d�l֥ZnnmG�u-�U$1`���!�l(Al�� �K	�0���(����m'�*<�?+Al�̘�c�Q�š��1���I5�!��������&˼�l�A�I�ؖ�4��v�Y��!�!9����t(��h����^����0�(;��l}&3�<�CRl�V=ip
tm�qi9)�YŤr&z߮�V@U�?��Y�/Ys��ƹC���*�y�WXsa~R�^�(����ո���ԀB�-��Oa?���t����]9��.X�|r�o�{@N<7�k�0GM�2QkXg�+DvՃ�`�#��k��2�0	;����.�b	V'�G_Y簲t����șC_����I1����X�:������0��7�Dӽ�t��vc��V�:��_ZS:]�_a��:@<uҡl��-�=O0������@C�Z���0��/����%���7��o00L#S~�!��[��K>�պ��A��!R�7�D���Iii+f�v>�=�HS��Z��9��"U�97]���Hhi���J��0�iq$�O&�����:E�E]����*��7\:�kBg;=ac���i��z�J�
���N���N3A����&e';1-��l����m}%�̜�X$N�y��?�~� ?u`��jc�0E=�IGaA��g���ŨXai4�D���s/)L~��O�����3���Q�5cV��)�yϒ��]�@� B0Ǐ焢D1���ѭ	18������@B���%��N���;�&��Yz�k5�B��]�ܒ4�yڎ;z��Z~z"�:]��vh�b���>��Uv�Xyͧ��'� ��Y�N*ӄe�zG��V�{h	��Ge�C�W�U�XޙYbW>j�
�8�ڱ�"�.o���ŐnHd0��O�	j�}�H���mzY�8e�<�\Ztz�p�C,��#�4�݀[�dT^��	�! �Bs� )֔.�����т>�\}���o�
��-��]�bh��TNoԑ���y'����W��b�>:��@���R���'Ed�${��8�uH��L(�?9)*U�eqp�&5���-��란����?]��m��`饀��Y9sǁޏ�K�?~�6Ԫ��~A��:% �c!������2CrȌif��UY���Rb>U��X��ʠ=���mS�,�_Lm�:xzqi*��G�Үm���:��v�\w��ϰ�uӍ4�Q,Z��
<f�JA�Q:�\�+|;�?����r��l],pU�����j��yk�.'�	K�;�L�Y�ǀ�yy6����Q��}�}qm> ��R=QCp����Cx��hbx7~�cf.�K���K��mJ�p螚��1��_�B\ ��?�����@V����`��*IӺa�/�����
�q "9�juNS)P[�a=��̥(|�u��l�!��~yŀ&�Fݲ`7�w�h�'�pt�O3?��)L"�v�G%,�i~��g1�b�5�{dd��b�ǵ⌌4G~~�,��Q��M�K\��e�I�TV����]OҜ<~�_�qs���9n��TY��w���4ɾ�9����@�}����S���S���%.�	��HҾ 8�V
uy�����g)�.Q���a:��L�	;bXH!�Gl�u�Y�ZX/s�c��{)�XC��h�����3W���2l�JQ��.�a�Us�z������7n��r�u����8�%��ė�m|�܃Y�@L�x�F+3��~[�8��E~�b��x�J`��E`؜BU�R~������s.'8�i�&�|�x��Ԃyl�Jb0v�2�E�P~D�f���)I��~Ԍ�R<���
����H3{\0a��Y!���s2g���q�����8�5�̽�T|��F�>_�ob���7Xw�)��]�����#� m�'��~�rP`�����dU���Ft~uš/Z �1�I�/6�ǜ��iX�b^yMk;�i�t2!����$ �b�~~zb`!��2]@_�}�69u���������_-@V�c�#J؄��xve�8���B����vF5sY�.��)O�#�e2p�X�	�Y+��uݻ<�,+*�s�����m)#����}[o%��XS��t�ܺ�$~h�8��2K�@�2�Û^B0�DJI�����X���>���^`�J\qS�6?;�J��1�� A�y�ʙ��͕�nD����L��7<ip��e�)��؀�ø�u�B�	���5bs�}��� �u',z��J�		n�h[�/�K��q'WAoK����8xX���\�xi�ct�pH׭�\>
��K�t���l�@L��CтB����v�J�$PdX_������q�l�`�h�Q�%w�E�7�g
3����ɤ�Ogn9����6\���!�a���\�%@v�!Y���C�+@���j~k鯙��)P4��#�n���:�_Dх֮��e�����ia�x�H{�F�S��5�|D����A"��9�F}'ҋ�T�@W�n��6|6�*�I_����C?\;w9��lE��./����%� .ݬ�A�K~,ځy�D���3�W��@�@�b^���`v}c���q�����QH�P��@9�E�� ��|��݃�5I{PK������F~�;������A6�HU��k���{�����9z�gx�B>�q���p�_�!����� �$����V_��XTJ�����߶��f�ޗ�v�L�Y�&n����J�q��ҳ�����Iy��Q�����K�sSq�=g��l$���,���)��8���q=�@_&iQ�6RbV�l�?řܱ΢���2m��P<�3��u����L���h��ޑ�s�Ʒ����כ̍�.D��n܊V������K9����Lg͐*;�!�( '��8w��`�5����V��GY����w{�c�%� h��K����u����)�+=]p���^��`߰���8�[Q��l�MϭH�8�w�-7��j���e2g�3�Ͼ�R�����Q&��2zhj�ǉr3��A�#�ל�`V���*�N���9z:l�6�[g�h	�l(J �f0daw,�x��P������:�9��/����~�~���!ݥ�P7��?�3$1�z漯�i9�ﻢ-���W}�0Q���Ԍ@$�l���ҫ���B��XJ�	�RG{ ����B��1Jp�`���/���X�M�j��Ϙ�
:��"�"��v�v�y� l�qf�l&E�o��b�i���@��S������)ҫ��CQ�ۻ5 �:L��ls-������nX�����19�#H��7�;�LLJ��_�>:]��/���!�5U�s�h��k�PQ-9{_H�!ᆥ�H�8���=��+�yw��%p��K�|��i"��C��=��]�^����l�Uc ����بHXl��ZDt@�u�����髆Ϧ�+���W�������i^��l�2�w�Y���k�z����YA�5�мE����'(�}T ~ |�;@�������[���w�#���&�ˢ� ��̽H�<�k#f��j?��i����w��#a��*�v��!񷃆_}�o�g��ޏĸt�̥Z��n���\]X���|)8�!�m�&I$]�I%�a���O}��C��-���?<h��!I�0%�xf�x�<�a K�i�֬	�CG5���$O�7�����&��Bgʒ4S�p�~�����)�lj��	����ͫ,�Y�e	7�9,��K,���6�`䱚�,1�=�l�f6,\I���2H���d��t ���g�"ӵr%��[�IM�tQ҃��|!��m��L��E�F �^����l�:�����W��C��� tң�zE�Dh��*�S�%�����<Q�rvܚ�=Y�p𢀊�
�5b�BgjMz�+\�[�������J�6���$�
�4HSD���\s�{3��k��O}6���M8R�$�_��N>&��K�?�8��w�$�-!�r�Zi 5��B�R1���QV\^+��^�<�}.��?Ni��M�6�Hۮ��}Y��
0�P��oέ5nJ�b�£B�2c#'�_Z�2���&c(�(D��98/�tOڨW�{�X|2DzU�WvU&���z��U��.�a|�a?�(�0Uqq<Ѷ��0��$�;c9�����S"cF�g�U2��V���]�'Qȳ��N�����8h�[�Bw�6��m��1Rk �f��R>N~�>�@p�_����!�}K��@���p/@1���)K͒!Z"Q��;��bf�����w]�c'� �qd��qD�]!1�r�R��Pt�5�1و�7�9�aD!X�� �<����H�=&h:�.i��,n��a"3�"O���9NfG���ǫ:g��b���:Q���Q�;W��d*ZC-!,���8,��.�\8�b�F��"�0�>�����q�]��}�N�n���>ŻY&n�1�j'�K��	��SM�5������]���+2�Q��u�Si���#���q�7B!.n�_���`B#��W�yhD��z� 
�����!�����ѫ�2��F�OU�۶�h=�%r�cL p�Y��̭p"�]ZEl>��K|����,K�l���XH���3����46���t|a�~゘�gmK��Gt��.�'��R�x��?S�hB�=M����)3C�����4� ��X���Z,:M	�"�����}��n�n��0Q	��O�Q<w&���T�$;U��c��H�d�C�A3@኎T��FlJH�.^��6�}��.��]_$���}	[�-.��ffv���Ǜ�݋��E�K�ѿ�����,��Oiq+=fL�����h���Jf��j�a�Z���],����t�{�|���sȁ�:�úv�ܒ[p�h�k�r����빸L�3"��.`�Z�N���tqظ�6=�v����\)��a�� %$��Ξ/Rn�(�ǋ�!��`��>b��r�Vc��7@�j2xo~���d���al,$A�`z$�q�8�oH�wQL��g�hF�8����F���S�1p]�b'qf������y�q�ռ���p�ĊKTW�k���m�	���&��tג=,JU����W��z�sq�<<��f[��@�^����㐾U����ÿ�^ˉ,y,sk���b��EG�@9�V���I�責J�s�u��I�}5_����HW��Ǒ^�6��L�U~���_:ny�X\P��!K�TӒT��*R�/��3�p�,I�^�ɥ����
�3�Y���て� x���Re}@{�t{���=���4r
=�Ņ�jo7(0�meg`�������ގѦVސ$`I'ȫ���t� EE�AO֌��XO[d/W�����3�2MD��~��<D������~;k.�I������h1���c9�W����~j�Y!�����8��#�!/J{��7���تc������1��<�<�T'�h�O��)�� 
��$��iͼ K.)�f�����I,����C\�=L�TC�̄$�P�I#��hN���i��p�1O�����Z�n����'�k�J��Įp��3��e"�<!QPp���%i�Mf~�e���Ք�jR
ĉ��_9�Z{+���$}���!7@����w���hwC����~s��Y��H[Lw�tVt�pS>-{��F?|�n��\���Y��>f��y迿��\�pkμ����-�)'�4�V9��hW�"C�;����T�\���B�	�b�wA7V����Ǒ��lx��+C᣸
4̈́pO�}*V��G��&��"�N/�v��R$������Ms��<�eR���E�il�CJ ����PK~-�g����bh}��r^�y�o�h��T~[��D�|mن6�jP�SU��6�E��l���vQ��i���m{x*ULc��=Y�)�ݕ�4(����s	M���x��-��
�+P�Z�x�s��* �Lcr�7 w�lb��m����9�IȹZ�$4XõVo�rR~��OH~ke�6Qx��E�x=r�-&k����7a�����8�?���!._	E�'���{μ�	-?���_�c5��k�|:۵�O�o�fNxw߄
�&U�4�]]Z�<Yoz4��a��O���#�]?����&�
�*V�N+ҫ�Kd99�x2"=oO