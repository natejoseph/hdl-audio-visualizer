��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��ݷ�����L�K=�D�W\ᮞ�a�ZC/v���؟��� ��h^�����vi��F��լE4m�c󠄱9u�i2@��
���p~��k\���"�i:�
��%������<�ěg3�Gj��yeXD���D�Ϟp���ht���Gv��d%�
9x����L�P���ϳ��K/	� k���46z�{���,��$�6<ţ�r�B��A	�D�}���$�.�% ��V~��yPq��>cw��zɠmS�J���2�R9�ń� �T��ݣ:|�G����Nb<8쳞GW��k�-T���#�����J?�����;�~�O+}���	L�b�܎�<�.� ��s�D5�ƒ��Mr���B:�=����=+~m�:�or�eT��i�>�sYu�D;�����]��j��~�h �*?� d��!	~���Z�K�J��$;�|��,+�=����F�iר�%���0g�z[�������� 0�h3�q(��N���.+�'��m����[<T���S�㞠_$��`�>��l��	�vq�n(6�q��4sM+��k�65����C+
��b��/%<3��6���Vǖ��u����͖R�	T�@%���ɝ8������Y/Y/��V��7�$,8�n��]i�6S�c �����\����ղı�RU*p�-n�w)�^�-ݸ�����bV@h}ɤ3��R��_��B\3�л�M ����`�ی=*�ڬӚJj��M�b��L5�����~�[�w��Cj��|��2�z��!�gl��3"�2�@m*��Kr�T��n��<�9N�g�ޯ�@/�B�=r�fةP�簣<9�!�Y�_��,��ُ�t���˒p�E�e"���ڍ���b��m��C�}Y�9�n�2\�^Uos����ҍR,�l��n4�s+��B6�$��o�M��g<y,S3Y�b�|Eޙᆛ���܂�9��b�+�\c�f�:߾��c���������`!TMP�Pf7�k��t@�S.�qwƛ�l����"Ch�Hq�d��kba, Zn��1��Mཱྀ��j ��ץ�R��?�.d��7�q�R� ��k��}Aj�9��{}A��b�ДF�?>���u�`���.H�{�z���7-/����-�諡.h ݷ�N�Ђ���,�a��:Ft�f3[�rwQ�H2W���Y��]@I ��2-�}��g�@��V���`�U|�:HIxy�/��)®DP�X(g��|�z��,���f<�� ��.��2���F�����MD�Md-���VRɮ�����~'�'��2��Ê`��ԥ��B&�|ݴg�����dP�( /���H����2��1�]`�{ ID^�d<V'�381H߂�Đ��p�TS� ��=�{��#؝_��N�T IY����C"�P7��V�\�7|�2&�"aha���g�ޘ��r*�!W�ql�pݞ����ӊ��V�kR��]דؚ�q�=�����1@:4��Cc���\��e/|���c'O�#��i�f�ICf��A���P��+��`�OM���U������dd��A�����8��.&�p�k��#���,����ŠK�t۽x���wڊ�� �^�Ӆ��q!�in˫�����ĺ�s���0�&�L7��a���<R��u�Xp����:@�o���>���wA��T���N0[���j�1=��x���_H~�c|e�Գ�-3F��������"�9�a���<��4xm~U���j�2pǣAg��X#�r��')�ՆO�G�2�)~�H�Pd��t?�0�P���:6�.n�b����b4�	�f�� ���?�)���,��LM�``�Q4��Hm{��(�A	i��IE�������e�Ձ�Ӌ�ڥk�ܡ�-�$�Η��A_*(P-��@ �	+M&p�b� ����o�M��Tܛ��GR���q�N�R����S1L�t��4���q����H�̋e�B@I����XA�o�Y��(��Fk�'h&ynKЈ�R*/��̺� ��~/�F�I,��ߓ%�^ �����R��ř��Qlp��� !$M�xB���͑&2�n�Z�'�~XL�*��`|��ba�}m��!`KC��~��5�󙟍�Av<|k\O����Uv>w*ugD8����W����Ŗ�z�,�����qE7;�:*�0�e���aܯ�vh����O�G�+"F��� �-9 �{ER
�Z�d��~\��>�q�3{�*EJh�����VK��Q%�����tD�U�O`�A2B����	|��V�� ���?Sn��l�� j�K>"�؟�.��Q���I�؃Ѳ�@*�]����Ih��k;R�I�ӈ�
���&���B�+E{��lI],P���$d�5յ�̋I$��>u���~�⧃�Rb���l�h3��⸿��[u���eL�;?hn�c���z��� (��&�!�w�	)�#u�13����5oH����&;����O����}c�Y3\uA��b� �����>r�+�a8(ڊ�W�dԭ�8�1#���ܦe�3\��ΈJk����oK�9Ï�vv]Upn ,�t��IV�`�1��bA�p�d�{�Ƨ!�c�� `VtEd�U�*�	fu|������]��{�,+�ǩ��bGz��n|+je��I@�<�E��3�w�w�'����6C�̆d��GE`�:ۚPX��ҵ4��}�l��jk�&�!���_p!��`�7qֲo�ލ�}��
�	[O�>6�R;���������y]�y?�+^wj�E7A@�ߕ�և]���i��t٥��
q�8���{n�xV����cѐ���j��E��X��kь���Q�f���f���&���h���	����T�����2:f:���k��(�^ 
���W~�#tz��[���DSnoK�j��=�AyY�§ݮC���UMD��]<�����.-�1ۥ����+U�n�,�<r�'��F�Dr�GQ����i0��2`�Q�-<.�k�Ꭹ�*�����w2a�Gmg����Z��0���ݧA\��>��x��Ү=\
��k��	)�_���>/4Aw�;=w��ӯ��+)�Q�gU^[+v�L�̬�0�4�\8p~�,8z"v?�uMYV�0X�]x�z,�j���B�>C.�/����:a'vֳ^����$��~�����,��/��O�HKcz�}\��@xM#��ar���j#4���-0ڛ$�9����;v Κ�-�;��j�S
a��KC%�ϻ�4�ݹ�p��`gW�CC�y��otl��@
WIV�7>�Cx�j[�C�D��n(�U3��lP��;�C�A]+<8�P�v���T�w�eH:�A�G��(H�;��Ng��J=� =�%u�|c�m�ޝ�x�2:��bt��3eQ�!P���<J|�X�o�r5{�g-�rS�$���}�\��sISoʧ��s�b4����k�C�r��20��H���DY��q�5�vXz�cL�z<�@yT��x&;nU�K�t����V'e�oG0�j�.%dt�o�&�F��3����F�~��)�l��;�5�,Gn�_I����"ͦ��L���m�S�I!V�Oo��2�u����Fp;�i�u&�cQ�����.��VT�Qm�����zK�n�_�B��,�(1��	��y�5g���X'��̨Tݩ����t�	n
�*��*�����;erOB.'�U��V��pZ܋�:!����7_g��!��p��u0�1g����K{��=iMM�e���}ql�l��{T��9Ɋ���_vt�L�;����(�a��g�|G�L�B�X!g4`9~��u]%���[l<�kb�,7d���K<���n���Լg�@��c�|;7V�IY�]Ȝ}�<�C]��-�(N��$���N���:�]��VE�3���Q�<2�m|6��E��h������`Y�+m��(	���7V���3�C � ?������Ӳ�aA�jt t�]ݝ�b�O�͛x�b�6�R�p��2̰������6���ԡm����!f�`�d$d�|*������m_ܥ�D�A*{cA1K1S�HqI�6"h�R�vx$�D����y��+�1��PF�TJ@�����=��"���ޢwX�����E?�8=�6w�NIS��~�u��VDe�|T��OǑm>Y��dA��-����맮����ȓ�U�W]�����ܒ��ݸ'�0A���I�����j���>��d�ʭy������ɲp�5OUv�&�x9	*��v{t̼�U^���jקּ𵴨����O�x��� Z{��`N�LP��t���)�(��Yo2����nU<,�F㱒GŴ���[�n	�@��Cw��Ԍ�-xrz�����P�T*�������|��JY�y�#Q�Eqll��ϳ��x������r���$c�d'�H\�Y{|�U\|\��#Y���ֈ����)�������+�+wzɼWwu��
��{&���Ŕ%7��3��C{
��,���y�$��ǚ�4JU)�{?�`����%��9)ݝ����R����l��� �a��@��hdY���n�5�X�S���{gVR"#��`��w_�{�7b��p��+��R�<W�IY�����O��o������Cԝ=�m_<�V�Ԩ�`�L��<���~|�>=h��qR^���G���hB^:�p�3��Z%�,�M�`��Ra�'H�����r��>6��4��uv�-vKץ4l�2�ů�ϭ�GN4�'���_SP�����^8���>���^�[���s�Se�8��]!C�Ŗj_ׁ�؊�WOgJ���j7��T�@����Rq�dhƚ 9M�$��F$�{B�_p:t[J.@�P��'���}@���@�ҦI.
m��sE)��ߨ/���ɍ��"&B��[�HH �d���ƨw7�i�n"����ܓ�2�>E�	Ɋ��� �d�K;������Az�aɀ���a�����j��}Y�M��%��_En�Y�Cc�f��C�B���,=�_�5��YA�ɱ*d�����ԍA�2O���z��P\?��P����|ڿW�<��7:�$�E{(o
�E.��5i��wn����p��}���6����<�^�dPt�KmT��)�6Z�j�u��K���p���O�ʁ31�
-H��]�]�`�Կ�H�R���>6��g�#޻��4�OdwBY��-����B����u~��k����������~;� 'z@de��nHM��	�u���:���wl)�ӎߘqS��J��3�]Ts�3����HJ���n�V]��������V�{���nFD�)�ԩ4��?�^�[�� �.Ʃ�*�9��bfTZwLP�oL}F��L�ZB���2���z�g(ځ�S��.[��[��M�&�2������+��Y����T�f�w�+�\���v�6꺺j�����Q�A�J��9���|�N���	����$P�d�W�@꿽� �L�2���W�`3>�SKnY���~Iva�:ގ}�~\�����)� ��e��[0��������xs��w�U����X�1�՛Ƕ��s���_)c���� �"7N���F5.<��u���v��L���>8F����s��� �~�j�S����?���1z8A&�s�nuI�\��_��~���2�5y��Z��6���`��F��-�N�at��P	��2�Ǥ�*v�ow�A* ���D�
��,�NYv�w�]
n���5I���e�ص'w�1�f�ɷb��\�у�R�I�_�yR���!e?ٝ,��Ԕ�:��.���	a�%f�Iej���Ǆ
���U�x��_r�`Z�//���|[�\��sibќ��)�q�ZQ�G��� p�������8S���0�c�pیhq�=]|E�,EW�l�:���#767��������g��Ф��h��Ƈ_�L��Y�?��h��0d��!&�>�ǝg�P�G����V��*2���[�<K_��f��,�p��|k�������Z��GgT鷂���帋k�2���Uw�rl���_@�l'US��P�8.<��O�u
�ح��G�ѣy<��_�ٿ�^����jM���t��F�3?�F�6)$��N6�u�g"�Y(�jF؎9Mw�]�f�J7A��8W���0�+�jt! ?��1=g���f*J6xC����Re��Fx��L'}�1~*є�j��#V��qS	��L�SLWK���Hψt��E��r�����ȟGn��&�4���+���A�<�ޤ3�绮W����<x��w�*�]æ�_�ļ�&�sj'��i�� i�����fE{�JzJ�՟M��T�1�h���z���A�ajDW��Z�2Q���]I����G����l!C��d��ڝ���8O������xH���z��M)�)VXh�دw{�H����v2Ͳ��d9�^sH�|�m1�垔�gl���ݔ��|�����Ey�$P�+�a��/����& �@uRYm~��C��}J�+{5���'�َ�ނxkٽ��[����w��S>��F�i8n���
C�zF��^a�=(30��/��<���Z�@Y691��֓huTT �y�S��I�%��N!�ܴ� �>f��ٕ���6H2�2ri�+�N
^�����U<FȗCL���x��`+H�6��02�7����h��; ]��\;������V@ޱSW%U)��`)�6|^BA�U6SW~`��ӛ\��NE��ɇk̩���� ����=0<���U��}�1^���&^F��+�Ҍ�����a��s��ꙃ� ���t�^��<s�=�8^+\��8[�u�ũ��������O�WTu������n�TZ~�2+M~Y�|"�������}To3^��� �(�MA�|�DU�Rf����6ݑ���!~���{��_��z&��G��(ś�!���L�R�{S�^E#T�^D�5���8'���a��B<��Ny�$D�==�-
��4��=��:[Q�F��ePyC��!p�C3!<�^P�g�	�|���B+�m��{h�1��� |��@Y��=�R�e����;����7`���hz������� ����o�ĐA�!k��g[Gju��	}�,��2�a�6uY�\���w׮��	8�(��f��%��1��۴%�Z�ߨ3�F.{�(��y�6�2��M6MU�-+�̪u��
�(���'7�2DH �	Y/�̴Z�������H�/Z5��?ʚ�oq�+8G�B��"]>j\������?H��r�X�Q��Ģ6V6��k�]]:T'*l��L�qPfS�eH�|di#{�aX�i�~�6&�欸�U���*�I�,�Y�r�}�칉�8AS�&�q�34�?SD�f����� �hg"� G�g�P��F`�1���*� 3�2^�t8����C,��0;���s��Jydu*��ݟX� F���a�KG��_�yW*l�[��� 0KzfL�X>��e�/+���1a�n8�/Be���Eq�M�<L��zU���YNј�D1x:�!g�Y�
�,�#f¢����}M���E�/�ݝ2F����4~��	(��R��@�-$�S)vS�r-�9���o�@�َ��	��BƸ�{�b��w}��n�/Q��Kq�=��h�zu��uh���O`�r����ї�#-�r�����A&��d� s��>�����v����d�a�k�9(���+:���FeRٮ�1'@���0�țPvT��KE��}����o������K�ݧ˞��Zxc������Y9h�xV�]��e�p�����F�a���oT 7߯wN?�9��Y`���rTM����A��C�;���B�}��ҹ����mr�\;�9Xz�zA�s ����ݳ�a�+-�o��"�
���s9r����?���N�5�l�`9���-��ذrw��O`j�5�8�ދXߛ� �<��X3 ,�Ք=y8�"S���ʞv�SX��5��H�m�Fꕲ�{��7X��x37ԕ�SR��%��.`��B� �K[��4�rWz�7z6�.�D��
^m&w�~�h�/Lp,�dm�iA���B j�RM���@�L(B�WkЛ�pD���q>qU��՚0������ԟ�Jo^��o�m\�P���Y�����j��e�����7���}��6�Pf	P��{��sK�H��x����/W*,�הa����is���Н����Bݚ��r������#u|��A�}�{
/���"&6lU�����a�P���&��H���������Q���'���SN�"��.����q��m��T�#,��I��Ο�n��<a��J���(���|yV���N�]�����5�#�dOA���!����<g�������ѣ'Z7�,i���Xb��I�¿g&��(�9�3-�U�<9WA�W��C�el��'p��q�9�������n����ت�xa�]0�T@-6�o\��^�떍C�����y�[��Az:X5�9�?��H)��F�K!G�o���U i��O����S��؊�j�ǈo�9��U�=�;g�,k���!-.�n�F�ϸ��n���)�L1R#k05�L��/o�K̸� 3E(�g*2��*!K^�����J�Wf��|w��M�+�x$J�^��A�J�̼�;$�ث�'�n�n�^��@Z��5N�iT�"�/�����N�'�z��ݹڌU�R��jT�#���e���� q��E\��(�k���;��n���e,h�y��\d�sӎ�T�Mƽ�1��ڕ�Ep��P�=vI�+P�'K߃�J_gD.�ʿ�~1�繇Uu8$e���tV�/��>z�;X�2�ʶ�F���N�αk�G��`��R˜`���OJ����C	���WL�N��̵��l��+�,�k}|p�)��	������L8�R>��r� �,��C��$��6�
�ad��Ht�}KuIw��P�,?Ff�#���Us%�#|���/U��ME��У��Lx�0Ƈ�6�FYȟ�sc���/�W���� �������P�s�8P�|?'�YTj�Ȣ���X9�X*bl��^D�Jao�y�r�����e� y-�B�����d��օ����S�`����9���s�o��#&du�Uh�pP��
�D>W�)t�'��L���R�4��~N1mw����J�*m�[4�.��y�3�X`��>v�Ϫ��f^��P����f�a��l��b'�����'�K�]d����߱�²��8�ыZ��E>���~�"��3����
4�"d1��3��"��ͅ9��X��A�}d�1$�n��N���D�v9�:Ң,��l�vI�1���%�lB�O�~�.�g@>}��t����.��&wP�j���]w�5E(�d�Tvb�
j����(;Y�$8��bJ'�DHW{t�
[xm��x��;39)��/�X��]��,[$$�}�,@�J��lոα�ir'^�f	��Y ��3o��L%���[w?&>��+��9�A��kŐ����!��Z/+O��C]�:�j���y�� \�6�ŝ�cVn^�-�L���^�f(�O�jBQ�@Q�[#���v��h�X%L��Q�"��'}itJ�%B{��g�bI�B����x`�:�T�A���cxh�M��9>$0a���{hꬠG�4�Rް���!��T�
e ������/L0�7�|BՖ9�D��6N����*9! ~�f�:��`b�?J��XU���B��G���f����y��1�0�Zd�	S�4K xQ�5w����6���#����X��azm)�<yI�	U�j��]~�\6]�y���D�%��&�ڪ&^�s�u��(r�x�	rw'`�i����j�
�Us�6��k�
sӝk�G5�ĬkE�Z�Ā�й�/��˦��rhhiy�;Yd�
�^T �v����ɇ�v��q�U�,KY	ݻפg_ �xS����!�8�@Y�2�#�e*�X3F^S%����FP��:��1��/��=L�	L�k�/�$V���LS�T*2�V���:�p�jۢ��N�-_�P�$9��e�D�:�$��7_�\�
���m��R��" �n{��B�r䖜d� w���e�&û��R��-��k���ܱ8��m����2T�SI�>��1۠�<;�y�E�9�̈́�Y�Yp�m?A�mg�������K�t���>W�{��eR��g���}i�5�#ޑv��� ���|�u�em�Rp]���b(���Q�l�T5�>���m��3e��X�d�_�o�/�ȴ�������f�)+�jaRu�y%P����Zъ�h�*��;�Qs&��L6�ŐdKv��
Ǻ)�aK�@�b� ꢲʔ�K�/�4��i�hTP���,8]�~(:_`Gs����q�!&�V�����[I��$�^����Fh&y\WD�e�Nt���������i��$ Po�S@�m��@���qׁ�.����ǔ,8�����'�|�4Sj��K�c��Y�ؠ=a��u��n�a�ar�D���5�U6Ms����i��1��a+�J���d�5�V�̠潜oc��z�,֡�v���||�ra�F��ɢ^�g�`U�K>h��P�h��-
��S�F0:&M�v��R�?�����A$p4K�5��{7"-�QS�q��ŝשc)�c4���n'���h4���_�Ŵ0t�9`Ȉ�AP�����+4<��8E�6Ŷ���y���5�M�.�>壻�c�� NN���
�R"��K3��x����>P5��G�`���T�/�;�Ro�u�@^֣��3��i�l�}����������7��ӟⴭ;�h����?$�\�\'�خ%H.tਸ�58��F�QV� k@e}*��<ز�o+�(�&���:��f�\*UI~�5�4�V8�9&��gT�Hֳ<����y�Oj�9�%�X�����'lH����Z`���'���E��\I����2���8<�szoئ��D�EL@� A^�{Hh�����@zs�)P�� ��7���F�4���%
;9��k9뙆[x)Pa�Rª�$���"��([%��h�~i��˯�O+r�$"�G�E�[�����h*���̶ř�ߚ�^� �G6���}�r{sLϔ���e�(i
�}m9To%H�8�Z�oţ�bL�97���w\E�f`���@Zw\��so��A�ۣ�� 5���S�
@�U��YV�����&CQVZ _ ��3z~�� �q&ک�{����@`��*��B��yi��+� ���I����ͅV3@�B��.:�C~ѸT6�c�5���֊��Dޘ�Mn�2�Jӛ`�'��V�QD$��E��_pq���ʱԍ��U�K*a |�,��0l+jҢ}�t.��P��g���T'Q��i~Vlr��[<�Gy��g<<�j��y����N����V�ٛ����:j�hd�9������~��y�^�S�3���H-lp��`�,P@g��<�'�s
n��N¦/��; \v�.�rՆv]y���zJ�����/�� �9ƅ�2�" n�GB {��,���3� ��F�H�C�p9`� VL����J�l"�������c��L�UP4V�߆��T��Ŗp�����b ����%��m�u!���<�V�UrH+���kd}!g.��	��䬈��C�����uX�i��I�
�HC����E\hpL�2#Ǎ��4�0,g+�v�&ߢc����y�*�z�ls�Ϯ��J�BN	��>/���V5��5ֳ�'�b�,�!Qŗ�~�&�1�Vi~��S:π�_{,� ��c
�!5!O�?��ZA�D���)�����"�掇Ԙ��d�U�:��9�#�$��B3̋I���5�������:���ݹ�=r_ }�3�b4*hS�jT�w��Y�kA��寔���Og~��V�����|���.n��m2(�+��>� ��n��5�W�>&��gD��L����~R�rs����rߩK$��Ң=`,?����s��ů�5�nP�����V/-�:�NY����u�6��γ��\�d9:���)_�>E����}Ա}��/9�s=���}��
w�8��#��W�lŒ��o)��$�zf��[�-��ʇF�^��<'��@�llτ4���*��NI��=qbѴ�f:R<�c	r)p�a��g�U���'�	�e����Тǿ�*�4d �}^�B�~�4���	II�����5�D��S�*������נ\�O���}��>H?�Hrr�"㳀���/���E8�(��]�v Rm���`G3�N��/[A�ə����nI�0ab�A7,���x	=�hS�>Q��C�,:����b�m�=\Y�]A�H;����[�SE���?~Yk[�$k��ƛ��/.6>�B�ŏ	T�Y����`AVp��P?mXu ����	R�c��"� �o�5���n�yz�"��+ÕY�ϬֺHɨf�����\�u���.�.�%����0>W�*�S�-yפQ�|P*[En(k�h���UK�]H����I�˩�Ls92�(��{�� ��[�Q�Uj}L|�����o�/!�3��N�_ɢ"��݁��l�=����^~����$ݢM���n��b�������qJ�=A"5�ɉ�.��u9/�_��ά/�B9����8�52�\k�t���Ly�z�1��y��-j=$�S��7"�s_�x���l�xa��\�D /yp��߷w1wJ��%(�0�u{�U��@'�S��I��R��)Ԭ_���wƆ5����G"�a�O�24L������\H�����T��d��5X �c�3�����xlE*
W���`C�(s��<u=Tt%��i?���>�Lu��H?Rut�������'�$^uu�K-��O8�э����/�)��E�F,�.�Q3z�#s�0�� ܯ�������vp�Q�2�+�Q?�@�A��E�.X�H+���EUO�s�*�D4���u��tnzA����BS�����������c�wɌķ��
�
^5N�̹�(�n��M����e��|�wb��8���[�%d�~1�c�(S�� 7W�HzB}��p�BJz����$�8H}C�y� � ����Q!���4�}�eTd�n����D��=�먓�̺/�K���'�j��"�m�7�����C}�b=����]a����h�E�h��o���w��j�߸>l$�Ϋ5�M��� UÆ��s����*�B7>�}�o�qU�pS	oe���6�ЅxG|IkRs�b��W�G�4�{�����N{b�L�b'�R�Un�[lv��D|3��t%�Q��5���eJ�&v���I�./�;N�N�:J��� �6����Ǧ���^���fm:���}��%��iʹ�!���������	��3�u}ay͌� ���j\�����'�[G:�	Ώ��C��y 8�?��66������<�C��:0�^�
A�;���R�1���E�����om3J��o��a��!��>7V��oQ�����PK��)�oj��PIy�b#T����Z���[j1!=�r�.�J����i���������p�/�� ,fqb��=�(:���#Y.L�<Z��|4Fj[8��(�\��宕	}�Ä��^�]��S��R!��׮�OA|&�^�=�%�ۈக�2ǖ.pl�f�}�ID�E���M$!�7Ӟ1�gl ^�����$ץd@~5�H��E��!'�J��:
���6�����	P�HgJ��Q�F��U���V�f�/d��+qw$8��ql\�Om��v�lvb�:���������ϴÖo�mHD���∥d�b ��-��a�ݻ��io���eF��1�k8�3�ȧ�q _��2i�f��X����.m�!�G�Ԯc�N�'�1�:U��?Y͊ݣ&���I{�f9\=��9�)����r�yl�*��^�Y��/RK(�'�H1����:�ZϮt	���r��[i3���Sv���z�JY��\�	r@��4�� J@8�F���;z���弚�� "��~���(FW�ƛ�8���c���w�ד��c[����B��,G���,؊�8��TUr*>8Nz.����T�p�W�r�������T���cٍ�Xೀ�<*������|;&ahT�"ZY_a%�K�w2���8������-!�(QI_��G��V3	 �
6)�z*�]DOX[����5�yKI��;,��!���3`�̃w��ؕ��%勏��S��(֬���w6y{�[��x�� ��
����tD��q��{ǜj��yn�j@�(0Y΅"���͕������i��aC�$j*�����z"�鰆���.�By$��
�2HP�J��=-2y�:���6���}����<�D��~X �I�`��,��f@��|56D�2ҕ�����@ɊIK�n���CтY�M�67�}�N��q��{Ϭ���;�\�+��ݼ~��S��2-����[ x<���I�hmtvfX6�-�u�9�5+x��dK��fx��N߻���٭7K�������r�[z4��k}QX� 8�g
��lF�6�m��H)��l�wo���΀�xP���i�9�n,�ǤU�F��QFt}/��+��S�%�E/Tu7��a~:�03�#c����e�o�\�9��DWu���d-/�E��킜Ŀ����
��`:o7)��I����0X
����oA�=�MV���]�9��7�R�
RF�菽��-F��[q9畸0��M>#M�k̐���'9%���ү�?*���DC�;�oFro�d
B*E���ŭx��t�rzE�y;J{���i�xz4V�0�*N���4�-�g�Eu3u��n4X�Q�=,�ȅ��/�$�@��`�����R,��x��)�W<���mЅC)�i�:�fsv�#C{��6�QL ~�a�+v�)@.���$�7�I�)n���\��f������9��l_v��p�٦��̱��ȩm.��e�a)�փ�jp5���+w��BL�Ġf�~�0�t1>N�.Z4��,y#u��d�o���\:���!�,�=��tDcA�9
Xv�+�F�+1^��> ��d���jE�
�j�(g���(Oq��jՑ��
#���SpZI*����6^�R�����N&)��a��\ywb��e��J��#�$�w����Fy(�i�/��y�t���7��UIQr=r)F3qHB�^�g�u:FK�$Y���E5��o�31����iO�.y����Oa��� �1M���	o��ݶ�f��X�J����ibS	���DM�8���4%�j,y�Ȋ��`���H��*�Sv)#��p;Un$.���r��m�Į���M'LM���/#N>�i��YVp{X�S��i��[0����s-��$�a�MM�Z5h{�@����=3���v�J�B���4��qY�^&,S����� W��s����Qf�4�*X,	�
0�&��/z<��	<O+^��:L@� �W|��Њ3=���Ex�"� ��O]����TVQ �:�]���P�j6�TL�j�H�WC%�7*�Ȱ��I$.�ڣw�ISCT�X���KO� ���Έ��X/�����T�����:�:k��a����FȂ;�v����?����p���9���\�9�_4)���$&�I���%��|�=X�����ZdV��3>`�X���8�j�jyV^�|Gj+���|��&��I��֛z��Su-��������/��,�ּf�����$�1��R�R~{I	6�3M�t�1Y�Պ2Dte6�/�HE�̖�(�W�A�`w�����暋�o<���ꔿ���9v�.��ي:����b���id��>���p&�B��QA����"��J��#�E�Z�/��:7��tJb��mR��zC�_����@���ׅ���kVZ�G-@�S�����m"�9!/T9wFuV>kN�<�`xOO���^�ᑩ)#��5Ҩ��op0�x�yE#���y�T�߁_��>�㟸��6+���WeU`�?��T"�fW,5z������X�y��ҭD]���&Y^�%D�ҶӦ�ƥ�ߤ��zN�L��(��ӱ����v��(a��۷A{�bM�^Z�V�_|k��q�UBf��$�s,��(�/l����s� I��|�0|��4��P#��6�#�V�?tJL?<ɪLi�U���k��l�Λ��	f������^=:Ī�]B:ʿ���50�����~���6h)ȗ�}]R�)�ž3\�AF�
2��ٛ����xd3�w����e21Qu!��]�����.f�7T�~sb�/Ue�D�#r6�4wo]i������Ԙ16	�#�)�A��*���|)�FP �&�o���c�m�hmLC�4)IF
:D	h@]QN@�N%Y�4�*"�SJ�V#�/k�aѽ�4O��ɐ�������Mi��6Ht�� S.mi��{I������w��ߘݙkչ�9r�j��g�9t���K�Y���7��G�dD�4@v5�����"54���CVNx|u��3��?x��\���aY�3��-�i��?C����A:�@����#���:�__��b�S�m��?��u8l.����(������&�KX�\`����yT�%�:��Y��f�_��C��<�~
7�C��%�Jś�+�.&m��F1�q�锱�D��������1ܝ���Q�i`"�A"��z�F�ݓ{wӈ<|Y�f�����9Y� 5d�Ǳʎ&h�����I����ȎȐ67V8O4�%�|܄M]�Z��YW����]�咄��&�V���x$(q=PuKԬDh}P֫���c��L���˕}���Լ�6o�ﴡf��&�Ő~<(�m�lM�⪷Wp�p��93:�M �����ެp9����o��h~*�,l6g���@���4�
�?�m� �G�V����b!6'Vſ3�b�(A�
�t �� nQ����NI�yzP�4sڟ�.�7�y�C�k�vf"�,9�'\�.H`�y�{����hK?�~�����	�!�Dk@��
z_�F~{�H�܅Gk�G~ki\Ń���y<�%�<M�IZ����S�kbU��I��8���/����KĨSb$��')D����3vW�;W���Z�R�|�>��/�¢c�,!��НD{x�y+c�:�ʕ�_�W5+��A��~��:��{!��U� $n(��Eg���))��4E��q�+�v���p�ѦF�^)0���s��f�2
��\x�RŦ�R�x���Q. o��@IM��+����Cy�ݖA� q���.R���w��]/�"	��$n���"�"�+g(�ԧ�j��H�ܑ��`S3�I��.��s���쎒�i�]m��s��������x*� �t=6�qh���.��C�$��(��S�$ɑ7�Xhb�,�����V��]Ӻ�B�m��~��q[�,��Y�ݦ�u�����}r�
�`cVH��	.!�1���ɍ�����q�,��K�#G��s�1��	���c�0����)N'��c��i��}x�������>(h���(%�f��p�L}`��+x=��+l��^q,��wN��~^��{���	*G�hM8l�vP�jIl�.���r�4�3<��k��pd?J�tYN!�k����XN�?�[�U�g�E6|�]vG$)Ǟ�m�������Ϛuo��b�it5��lX������
�w����8QT�d�h�8���!�Sf�]��I�r)n�A{�<�<e�?�w*R=��XbZ�q���-�%�`���rs�|q~(C��m�z�C���V��'v��E��f&�x�c(�=���>Q\0YY�k/̗7RV�6�!F��U޺p�jt4��'���":�='jf*���R�ܡ ��l��9�Mon�F�a��ӗX�*���4����R�X��A�v��ⲃ��LC�)��Dd2�1�\p��u��SPV�(��bF��g�
����k��ZK.Nw��B��3�4(�)
 g6��yVqA�AC̹y�������ߺ�n�p��9��M�T��c_'�i���fr֏>�g����֑�,��p�Op��$���ȶ��y�u�`�c���hdaw��	b�d,��n���7��D;�kM]Ip���?@�[�8e�o���L U����DLMHR�W[`­��C?��^�C�� ��b��iZo�g��h�;r�^<���C��y�M�������n�"��Q���Hί#A���ť ��;Q˾��94�-��[�yh�8����� �Tm��M����ڷ��V��5-��b�{��{JT��{f�]��*��
z[��K�ٗ)���Ks����@������*`���t�<�<
�-trE3�7�c����� �w�D�����A�ߓ���s6��%���:��;�o˗L� �a@=�$M|�{ �|<�R�\8#	Fw4e�Q2VL�~��7DM9�K�/�A�:w�'�ge46�v���$P�s�u�x�{���JQ�u˵�)׋x0�w\����F�L�(w|H�������k���ܓ���A�� "V5�Z��՞�4pMQ��z�ZZ.3K��2=L�I�g��&d~�J��1WT|�u����(b�f`�]`�NA�>d�}�=g_� '���q����9e<�+�7�k���H��Ui�k�m-�ATT��>I���v�oD�Kc���>XU'� eJ~O`���y'	��u{N2�������c��,���g�m6��c.�WWF��������ۃ%L�1Z�?f�ޝP���������V^U��R�v#z{4����d\�s�/��T�e~�G-�-`�^A!LE�G��"vHF���h�5�v� Y�gƛ-(�=�U4���+�˃/~8X'��ɪe���硅�����i�^�VT�#�
;Ï��,U���@^R�@
tg�3F%M�w�Itb�������J~1�J�)�@Zd�w�ʶ��6��=x�n�̶�q�R��������Ӓ����
�˦<:t;|g���5P��3��Qzλ~ ^ם��zrD�ڭ���~�b<�˜Ԅ��E ������E��Η��A�<uk	���1Āc�2p\/X��5�Ľ�"���o"^�c���O#r�-=_iE|�d:K�&�6�K�iF�1�N�h@��Z����2�yx�Դ�t��VƼu*���w@��,�5������¢�8�ep��Y� D���%eB��G%\��M��%$糀������y-����C{?ȯ�>�J��60�a@�fɵ���!�������%S��9�gh���;�&�CR	��V�b��s\)W;�����F�XD1����
�t��jP�Nᝳ�Ј��c�}�_\7z� �r�BC���*�z5&u���ӣCE����f��ҡ�"R��;}�z��OF�x�ώHu��k����-L�L�rLc��@��ȑR����3�V���!�G�A^vff �G>�oӐt����|> n>�F�H����6��;�����w#,6ɞ���_�� �������Xpנ�b�O��Q9@XҪ�]�B�C�<<��	�4��1��h5�M�8�F��{~:5��=K��칐���+7��{�����E�!��%�S�2D 
�|���Ӫ<:�"tч��3�]#"�ӷ�Ȳs��Q��D�ױQ팗�!l�,[������P}��jL���ΐw�C� ���a�Zp���5F8K%�8\3�K�h�9!"ʭ�Xe�:�?���䁸]���4�du�#tȸ�r=$_md
��6c�x��K��|�N�}n�f��[r$�S��'/rE�:e��9���7����W��Rh���b�'O$��;�
c܆��������G���P���j-'���B���̌p�I@a�z l�&*{ʷ��9
�	A�&�ᑾ&<�1�Q��$n�`05%�]ۘ@�'�?�����C�y�6�dO�<!�%��Hڡ�G���Eߕ��E�hW1�\|�<
WJ�b-	�U}�d��j9;E�Q.i8���3EY���]M69��.�f����B�>'�x�|F�Qk�j��L�Zw��B�w:)A��$�Q�����Y�j��IK�Hc����s4en��X�6���O��j�c画�w+|x�=��J{�>Hf��� fhZ|z��u�W�g�i��5$%?a���I��f�o���_G˅[���B%���&=?=��z��2�r�!;\�/��3�xM�9��ڢ2c��:P��{�LmawKb�z'}�v�d����D?~?4�,�.�J?i�q��G��E,��V6���ex���;�2Xf�����"�6�3�ϐ<m��v�:�(����<=�Ce��m����*�?�Vx�0',!�v��<;i�D����������*tL`��9vg�V���*~Ɛa�g��o(���s���Y�1�ˁ�r��i�,q���Ŭ6Dv}qt��>��R�k�BW9-�i���i�D.)��o���T=���]��E�Q���řٜ�v[d��jRj����	���RJt���*d�'���%KD��*�!{%4?�{� '�q�a�C&?�����L㎟<%�jF�8�<�9B�pt�&}�����s����[;�1��*� �If��^��w0_Z݂K��I�i˭n��$�|_��!���b��Ω�+]��Q�� ��Q۹)�D0h�2��*�2M:m�T�bx�Mi���q��o�cg�"�VG�]
��_�Ů�믒a��|�0�;��������%�}�3�}�쒗��ԡ���%�m�ђ��A6l��V����Cz��.t�����-vue���X�v�� ���~Ϩ�rc\1�u�j��kx���@XP��8vʩ�n\������K7|�O�����l��Z��y�X�R�/G��g[.oӾ�%�������=QFn�h��ڃ[za]�jҡ����m/�E��I� ��]������ ܡJ�F:���#.�	#���7%�����2ֲ��ߕ�� ���N'�47��[��-M�
#�s�Z#u�����a4��ꬸ=�A�A��d��c9��o���S����	v�]������2�6��fK��g���� �;4+�*f�ZO��t�,9"11G�g=��$H�>�gV��6�ؼ'�;�-a�����ɭ���l$�E]+]���^Y�s���AV���G0���1ĠK���ÿ�]��Д��ѥ��l:,����ųE���KT=�K"��^��O��#��`��p�I�sr���L%�N=u%1�F�m0l����v�[�5����0$����l��!�H��L�_J8
���I�0m��)Tl�=.|
�aP�nN�J(�t�R�e��0 ��/YKKĜd��(:f����$�rL�J�أ/�sCS�ՉR&��Id�w�yY$�r�@%*�<1�G���_ �s��!�����`l�a��i/$��)�,U�X����Y6q�����7l��R)ʖ���6���,j��Rw#1�������u�"�	��f����A0�k>8fB/.�IB;�zʇئ��M�)~���Q�a�1�x�_��
���I�q�[j�D���Z<��qpב�A~	h�jA��)��f�amw�vB�dc���s���222	SOOq�l�SO�t5�~`ߵ��b��?Ǩ�+�.U��q�c������](��LƒN�����9*�$V�	3�蜈���G�.�L�u�^�9�ƛ����n
���qEyJD�� ��-��������@��;JƱ��mSlL	b��VI3��� \>�6�ڍ# ��V�O�=�Na]
��|D��6�}��cJ��;���r��*1q��!�p#��oٮ@�	�#�ϟ9�P4��g��r+^��N��YR&?K������A��G��KP�`ʯx�1���k���>�X=O	�L����V�=��*�K�������O>�o��^~��^k�ds�tC���嗶�7a����{�t*�z�Ο�:���No �˻�F~��H�O�'�E�g�,�����.���׆x�}#H���K�"e����V
�9 ]! ��b��m�4Q��7v������ϯ��h�4�9����z��(�]�@����t*@�N�z�Q��g�Y(t���1PU0�,��Xk�>Z�]D�5�����p�g�h�(ѽ1H�ҕT����{Ȏ4��g��bٟ���8H/��N�K�#�I���[d�.$��_w�g�A��@}������+;�o���[��o��br�㐆��n�M�3��� �ޟ=�?�8����t[�#�nl�V�
�2&Z�b��6�x��2�2�����]��35�(5��t�����TA/r}�p,���L�Y�����}���c3�7}ۯ-�03���P��%�g?>��j�&n-���A
7���SY)\�K~���̜�n��1���8ԥP�r������%Ь2E_{u��=}
�n� �G!m��Bs 8e�iQ�ne1� �����r��������Q���ߏ�-i�=qͩ6�B��R��*�X�L���G(���^ٙ*-Z3�B&˲Odj�S'�ǩ�� �c�zU�xH�z2o���6��K!�u2������(I%1��O��x���Ņ�����#�����Y+6l�3�bw���Xc��-!��5��M���`x�6���	Sךx��^>y���7��Y<~�r�_|9�X�c���k�>��>���zv������&PO��9��~��P2�jt��LnK,j_���[$��c�<Y=��?7����+��O��1�ڸ��G��9	4j�A��X��hP���G���ğs�{�����T�4�����������C��a�d�Y����OY�2��"����2O%���K���HsZ��8G�͛�V�f���;�T<�[H�]�����2����^��A�~��M����'�A������h��YJn"�$_���F��q<�g��OwH&b���������r�iX9z,�i��� �l8�	�7F-�)a�8��q�Q?�)C����yJI�HøÖ����q�H�(!˃�,����Jaon�N�!���/*�n����0�0[�J�~�_Mc�Έ����X�����X�ҁ�����P����l��i�Q��������'�i7�m?��]��kw�dأ�sV}�E�4��+��	��w$��٪�Xq��9Di�Uyo�/,�j��&�j���i��q��r�U�O�V�H4�{~Hi���~��os�Ŋ�$�G�`z������D���k^.�"'O��MǾk'��wj\m ���{�p��zv�Աj镔�qQ��e��k��7�r	?M��m�'�����d�RX�]-��5�ꬪN��53D
���i�)gɞ�}���!S[��#Y?0��-H�$�a#�)~�)fB����v���f��]UT) �Ɯ,�C�8�����-Jm�����L�b��<Cw�6L�T����
/�`O�I|���y4q�5
M3)�Olm��my�u}͕���M���
�AOENRW��cF/4aM�:��"�B�2����d���s��&�w�dPY�R��F���&i�K~�z`ҹ���!{�4�ާq��1X���q�,*��r���U7�dlW�>Q���5D讷���'�2)J�&�R:��D]��!P�w�]�,�z��y�2����	�!j�$��~�H�z�ow{6����Jd���m ���O�a���Ї(.�Q�X�����w�⠩i���t_���p-K���=p_]�-���l��ܽ{s�б7'���T�����*w� ���+���F��5nC��%��ǣ��T�0]J�f�d_=���lV�g�%��[�N[H�٫��ɐ3f�^��<P��~�kq9�R@��ؠx7�z]��0%ks������%����/��R�:N�p|υ�T{c��J��@���"�L	�@��Y��/yDef�u%G�l��f- �OMd:C�N��'mC��h�k�/0��g�_�^~����W�x��;��>���Ej�!2�7��nD��9p:�,_߶J⤕�ma[�:�ظ��� �{	C̍�U,x,���\6OHtM��Nq(�U�j��/}m���Fm"kE�Ok�ٞ/�m�g�10���J�$��4�j�3O���E	)������Ȟ�,VE[?$��sh�tR]nNqp�ρU$�2��3,d�h�ױ}�Ch�W+�ӔX(�"�2�L0�8�ԡg��n�[�O�mޅ���n֚
�����/��m�>��P(�#*ll��6fI��R��
d���q\�8�!��p��W�=Dh;F�3�Nv����W�"�6!8���52�����d���gL�Ϲe�)��T��V����J`^��s�Ӳ'�}�=,/7��M��/���qd\�[Ёw��)��"s-��aB�8�