��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|CB��na��ۑ���O꿇���0�)vUn�~�<�{�ߦz����춊0���떒=�]���W���
�7���a�0�Q��s,�4��`���0��I#���;2f��[��9�-����J�D��>hY�����f�3���_4ko�@�%�Ȗf����ĉ�u�(I�=&�A�p�o5B9Q�9��<�U���s���@;��)@�}*���K��@7*��_kg6����"sq�8�p����NGi['0Q4���G%��y�sV�2�.b�
�t>ȇ�·���ЉVm˗�)KVk:��,�܍2lv�b9pU6�u���x"�� �|��d�)�l*%��iV�'zUY
�=�f�����ݔՁ]��a�H���앿�3�aF�`�M�������x
�r�4( +^��rR�^?�J�CS0@OL�kv��eC�s¥��x._��b�u��I�H|l$bS�[l��ۜ���?`�x���׉���Ǿ$*��� �Jp�3�Lpl	X|D�ѣ�D8�Ŝ]�:�$��uf8�3�ɶ`�e�Q�$0ⓕ���s�4�y�U��;Î'NCw�ng�|�a\��������wi�E3��O2���E�S�`��#�'?��ڤ�%�?D��(�BP���~ۄ���m��He�f�x�e�X���^����3�� �.�v]�Tf����^:j���qx�*�`�I���o�� ��G��4eu��,b��Vv�U�>�����4��.�(�,���`�vׇ�X�;���M@��>�ܑ
���7��0#����kSa��-�g]'�����XM /l)>Nf�NF�Ԣ���n2�~�&�Q�T�����ۯ�]��(��:�+���\��5����(���7���c�0y!N�ͤ�Æe�h�+�H��~
���q��8�w$qȖ��� 2H}Y����	K�����d(���XC�=����S�`]�����J��Y8/�&��)�`��|"�<x�0,L����Ȏ��u?���(������7`J�#`�EA���$��҇�2ǳ��,�!?_�S2�凓3?�-�&�#=ê�Bu?��@�~wNg��R6��!�0}I�Xs����E�$�����_mã@�����2Qډ)�X;���oi�_�`�J�T`�1�J�ʪ��{��1�A\1Fy�yo�7T�k�G$)�-����e���ȟ�~7�j?\A�ݳE�[֝���d���z6���������C��� ����'��ؑ��'�}�����,)r�>�i�^�i�i���`��S K|A��ϫsz���Fp_\1���1ݑ��)�ؽ�����h2`V䙲g�m�%��CȘ���~�J>v�\P�ê-C�z�$�NbI=����a��h����M^��G�O8��nW�Y���]1����d�~M3����v��uPIZ��LUUr�ӫpݥ3.Dg�yQo��Q,tpfSr����K��Ʒə?z%D�57xA\WC�|?����O�ΐ^O�u�!�ø]��[�Q�L3��0�D�q�U(:�n�,�V�XӾ�=���MK
aL�l�Ud�&� BB�f�qa�[�Ɨ �S����8��������.���Ͷ�&'���񼋾�W��=�̢"�Ip:O��
����EK�U�ĭ���9�sZk�����4:���Y�-i��2�by��yi������M��㱧����xv��8�,^U�2�p�V��@�$��>r"���:��Y�� ��Ѳ�#�MAs22h|��=T�l�:�,`~%�of�_p*N���c��?��-o����2�_y��ɏ��hXRQ>��"ܒ��(J����L��r|6��ή�{0���V�r�XPBz�_6Q.*cK��G��P�x�x�+s��$CG@�tz'��qh�1�&S\�F�����O�ф9fאM�/D�Od	�qh}V�^�uJiq?[D�$��%�eu�CO�=�/e�o���w.�?��x>M��$�zInX�tj��H��
ߟ�/�7�����H��\��#��\����5U���S�V��XNׅՓj�ٱ~�z�7��ƲZ���,V��{�J|�۾�;-��6��������yr��M�^���aj�ً�k�L����n����bv|vpO��3�gyP�L��@qE����2�B�0���~�*�0���u�Â��oe�{�q�����9�EGu�T~�\>�k��
A��_-<�Vf�ݴ�"�<5�w�ƚ3i6�X)��E�����VO�	ӆaX xX �ظ%j�(w�*�id�^�x����Fw�|c��{mQϣ��q���-)��#G��PP]<�C�C�T���@����̣��X���°sq �;�+����9mVQ��B���<�܊�y�]Mn~ߣZ�pur�z=�-`"�:\�e\1)��Sj��S��w�Sᔹ$^�f�̝U��y�'59KEG��,� Ƣ���4ZV�s
�u���zE�}�-���*�)�ҏ$M�R����N����3��*�ϙ�p:�S�%��\P`y���#��Ř��� �|�qv\�P��lUt+��K�3�x\����-.�����4���>�u7�"l��<�Z�*�e�������!T���z�~H�3t
���R	?a������E�C��nP}Wh~���$��D�o�^���fqM�.��O���;�)$���f�/���,����z���Y���ʫ)ԵS ;Sm�c�jr2KkRv�K�yV�]��G��擖s�ú����LZ�8G��?K�m̓�N�.�/�U�5��ظ�������t�/A�	��M �Zô��m�kF�#�TN�7P:�y��]w��-j;�rC��"M�x��o [�a�9!@k���}��S��vt����A��&P�OF�􁱼��q:�"[�n�@Ԍit̫FF�
�]�EC�W>*��
M�{�%�P/�vt�)��]ͳ��:�1�ą�Y*�M�C��TҾT�g��s#���o�|d���{��箕-�s����x�����l� �FxT.��6����+~,��E�	�Zx>�A/�u���&�3��-<s�%ī���u��:�Z�j3瓇�Tn�e��!Nm��y\ϊ�5���f����2���əX�^�ɒ�g���O��o���Ȯw�	����HNGª��4k��׆>�gX�`��/𱁞N�T�|�T���Ԃ���+�&W� u&����N,�@���!������{���^]Q����Hݝe���JtƉ�B��T�Օ��'���8��
WR�]�r�G�D�ܪ���xe��,)�YL���v���O}��/R��_A�#������yK1�\��iRn�m`ߨ���R���N�, `7���1?taX���I��W���錕+����T�>%�p37,���i*�~�9�>�K
�R�����X��.�?�e�F
��ɋJ(�Ā;=P
ӱ���
;��_�Q�*{[u}�Rid߿1�#�Ud�>�ʻ`f2_��l4��0�m�A���{�}������P���X��[�+�_�Y�+-�N�Mg֡���R~��sf�d��=��S׷��ɤ00%~RH�9t�f��у�2`�HѴ���x�9Z�P�c��M����������<7|������ȬJZF��#B��y'rW�c��c

|��/�JJ*	z�����˚0�ǘ�=��oj�k;��.�q5t�4�zj�9:d�P�g�+�V�W7�������cVX�t�g��#��6��!$K�f&��|�$P��J6D/�G����%�rق�2�h	�"h<�q�A"�0-��R�����Z�P���ܜ~FKjO�F]�N����1��F��:�8�w e��4G��,�U����g��mN������%Ii4����ס��E�x����"�Q-�c�iߕH���f�x&|�>>��>�a�OJ+K�l�"��`t�"y�٣�ȟ����ޓ��c�)L􍫽C�ՙ	B���曑���Ë��?��⡳�/��q���N�du��l��p,L>k�6 ?A��^�QC�����'����Ր�8�R��A��=HF�-�F��j<u-�w��,�����6'�^��\y�Ǯ���&����i-ord1�úM6���i������a������C��Mǃ�*��X J�������n@�����9���bH��e�@�<�3���,�Ʊ('�jO"�:N-֬؍�G�U:�F~��g�n-p`��R%m���{��ac��a<M�G�W6�Q�B����B���Ӥ�>��=���J�u����Ų�!�����/gƢ��0�&���Y����3�2�t����
��gsl'5��쪅mݬ���+S��D)UQ�ZM*qHw�ו��p=��E�-����1ش��:�4]�{��[p���JNt_��/_���q�I@Ǧ56K�x*,:���U��]�#����\ K
%Y��~ɼ���	��>��!��~+h[YK��^^�����߈$�>+�"'KH,���G�֫	H�_���+�9�jf�5s��(+��V�Ȭٌ3�>��C��aܩ��g�f��=v�����6ar�T���^�6�N �HM���oB]s�#ݕ$�U�.=�3�q���뺥�K�ٗ�Y�K&�@i�(gc���Ku�T�O07�2���v�U�r�^:Hz�Y0rYW�����D����E�wr��ϔ�}Ԣ�t��s.�rQH���w�a �1E)�K -m䥸���+�3R���"`O[�ٕb�J�G_z�<�L�56��E~�v �S��Ɠ���Ŭًr�+E���,����ǲ�Zlq�"5EX H��B9�_���}UH�6Q����#2��E!�4�M�m�" 2����[�B��6­�"��/����4��������A�~��R8��Y}ͼ�=���ܱ�U@���e�yD(F���$ d˥�M�����=!ѡ� ��	�'�3?g����
aX�.�ں��{�}���O�Ej}���9�C�*��X#������>�9;����S�a(پ	v�1���%�۳i�YifV���G�Ј��t9=}�r�s�9G�7G�Dx�fA�����-Jt[�}�e���<����San����BW	�Fe�2�:>6�e7K���H���M�H�m]��$�t=�^���d��Zab��@_ƓJ����]�����*���nWV�`�b��6%�gmr:i�g"�#mQ��@����:�%�ZQ`A٬~�����a�x0���:���ɶTRJKKߣ�N�F6��E���J�������?���#.կ�ޭpZ�C��E�R�d��m&)�~ݮ&S�$,K��xX�D�͕�)R�$rX3�2I��?��甽��@��@C0��|�v��䝧�M��U���ʼ�r[>�x��/�҉>L�g��ob:�̍&�m�vO/��7F�G���JW��%�[�L��w�����[�e�f�Z���uI	�G3�W��4���xJ�z�k.���e]G5�z��oj�zz��b��Nz"�d�=���l�����U�f�u�)5B?|�@˲[Z�Y�����Цu��q�������En�X���^��rw���@��#Oe7#o+���~�
ϫ�K�5����}kIHyś���A+d�K�,��~�i+ `�8���� ����\�M�,�A����Q`�������Q��d�CZ� =�ѵ����<���2�����}��i.5�;K�ĮZD�֡`r&U0J��A<C�ң�dzp>���;�:'`�Z�˾~On�?)���I����M.���ԇ����ੈ�S�eC���v!q�����Se�p'!��2�ү�����/(�{+3vɮ�Q)��(֮Ӵ����-a�Qÿg�S���������b�n���w��#y��� ��R�1P3`������!-��Y��!���ɿvf��j�4YC���7"�ԣЦ�ݎ�33���j�g,��Q�[#��_�K�����y>P�k9�A�i�<T�1F���� �dB�����'�4�x�ڝ�~h>���e�\
�n�;�ʯ0�#�7�k��c��-���Lg��S\xy� g��c0B�׮��4o�D1�p��Ŏ�'��Z�G�Z����G����׌v�����Z�3����1��_�}w��UB�%�/{
�;��Ui�Il�O����%4U|JYe>�V`��R���/0B�*�H8ص��bq���C,B�L����<F����� h��P��5m+�)o�G�T�Q��cL���ë�L��({�`�|n��&H懼��h��^T����� <c���X2a�$5�X���{o�Ԩ�4ůU�}�i�*�����rQ�� $A+�ؠ��^�1ؓ�vaNh�(���i{v8��{�nW����#�	\*j�%,D�j&��XIz����.p�+f1�M�wp95Y�����^���4,�𹩡�ɴT�A&�W.����@�]���p'��X�*
�ko?MuJS���w����ɚ�����U��Ʀ!�~����ߟ 1���"z)�O��fٓU��.�����=�C^k1�I���IkU��˓q�r��$�Qn_8'�Df�K��@��ak��8���U����p��N����<�k0��(p2���n�(c�I&��b��+�9-���_�Q��w�Z6k��j�*A�div����6xne�l9�<�JwV_����m;p0�Da��+,�k�o�t+='+m=�6>ʈ�FH���YŠ�bb%@; �4e?]<�jW:���N�}1� �V�ȟr�7ƭ�"�8�2h�N�:C9o顏���������.mϭ�x�C?�Z�`�^ �]��R;���<B�@��iڲ�����ƞ�*��n5���U�Y�t#��hX����(x!�կXza4=^�,<Dk�B����a��\��1�<��t}��E������cq���O�:����[藆��\Z�q[&��]Z�����:��8"3E��a|K�酲tE��g�>�;K�\�E.�~x��l+�<�5A�<$���������s*2#u�Ҡ�K'~��L��kR�����`���<�ý����K��i'⚲����.�:!sر�����r���-�mͺ�i��铞4�r~�"�(5�V��7�s.�;���3�%� g1�Eח�ߣB�L�����f�|�fY�N�����"��*�}s�T	�xBFZ<wiR^�'�����;�O�FfĔ�3��}�AM��x�k�cu��ެ�ݖ�����d��3���L��T�>����}H\I�>#�H�
t{Q:���yu+ף#�x������g��Cm#{G���x3�x�v<�
��r@���1��9ftzp,YJ�
:pf�oz�u=��߮rQ��Aי�&��w����F+U[@n��#���2>�3~rx��t+Hy?�Qx1�
����2�z�H�w��˗�&(���k���q�_x�_��_g{�d8�dhU�i�>�ͥH���12A���69 �QuC�����ِ�����,��>E|���J��l���]?�T�6�(��n�=_n��/E���,/��"�&4MR���?���J4�~��ܱ�$�х\�u��T��W7{|.8�X�0T�%W�H�w}�j`���]�k��)"�G��#�a�bC�E����O�N/P�u.� ��B��)#���8viV��W�N�rz|�:��@�E��a@�~�m/!h��"6xCn��W���KL�dĈ}��R����c��������}C�j1�^��;�?FO��0N�����Q�V]�����U�	%9���9���T`%^ʦ�%��ܫV^�.f���s�@9Љ�X(�N���rsG]+��^�P߿Ԗ��+ţȯe�C%��@Uf�4��nb������@���	ڮ�1:]ёH�ԫrB�A$4/�Т�n�]��v�0���cq��|�m������mQ�D�9���j+�mj������NVY�z�&�������xXh3@�L�@�Ce��h@�-(7�G�Bk��0�Q�X�yw��n�$�?�G��@s�)�7�k�x>gU*ήl{���Jꎆ(����Z�?�U<� ���":R�0T\��;	@O)+q�-d��o����[[��CA�|l�4�=B��)��BN���͞�x��M��#���gJ� �N�2f G�%��z�/s��w�Z,/�ڍ+�;4�1�D�S�c�[r��k(	�������昻Z�kY,�]��b�I�c�Z����/�J����:�b��^f��.�m�7����DT��mAg�H��(��f� �$[ۋ�{)K�G�8�=����[�c ��Ϗ�ކ�,��"R0��o�lC��o�/�2�!�_�ɦ5螝����ݒmD�ޝ�1Q�7�d]S��g�cs����=��'�'�Ʈ�]�ӑOOӆ��ZԓZA�P�d��nR�,��{$k���[�efUasݮv�d�5��f�q�y�lP�<0 Sq����8��d|��nγ��Ţ`�%��v@^X��;����w�W�Z��7����u��x�`O�\��+?U��Z~JM�������n�Ӭ��FVι/�%�ex�
�G��槫).\��|J����F8䂠��,:2�ž��{��^g�FkZ�w��{Ś��*AȀ���JR~�`��i��b�tz���.L��_���.��8�
�=�3VG�,�x/ ��uPR��2�gl&25衸^�:�����v��UT#�	Ew6h5
�������q3����U���U�2��j<ͽ���������O��r����rw����1v��HW��V�e��U�<����9O8v���o-V��į=�i����`:M��Gs�f���W"���J�Jً�V� �p�S��抌+��*�+��N���m\)��SM]�r��!�E0bL10�E�J����� ��B���ˀAڜ{��|��>k�rR����GE)����U)�grZ�Ӧ�E^W=��}|�QԻ��=��5�5"�ʏ����ɟI�#��ŷ�o4�*��:�έ���x���� R[��~^b�G��K��X� "�G�1��y��{�(���Y�g��[ϒ�(FƝ�VY9F࿘���9Gh4
Πb��@�~Z��{M�yW�}MSZ���y@_��ԁ�Z�y�e58 �!6�Z��W�a�*Ļ�O�_{q�k}�U�c��̰D����ci��;�
,w��0���Jj�K��4%��,��UV���z�]���5X�Cع-��-%�愺�0j��6�{
gWOƿ �)���)]V�k�jvc�&#��?�FE��^yp�YwDZ�

gW�It�O[����L��L呺�|��A9�їD��9�F�S��ۍZ��;��r�w�IĔA�3́g�0�����vŗS��3�ذ1*-�rw��D�)5����̀����"�v!����l�����OM��0[���.�c�eٯ��-�xU �hs��5����G��H2$Rcc�%��u;D��侬��Z���k,�Q>�+TsK��H [�����ŋ�����n5���������	���Mc����la�4Z��>e��A�>��t\������`�EV��R��% �RĢ����R��2�+�ӯ wMf�8���֠&R�����G�v��~�W
RҨ����N���.��{O�����D�K�D	�P.��R����d��Uc͆��7����������o��	>�=D�к��=hfa�����Y��8�CN�0`��'m�ˊ��>xnr<<��Zl����������Ҹh8�W�b�^uH�X������ң�����rɮ�Q��@���O:����fϚZ�
�)̛��r]w# s�D�{g�o�)���T�����
�����2����� ���m�����P Cڷ�r��j�cKv���
Ry��9�*�ត����إ� \K� .h�~�(|:1Ëi[�~��O��R]�%I���o�ڞ:������h���&�f���5��[�kA$@��#kZEHGGS�A��: �#�O�R ً,�p�4��h���e��y�@������;T�=��M�i��8��q��.d�4#�)"�Ix�R������^E�a��3~����n�I�9!��O�X�h졫>pܑQB���D�N��p�Ƚ�dظ�i����3�1�����t&j �Bi�RLfb��pI�v�9֪̔���w�����U�P
q���ٸ�]�f�FV��مʝ�p�?�z���ŀ�U���;:�X"�E ���U�0�_�c�'e�:j�"�B��͵3Ԛዲ�X�e�	�p�7�U@y�ƕ� Ɲr��Q��B��N
K\�I�]5��l�X�^�Q��"j	�_y����"G���#koT�y������5����D���
�`"8;��TY�7�brL�eq4/�n7��4�;������*�f'^d<��l�z����[\m�	�q�m���d� :�Z;\��V;s9�؝m/Do]DM+��@E}�
6@=�Z���.�ɪ��ǂ��F��9��� �s�o�+l0�q�o$J'%X�&$g�,ԁT��;��*:5��s!�U��Y9vP��zk�Ihͦ�I�vx@���Q���
��Q�7��BN���������k �1��U�>��>O��-�M���c�&�8�5#ð�`P�YR��k�'��N�֤NTRN����|���cp�-1�s���#�9W�W
�����P��䔘�,��(jha�����P] G7���A�^r�0;���"2���c ���gú{&��h'��[w�!"�#� Х�\�[������dt���ň)�O��:��)�U���(�x ���@E6�C��ц�h��y64l�r�^`��q=�݃Y�
�V�Y e���ct��X�R�K����:a���t}`��MB��P�]4�z�j_p
ro���^_l/��Y��#�}�)�����~;�2���{<� ի:�('i�;�1G~>[��f��i���X��Οi%�EM�/��!�	�5o�73݆vn�>�jO~�����_3�"�m� ��{ՙF}��j�[
�U���X�d!�g�C�� �'iG!��u��Xo%�]V|��J�K�{l������\�/&��!�H������e����A�עb��wO�軫1�j�x���1�����0��[Lrt#7�0g(�CP���@�[���	��d�q�'ϑ�>ڧ�N��$���������U�tM���M�T������c��N��+��ul��іW[д�Wj]J!2���~�^��,��U�����'�4�1#�sKz��L��dI�'EH��F�Fpn��~��m���TުsJ��DQ�,��Ǆrɽԡ,V=g�g�!eX�󲍇�{q�`HOb�G#ìJ�J��({���L�γh�RΥ��P��`��q�8vv�ws��p�כ�5��ݱn.u-���4x1�o�<��IT奉��Y�L�4��{j��Xa�t�1�R��?��~���j�g&f��f��r��Y�P�C��ݰ��)��cyA��.r����{���{
�r<d��Vʯ�F�k|��d�X��!�"�[S8ǉ����R�"|d%�3���q,Q�E� w�FW�J�[����g�!VY�S2����6���V�F��̄,47<ɚL��.�����-.fڶ�uu���բ��s%NFϨ�a���R��3��vM#l���	���@�Q�ؑð�h��(�Ww�
I_oՙDY⧌0ir�N2N/��͓!;�Y'�1���T���y!�/ %�ݐ��Ak^��}�8��%��ԡ��CP��!Ĭ��{�����\N��F�ζ�˔��?SQd�x^� b\f8�e����G�wc!�����)���e���� �^�"Q�;t��P`Vm]�+��J���ؐO���'$��m��S=2|��/�nFi���"���\gx�6��E��&Y�/aɜ�<_�ݭc�n�XS�n[�������^>_�<�Gs��!��}``QW�/qz�6y���=U|�wF��{���BװA�q�xR�i��Ҷ��㚧sJ�f�F�bY���*]�)j�H�RBW�N�)#��>�W�����{OK!0�)��kSY2$6&��jD/����έ��k�24��,(�&�<���)\x�0�����h��J��f��Q��l?�L+�ČG�?�V10.ع���N�&�!յ�L.�
@�;p����V׻�<.A��V��9�j�����١9�ޖ�7��;/���-��U��w�>m��>����6g��WԽ^�(<�-{T=#g�$1'�|v�+?�w�|�7oKTpըQ��u����ݗ;�C��
Fg�Ǒ�?4ÏRۻ�t��^�fl��:�����y�vNHa%��R$n��=����Мj,S���E}E�c��㞚���a���#O6o���%�!�@�K^ٜ{�i�B�c���B7��,I�`]b��U�t�~��ڨAɻ1�y��w��&�,S[S�>�@��B$�[�f�p�c���)_R�%ˎBD[�s1�;�]jxײz�*��<��f���~݁p��J��x4Xu���Tv�6��^���`���mѶhtQ+�&2\bd<�tnK�_��4S�K���}�q`yP��96�Cm�� �_Ϭ�Rە�*�~��>�qYv2�����	�?P��'���YYI�u�U7�ꔯ��?Ǳ�r&�q��!+�#N[��>����%S$HLm���ٚ��D^�vu�_��>���$`�{����k��z��Ҹ�Q�z��/�6w�*�\�g%�А����$%\()6'��U���"0GTIP�{����%ŵT�ɒ|�o�?����&�f��8���4�<�H�o�,Cq�r� �w3!ޞ����"�Ri��h��ǦH�[��ￅ>��7g��톾ǳ���l��6u |�R+��+	�^\��| 5d��0�bw�S�io;&�~a>_�F���j�	G�J� � z�E$��@�����<C��"9]����}�l���>�x����팽�����{0 �v�"���|Ze�GIX�0V���i5�D�\��h
�V�?�-�QM<�pL>͍ٕ|��3nS�1���`��ɠ{(����/� �f��i4��/
�����b��,)X�?mPg�D6�]B'���z�j퓺�+�Bv3��a#��f;��{zr&*�#p���6���|}�*:Sm��`� ���ěNk695� ��M�>�p]��HY�9ʛD����|�L��Ch��!����u8��͚�0+�S��}{pz� ۉ�1}Xj��Ι��n���9�;�����2B8��5zK[�K	��n�P�������mp#�
��TQ���U���*�����fW��U�j���zUͿgj!T�$�XҾ��)�+ڰ.���_�鄷�`�cU�B BL`��jY(�|Gk� �|<�˓B&�=�F�l�&˙�iu���@T�
� �&�g=�=�
Η ٫�r���~5��]�V-55}��>Ҟ��F�u[{ov��=
=�cr�eŇ.�4�����wd#F�EQc�+P�������̮�/,�K	!�'h�����I?�\P%�ޒU7�f�M!�ι�j�Ғ�l2S<J6��s	��b�qp�3Cϴ(<`B������5��sa6����i�/j�����gdbGuݭ����� ��TJ������=d�괏)���8����B$�v�ػ>��Q0D |�TuDy�2�w�
��V�����������BW���ڬ����6��xe�q�{T��E��Y:k;�=ǑqѢ�e"O��#"�@���)Hi~�*R'@3�20�_õ�}j`1�A���1IXK���V�풭�,o�;�!����^e���5�8�ơ�	�����/,,]� �r�9�@d|��ݓ!�gV���S��ۙ;�9>z��Z��£�p��L�y����8#�l���i�#�����v�:,�E ��Iq\&��Lwa|���ѣ0�]A2�=ݧ�74����]�kƥ�$ͺ�ȃ��Ԟ4�4z����qׄ��T��ˀ�w$��K��Y��B����@���� w���yY�[�@�?H���U%�ЕJ�ʄ��1`ꌣD�����<*O�?e����k�
�K.�_~�w�W�e�u�}�؄k<�^6�Ȯş�ƯnFP��#BаA���I�q*w�o�7����٨�it�N�:�=MK ����x���3�2��Tg��]!k�,V��EyE�PG�b���g�I��pO�kE�\'3
����:��П4��h�����T�K"�����T'Ή�Q��>Q���_�����|��͇�k�cr��rЈP����\2����gҾ�hG����\ ,��sN@l#��d)4�#�lL�܍43�n!J�Nim"���l�U1q6�O$a�V�DX�ʤ��M-E��lav5��<�����n���E����ؗ@�P{qG���
8���V<��.��|�w1�UNg�{���D?D��ǎj�ݢ�2f#t3��O���G�����eO�����8(3�S!��8��(�i���>�)wzEjE�J3����nJ,�#�G��+]P��קi�Qc\����W�����,��S�$N.�O^�F��_������3t�h���}�y	Ƚ�1EY��6a=p�.a� ����9�����΢L�F�Y6���sQ�gt*1R?YwN}JoaYb�^���q���5)�q�o)� �B�܀�=���5N�Z���o�2��.��U~�QJZaY6���y��I}�ڈ6B:aO��ir=��//�{�ϭr��g��5����p�JK���1�<���<�9B<�f�b9V��d�-�*͵s�sLM��H�'�ʁZQ�9C���5�g��A=�t�:Gm�V���:�����`���2�R���uc1�w��
���O�fN��}`���=��E7�@C�u��"Z�6���A����|���`^�l�
�p��/���)u��3`�L�U=׶{7�h��R�	F0�P��t�������HW�V��[�
�9x�:bΆp�Ń a�~kA��T)�D�����~T��':���J�Z�Pqi',8��[�2>li�,��;:(L�j:�i�'� jK �k6m��l�8,�y��<.�����G�v�aa�pS�e�@��嘺��6�@�V�>�@]-�h�rq��Sg���}=_&�MN�|yz� ��b#3��1�vyI<�$ż���Fv��aЅ�?:8��k�T)Ź��r�Ǝ� Ru?I͗��k����8F[<S����Η���H�N�2�zp#���t2Z�j�	t��c���*��q�I8S�/��/mD�ܩ�Z,X��છ"��(��J\ɑ�׷ůE�� y
z�b�{RW�3�,�Fr;/��۱z� Q�	����ҁ��oY,��9�ѷ�����o�^��s+DK/�͠�g%��=?ٚ�	�'�Y��Ǖ�y��K5���2���M��+n]͡;+�߬����}8���:��z�B��D7C�EC�l�:®����Ѻ�$�V���-9�^��y����a.�.�p�m�pX7 g���#Br�&��pp��E���7��CW��Ee�@@�D�\�FH����d��`����n.�����]���<;��v�mյ7����4��XP�,�p���@r�{�`��H����'��su��m���ۯP�/<�?���%�@�_8�����3�<)�S/�೎
���k! ո���+=�v�����_� ӷ;�����Ld_��B]KAs�U��ƮJM�K���3��,u��.ϕhK��5�(#�T�����LV	&y,e�x_��'�Vu�pE�ԝ\q_F�x!�<K���.�V�2���)�<�����u_�6<R�>�n?�>�����X,�{n[��~��М<�f_�2Q�(�����D�S�7)1p����q4_@?H���v�!���,�ұS[�;�}��ws���Y�l�������6hS_��ܺ�a������N��x�(�ԀP�
�$��s�:�%U��m���hל6����v��� �$�\.c� ���\��I�k�y8B8����i�G+ם�ǈ���̱������CW鮵Fԕ�0�Lfbiԁ<2��3"TȻ��.��c���i:�!���V>Q6�� .��K*c���!�;�8��Nz�?�3r�w���]�"ί9X�v����WN�����o�� ��}%�	����QSm���]��c�M��ߔ�o���+	kU���ƌ&i-K��O�ݖ�g�Z��ζun�#�Xm&(.@��QT=��o�xp�E�5�� a�����'[#c����j��C�AP�r��:�Q��z��!�i(�"��o�"�M;��_}U����7��=H�)��^{��*O`��UJ.7��OY'��	XؒLCq� ���I[�VN�G���dYQY?��)�i�{0Q#���+�P\
��*�w�Pd�O�ްH�C���;W�h��b"��JdY�/�k���?�O�8a��V"��@�5Z2���f7u|rPc�aTV+��.�Fż�����r���� }��5�9��$ؗ��>�B�Z4a�p��7�j"�f��SW�|��F(t����E�&��
�R�mDEԳ�J��4�Ss�O����F��7�{�gޢ^�Sx��Ǟ���ً���f��^P���'��q�%X����ŷ�����I5��;� AL�k�[��莄A���f�E �YG�*U|q��?E�!�;�X�\��@C�,f��U������>4L��6���
� 
J�^[��h�Ë��4��/�l�?�Ð�)��={����bv�[@Ш8�������f��ݎq��[t�����P�^u���X��BC<8[g-��߄�i}٤ _;a,�iO4�̪�׍���P�jk�=����D��*�0�K0�]�pn~���Gv�Iu��/du��6�G��֝�NN3��9\r���g��t#��&%��`�-}?�{}0~��ya=�VT���=�`�GLܙc�a�x(bq�w��L,r%�d��+���R�� ��Ş�VY֒#����x���T���,֙��Q�<9�LÖ&�U�ݽ���E݈���P���+�H̪i��S�s�!��縍�1���>H�7i@J�8~@k�75�օ�| z!��z�s�ӹ�6���CH�F���2��$���h/�]l<�ʚ�_�*%}������Yf��(h��z�<��fժ_�FrfS�e�
�`�W2|�{
1`,uߚ�$�V .�R�U5����#�k���> ���&q�a �0��g0�(+���$,kBU�*�K��i�{V����O������@�I���ҡB���ow�����[A�����٘�8�l`�ԸC�\�D�L�D=��r����"0nZR�M��>C-φ�pTGf,���Am���f��d���T�F��((��/!=H=M�8V�����y��^�ec\��`r-��)�>}ʫݬvCp�:���(�}
_�^��F�h�j�]|%7�n1��9/>|$���Y´�q�]_{��x"��Vp�͗�2rCg���x8Q 8ZZ����	Es�J��׌�'�Jm����V��}���(C��6�+�Wi�
�QP��/�
>��@P���!� �
��֛��]+�d"4|;j�r[�v/���8�#���8}�̐��}�G��������J_|�EJ3�+�gBDIb7��36a���[B:��	d�G(D���}����h��p2��_`ϸY^Щ҅�G٢��*�� U�r�މ�VV���9�z��ǻ��қ�W�q��؍��ܯFV�mb��߫�$Z�2�>G9XS<Q�^R#����*�_��%��@�<w�ҏ3%d����I� �yK�E��")�(�c�!�F�b-���6�!UK�ȹ����L��!��Y3�\�_#���3���4��g�6aI��u梏�{�ܛ�@z=���C�D��Z8U#���w�`�"0��fA������<f�'���	MO�3��O؃:�8��\W;L�xJ �_��Ĕ�|Mz��l&=��9�ԁ��̦��K���0z��%m�|��'?�O���&籡z:UO<|{�9� ���N�`<P��O��4vH��!����*�� e�����EF���n]��'v���4���@J��bi�н�&b{��-߽60�P���/��wp�A'[�i$��h����rH��5��u�������LҩTN��:h����:�Su���V�J�L�5�#"c	�5����zK��t"v�dI+��*.m���i<�jz�� N�°�Y,�(�q��s�%�%�w�#Ef_H��>uq%��c����������̠"Mv�8m��u>�UW��ē�ΗB��&҃\�J�9aK��!�z��d��6&��a�����W��D��>���͋�*OkV������FI��W�|ޣ6'�XD��Z�%э����䯇��C��{{H[���ֿ�pF"���n�]�R�wB\)氵�:#��ĝp��:fz\�͌t4<�@�D�=��r�,h-8XD�r5P�	.��qT��#��B�A6Ru����á[Q�(eQ���D�!��h����q�	ؾ�rI�G���ފ1�t@���b��;-�9�P�������P�72u/aޖ������b}�������mR�g���P�>|��ڳ�[,��X�\�T�Ʋ��5"	�W�0�;d��v��-����^<~!��s��]�b���٭��/l
��^.z�e�!����#��]�9��i�&��j�=�y����b�-��I~)�M!��m��j��L:��PVE�G��k���a0D�!�9</��A�'�=�%&!qTw>N� HhA��FqG�:	u0�;fV ]��?���>������� G]r,���th�5o��Nce���O����6���)�ݺ+0�B�B��k����ĵ�ߩ}�F&��f%/�چ���Gt1����x�>�`���@.[���H��Ʈ�3`���(�,��;�%���O�y8�#AQ��L�hF�W
$[`�JM���rq����9O�ǟ(���0SQ�̎'U�?,�����n�Ė��x!�y���\��a2@�����x[�l�6a���@�o�!-`1�3�f6iU8\G�'22��́��C��Ԗ�#�f�1b	﷐6@�)|��P����,���}f�C�-ǐH}�*]�a�c?��l��ɽ�r�32���b�_��GϚ+K�����{���)T�W��o�w�'Yl�dcz�3��������
2H毐+�g�)�\�1�9r���]� ���v����w�l�[���u����s�b喋k�S�w�3�e��ҫG�-IB� -������]�G|w�l�-��I�^GF����8H��[0���,8�V���1�}s>�������g�^_�.�ug/,S��,jth��b (WU�m�<w�I0���r,�R6�����/��4�"ya�Z�鴟���C��s�Ї�WRlJ�ݞ�)�ߺ�b?� �=#gu�'M/E�3jѳXVe�;��N̻}W_�wW�62�q����e�+���y��v^g\s�!L�4YQFf*ċꑸ��s���P��J���#�)b��L��������%�~3S�T� ����0�x6�:͜�I��ߩ���+"����%Y&Q%WNನ�+�OSt2�_�����[E�p��b��#�N�dh-:>mԳ��������gcW��lSu� bW���"���;�®���;�a���E�Z��ǕX�)�~
`���W�M��:�(lA�w�}Ӳ���Pn�Ѹ!��a�[/�Yx����P�	�ۓ��=��A�7`�c�¶�Gk��k��+υ�#�`��[�L[�,hlB3�,��zԛ٥A��l3��W��Iֶ�� ��20�hK����ݑ�C��=�_i�-k�䊱{��(<�b߄c��|��=�~��G��)f�z/s��7hy����q�y'���2�1�Z[|/WпTO�d.�'��n��Hn����L�jZ��Q����B@�R��MG���P�@��3��]eBfȍ8�~E��~�s�Ɠ�ק=CD��
���?p̯;��^�>�aR �����BM|:�N6,M5�Dvщ���㮢##$������d:��\�J9`��W�,X�Z	U�4I�,����	�R�J��BӫH)q��u�t�B���,&lϚ���|R���/m���*	�X��&3c�?ht|�iX�MlYC<ox�|�ߒ��ִm���oy����B'Zo��G1H����KI�X��w�ZJ[�����x����6��7��1�FJp�Qr��pD��S���@���W�u�����C!G��g5����� Fub�GD|��S
j䤝�������ut��I���0W^EV~_g}0�zVr�ٱ�I���d�Μ6�����V<��n�N*�	.e3z�MmQ��3sY�	�Z?�i��u�������)i[y��?��B��������� �L�o^Ĵq�VƎ��w����)>9�dIX$�ir.��9{aK���L	�E73h\ecZ&����׆���3�X��[�A�b\~���ŋ�C�L��&c�(n#hP�o�d���X��N��{99I��%E��,��b�[*U�GU)�At��Nj5X�Ȯ�]8<�4%�a��&3ȉHu��]��BW�x��$0��7�-�,'_;3�v�z�щY�\�lcI�*<܌�9��!�D7����]圇�sVɣdgtU�g�$/3ae(�x_������MrQ)Z���˞^���
f�%#��K�"�&��_L�3[y�c�����Ad�,�sY����a��Ttv́d\�:��
I�,���@3�#� ���.gԩS���>.�{̙u�5��W�b�A�*	=蚴+z
/�ZWǯ]*��S��{>ULV�{$���K&�{f�7���$��v��Z�~�Em��`'P��/���k�߮f��վ�7��&� H�z6�X8�r�r,��t����~hS�g?���t�`7��A�V�M��z>?`\ƪ1�M\<?���r	cm���n�ȡ�䮮�q
���1�� <�_�,S^(;L�3&�b�)+���R�����C�ti���(�ɸ`'�3<"�6�h(l�74�yF�P�4
^�"`�.5ں��#WI�_96��5��o�-l����;:N<1���Ju�����Xas����e��[6�_N^�x����|�:���U��|����*| �s�㝽�a z�X�
�ȏː�<b�����Nm�7���h�X>�a�3��r�o�@�1f��[���sp�~ɫhr�:o��;Jl����n�[�߹$^D���v �t[|_�HE�}�8��A��g��^0���S\y%�G�R ��d ��~@{oA�3�9BRh��H���⦱����1�{�[珥��Y�(�Sf*c��q�Rz��%�,�t[A�H�����WI��0R�9�=4����Bɔ)れc��Yu�?Pa�3��N54S�G,�Ҽ�����j�Z���
�j�sq�&��CQ}�Pa�d%@w�M�"�B�Q6�x�c5���_��o�{�U�ڥ�F��"��B����������/U6�f!ԶΙ��T��3�œKg5s�����a��=�F.}���R�b����XJ)6�2_�#$Vb�3C~*����`�"p,�?g/� �
:sT�|m���RV�)��v����r���u���~�q��T�2�й��i	�}��	$6QH��쓺�~�;H�|\�?P�m�c~ԴN�I=��A�Q�/yX~~A[>�&����J�����9���Gd�Ҵ˴�����
������g��O
C�An޽z�
	t���9f�ϱƑ#�qB1{Z��y'�!\���7X�މ�~ԥ�R۱��������:��3�	^��)d���P���ǥ�����5��I26��7+O�� ,~M�x�D+-��H]�T��c ;��MZ��=��B?�R��.k�K]�Zl�#%V��2E��j]�P��!�M�A��s�[�V�W6�"t�� }f�'h�����Q�d����خ.O�!���_�\��q8o�|��rJ��B*���MJ���������h�{+���>ޣ{��!07M�������w�Q�:��Ĥ}�w`х�%��'�;t�R̺���]���t��7Y\~n�Rn�(q������^KK�?��Y\e&��D�T�ϥ�\5�*5}��%I�3g��Jy�3�R��oS+B[�\� 1vm��ND|Ի��`�@,�EL���>�E�����z���]��҃�[���+)}a��N��n�s�3P�`|A���!��� wD�e{�N�oS�B�ˉ�Kog�E�DQ("����-�_�H���B�6åc���^����.��X���{��;ۯ��ꦐ�+-2������"�w�6�5��C����I��QB{nU�����"�O�����g����@U��R=5��U��|`�_y��rz���j"��a]Dk�B�4�!�|�6��5y�$9�����5�yJ�X�'��)��.p�5M�;Am«���^�G��X�<N��$���LϢ7:�dH�`�M��<U��p��bH��ƶN�/
�����1�u����or��MazI��=�.q�Џ;�8hL����%T'�8k��NZ��A�5k��`a�r-8�Ȫ�84���4&O����s� �Ǔ�:��ɸ{��М���\�4l��ރ������t�rc5|l\�j��H�u�:�g�Dl7P؇~���N��}�w>�#v����e�i�-�ˈR���F���>y�/Sd�`���L�Y�{��_���ǰ�]c���S�bu_E��D�9�2�S�#�k���4Z'��ܔM�CB_o�Γ�$�[���+���zĖ������R󫓷��~ز3I��k��c'����OĆK��U(�6x'��E�ɚ��3�F��y$,+̗��2�̺C�خ�I��:���p��؁����3_/iÈ�M^K���`{5����q��Ѷm�4rDR�4�"7F#&V�w�v꼭�½V
��GXnA��#��k/�����\��f7�^�g�_%C�P��|����9O�C"����*�Fh�+6�P�i �=������~6��V��߆8�>���Ƒ�q����{��^�lj�!<��9a6���P4��~�����̦�$�l��z;�L ��_ ��ҹ�*���&�#�]���@ae�j��*Rձ�a�㨃�U�Qi3P\���+Q�H^Ȥ��һqgT ��<Xu����oۣg�j��/���}��n��v�����nG+}a����s�D|G�)w�ds�I5j��6m�qU4��.:��\���.��S�J�'/�Ɖ�++�|�����M@����H�X������4MZ�v�:�Nk�	�[�aH��g�O�*/�/Zj&j�=��Fmd�\�ߑ����
�H<B-����I�Nw�3�2�'��-g�+
/��Ż�Gdl���eq�$�� IL�`)D�H��S�U �H�˄F�U ��g��X�ɯ-��ࡾ�;�E��e�%���`�n�>�F�kBͬ�E,�at��)ꥹG��Ѻ�u|���I��(z1�dd�m�S��W/4�i2vQM`�+� ���4~�Ü�^���
�N^��D���h�w����璘3.	���JDU�QJ1J	��˕����˴�p�`���r����ҀUiIrU��u� ϰ�x��No?�~ހZ��.�MDZԊjN���m�+z�z<�rܒP�z������`�<]M
�k֠��	jE��nlJO�x<#�ӕX���et]M5�5���6
qk?73��w���Zh�[����Q��=f�ɴ�W6������؀r�@I�w���B��w��U�N]�ɲ1�q�����&�3��6����{	?���P�����*T�2�a�D�Z<�<CT��y�������V��xL�#n���)�1)v��!���+aH��Βa�%  I��ͩ&�U#^��Kw����e����s�ad����ި�	?��O��`k�޲�sa��]: ���g�m)��l�+
S:�cޥe���]�0�_�yn�X��qδ 9q��pօ�`��t`n6��S�bZfr.�5u�@:G^����ܘS�L�]F+P�.�;�+V��W��:�K�8��=�D�#&����a����4���	`g��
J'v�W]Y 6���N���Yu�a��ˇ`"�}�W�#�x�����f��!y!r檬~��*k��j�fl3�n��CN�ݙ�ު�́eW>m��)&)=����{2G�͸g��C�U�>��pR��=���N����-Y���Z�K�oH�^�Ct��6��\�.E���EO�F����^��a�d���L���N�Ip���.[�'�?�unD ьR��}�Ը�|��HT�B�1hѰ䎫I��uu;���P� J&���K�i���1d+���&D+��s)~߂��U.Qs� �զb��`ڱ��&0�q�
9)��G�#�-��'!��j��_#�%	NZ ������ݻ�5d�<��>c�O������=Y�ob������:�uC�5�m�T(G"0X�(�صђ�y��"_���^�Ʒcɦ�*l����"�$�����7�q��u�x�WM�q"ZI��0�x�.F����K����}���fZ��^��W�?aX�L+w��h$:�R%�2�����٠2f���<���Q6FJ?�%��*�a0�vƢ��ftu���D�x�;����6
�΂�?���Jm;��65y�<f~�N#z�/}"�V6�ũ�>��+�h�w����9��z� \�:?�5F��ϟ��C�p���ق��^l'���Z�ga��@2�|��y�����w�,dv��G| TiqVfg��~���]_�ŕ#�ɺ'.(Bە��Fk��y�e�r��XQ�b�(��C8��=�7��d�NТ�\O�CĸڦmlHY�4{�,�j8��У�������5`W�9�~zzc�,y�l�/B��s:-�1��TЙ� y�);��}���}:���@/�����"��e���N>WF�$����/%����&����\<L=n�Q'�_�ZI�d�-�u���,M��yv�ppYj�Fz|*����t�<2�2��g7�k��|��A�~v<�yӐk�,��ľq[�n�2�y>�Y�{��v����V���_4�K�Т�GTo*�c�� �d������Z31�rߙ�E��i�i"���-��@1��)�
U�G�4j)��UJ�4 z����#�k����eG�
4�]�{Be%�s�K�M?v����c��B�J�@�?���!	���@�Wy%������F�:�U(R,�6&h]��oܵ! �6�$�0��M��4���\�^��c��㾂:_��E�R�}!'n�ӧ�F;a��t�l3?e�\���G�h(������8���R5��MK��yX������8��-���y�^>L��|1�W�w���_w��Tfo-�e~������0��dJD��aN@u)jbZ��w�,���\)����ÒM�k�L��SW{����r�ՙ�5T�
/����.�ON�d�2<\6����U��٢ �QU��w�د�nRj���	e#ɀ�A��ExkHÓ��!�p�ϳ��ѡ����;�{��SC�	����*�4�1�����M˴=[\���% �b����>� ���� w��w�ɽT22R��9۔��٬cO�� ��S���%Gre#zUs���Ĝׂ<���h0��?�Rk��`:G�Hb�NJDr����9����6A�M������sֲ�0Ș�uT`k�%ˣ���z�"��`���`���
6A�mo��G�Dd�R���,�N�U]P����v�j[֚�Ŝt�+wc�E�ΔP0g�,�n�o^�j�I�w[��]�����E���Zb,��j�����RHCf$���N7��طۖ�Ê~j�����\{�V%J
B_���✭b�����>���ͪ��*7�"G|�H� i�0���J�%jt�jܺ�_]�4�xD�i�Q� Sό�U��Ej���W$�㠨�F@�f����zM;G��%��"���+�KP@c�E�: ���oV`�9m�xtzs#�8����{q͸Yϙ.����gw�`��/��%��_�1���b6p��|e�)6H4"���$�1)�^���N����2��*Ҙ`����*�*��"y����G�Tމ@J&��?E���\P��y��]�QC���Rbr����U6�tt{s}fu�����aG9M��O�L�g������qf�iOO�s���$Ć���U�qDZ�x�4��L�֐���y�oaT��!��
��YYbv`�p0�>�Ϲ,���}���K!��h���+�-G�l���]^c�(YA,3�0=��Z���������!:�r'���LB��;�z��2��B�� 6$Mʖ,�[�Z��{�3gW�g�^��_��Kv~1�ڏ�,�ɸ���|�2���8)lAP��(�w�(WL���f�?�O6�|N�k�0hŢ�p9$q�+G��߽I)��qo+����H��� �L")�j{�@^`M�
�MN!�(K紁.��2*~o���t�°�T-MVD��hd�*���&bƹ�ٰ��$�ؓ���׊\���G�ݨ@$�)���]`vhM��u��u�`R���r�x%d��b>�ӌ�,v�'��c-pm��v b_ae����n���kf�ag6ۡ���LT����&��u@����v���������b��]��Em�]��z��i���p�MAp����;<�3�`�%ِ�̵���?��t�q/կ�d	�;5XBOL"]�Z��|׃?́���;����&���zO��!� ����wBT��O�^���WMx���l-f�/V�ڔ�z�J-�i�+�=�|�^�QX�����n��4��g�hf��2cf�<c��`������i�D���d�-�75�E���YN��d$g �#�4k@�Y� �r��_̕��<�c�bJb��?�o�T��?)�x*�k�N-3y"���p�Ø
./`	<�3�����r�B�Z�l�
 �A��}{Yi�J����Ă˩!�8��cE\N�@�MSKr�"pQ��4⋥b�����PAA}ti?f��k-x1(� ����#;�ߣ� m����d&��SvS�a�}� �GJu<k�ŝ���UV�q+G��TO��}��M�9��ŽE��H�,
�	�'Qw8��,n�8�lW��m�+.��_