��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C{�����\��1���O+��Op�L�2.'�x�a��R;m,�(z���<0����BH��Q{�ـf��y���f�
cx�}�щG�;������:��L��sB��V���[:�~��^\QYK�~�r�b�:Y'��U�r#l�I�5̣((��L?��l�M��\P:��l�k&����6�ķ�QɂVg������PX��G�?�o�bHo����4��e��hr�[������&05��P�K���Xz�S_����	M?ٹg|{��|
��'��<?=b��1%#'�R��J��A�"�~�Gg��4c,����z�}�R�2�8�?��1?N�j2����x�M��v��/��Uet���|-z~п"��$�WI���H���^f��'��������oK��˥��=�[L^��D((�nB�w
[�d� �pX$�H�>s
�ٲ=�w(!�=A����꦳E @Ϭ1�8/]4�Zk�r�c�&�ϱ��E�֚�rÍN��w��~.��|4��aq��L@P�v^�Z���x.]3�`�����6�r�)4��1��#yR%7_�n ���� �BE|�<�/#�vəkg뽑���o?�����T�������S��z��f��k����o�9��|���کĈEiGS\�vt`�a�e��X�NShʼ<��_��&Y��5+D���\�������q4���v�t K!w��;i]�mT-�Vw,�R�i�ON+���$��.�X������ڊ**��͵S�����H��J-��r��fi��>��q��+���k��_C� H9���z��%
�í��z�-�k�ju�ٜto�-Ow�R������ ��Z1͌d}�y�a���Q��w3I[,8����sڝ(+1���9f8�oG��>�j��B��M����a�Zy�������|�z�-��5�S�k]EԽa��_r.&)0w�91E{�nE��f����]W�ֿf|w���[El�g1��N����c��?=Ys>h���V�����op�|����@��J�Ƙ�Q�i����	��ˌ���\��>�L'�vf!�Y�5E +IY��'+�rCn�;���a�3�p�8zD�]�.SF������.��M�Ci��k� �Zf�޶�ec��+\�9���e������4���a6mv�����g =D���a�{~�sL��������S��J&�R��3t��]��'�jG�fRi �Ǟ>�7�8���xHF$����6͞�4���%��0П۱ɞ�y��C$��q5f������e�}}��lk̄ze��.�2��}��3n�X�C|N?@=������ oY�+YɶO�Y��{���ԯ�_&���^,�����h����1����8��D��>�v��d��zKQ1�:��1Dӻ��ԭ�:ng�#ZtJ;Z��O����
����O?F��2cc ��s��s����hD�[�`�j�������#�<UP�+o1��W����ԡ'p������HQ�AкH�ӻS� <̎}�[9��	6�O�خ�]���S.-��3Yx��&v����*M.ʏ�ku�m�y�:�ɢ���F&�P7���1c)Qsb���>Ӷ���Ԃ��Z�hi�E4�ff\z���Β1(���B�VgǨ�ސtZ30.���Yʽ�<|��v�X��1D1��t����lh���9��o�{
��m>��4�g���c�GE-�	Ձ\x_���=�Usּ_݋�_S c����?Z�'��$����1Ү�l/��,��S���Q J���mԞ�$[���X�B�D�,��RB��=e�I�_F�,7�t��M�W�8�k�ykf�[�ek���B���|���y�W�Q��+X����w����ajޣd���5����\�ùW�;�ˤ)>���*��ͻ<�N�u�;���~�P䭩�væW1�i��Gն=��n���@M�}>���h|D�GG$�c�7���~� �
Nb�㣌"`�t_��CG������UgW�z+�#�~)Ao�O�8%�ĺa�ȀJQ櫦��D�_�S�����}!Q	LXsV1=P/�X��I���	�Y�*��c	Յ��&��P^6x�c�5�w���'�LL�R3BC���1����΁ Q$�ir����a�y����1��q� ��#'��S����٤m�,�$ow��I�m���Q��i�
#͟ꦍ�����-�^�O�Γq�G��Y��T�����l�f���எ�kn�$�L�vҜ�\��Q��|���O,Kw�8C�IT�e0�|�J~�2�wLBo�t=�3"QXnK���z\�.���A�2&%�(��hΖI��}�&�/��r������Z��le6��<0eȵ![?2��q׸�>*Te5G�J�8�h-��Q鼂��0���2x����i�^�&���Z����8��9)�Պ +����azS�[Zp���y8;�=ݻ�u)M��rb3��"����³Q�H���fE�z�
-P��$�����'�8�ǉ��*xu��p�Yy�^�)m�Y���ږݕ��ӻxAՎ3�B
�a��bg�}�Sc�Uz)l�BS�K��}�U��c���9v%�`�vz>�׿��rJ��Mʍ���T,׊��̕�z1�����bwV9i�$��i~��G����ӵ�9�f���݅2b��jc<��3��o�!�@��t;zH]����`�-�������:����鄤;/�F�����5�|�:���H�}pG��m]�4�S�y��ё�����H��:�ԫbD�&.s1i#ٝW�8+/k�<�h8{�E�h���E�K�q��"^YI���g����ul7S��7��������Q��g��ʉH �ҩoŏ�U��n5��,0#HG5ޅ�o0V��o�A푢g��w�)J��_/�������B�G�:����	����	,<������I��������p�44[ox���r�9�P�	�y
�iZ��������'�����2��Ӻ�>��5�v�"w4!?^����S���l4�x&6�-^�3F\�}c�uuC�d�:����1u4GKٱn���*�t��ԩ��Hj;�
�[h�V�Oي5��ƒ��ޛ�
H-�\Zo"�E��ݢ��W��ݗp)P�T�&�/*q7)@L\:3��Ib�}�;�y�'�L��%�?��gTo�[�UCr���ߜ�Z��mz����C*�U�`xфbN�v�{��9ǿ�;_r {ʕ$D���֍�e�ud��JP�a�v���i-�
�6ث�n��QX"����H �8���R�i\���3Й��,�9��T�?a9��c�U�r�	Ȝ���CD��/4����;]������bA���/J��2b�U�݆C�kїk�2�_;��2{ҪD+m=��*��{����[�^BD�S�&'Bb�����z�ˀ����ǖ��$�Ni�O�ӡq�i�hti���v�p�1�f �t�'�����3��\���[e���k�AZ��@+d��Y1�US��%�!�eG�K�մ��
r�MK
'��Q�+f�����G�u-�X�i}�]����^�A��J���)��ȵ˽�MAĄ�$�/;Gӡ(i��`/� �=��-:^�q}�|�^�g��m��CEv"#t�鱹.�Ӂ㙗�ĵ�@�n7��|�qL��qp2���e��a`����䕞v9�]���Z+o�G�|�]��mAD{����7�k��г�Ȁ��̤n.��a���D�v>�����Z��? H��<yo_&;�%�K�4�e1�����F����l �M�A:�?R
�;�Y��c��/ꫳeUBO�#x�3����4��/L�n<����ƙk ��[y
�6+2�v}^�$����Lx�Ou�s�b�#Q@�=��O�X##<�0g�ż����r���:夎��.1�v�����DB�74���e7Ţ& ;%ڶ��UΞp͍�󡌅��8��������p�)�^��'�i&�$(0�$�\~r��wӈ�#�e�Ra8hU	��Q+�q�
}#�P�
��y�~�o��7Khc4Ss��@rqck
	b ��5��vW�j�����3��g�M�]{B����5� n:�=%������a.Pւ�G#�v4�ie��8�:ĜV��(eQ�1�UJ�
��<>��7la�t&�j^�6~�� 4uq4L�K\�)x�<b���s���ƿB�*�<�f�\�G��ܧ��("�I�C����=�$�,*[�T�~�;��B�#Z�q�p�$嚨өx~�i��j'���{�zYb0�.x!�� ]���.��� /`���/�,)#�^�C�/!�ok'�Y�`(Je	rTЊ�~s���������N����-�t��	WF;�=��6���ԢA�"�ޥc�0FV�>�{D���6�sP��2;\�z>�2ԗe�]�e�c�,����;�U���@���J�F����IO��m8�9p����:��6.��g<b3	n$����~�`��y���Č�Ј��b��T�Q�U]���rd9���S�^��r����ױW���\`�%�`^�����,�8HP�`vN�nD��C����|�T�<�B�OB�26" c���5���ȁ>�5 ��f��^.���z��!�䬜�&vA2h��}g<�qOW��	0X��5�=]q'�y�IͶwtP��9�dԿ��7�+J��l�aN5h�@�7A�������M�(��WAd��j�((�A�V�/<��V�Zg{Jһ�r\&wi�>+d����yn�p��ǵѵ��+W�)؄�rN4��mbOV�z�*��:�����_�,��u�v�fy���?�ԡ(ۘ*�퇱)S,��`N�;{Y��Y�$,1s���_v�T����	J��N6�ܓg�Sx��U�+R�hFk��^&�
�bH�4t���|Ց:Ni�y�����[x���^IF4,��|�)ԡ�f3i��\dAQ�i���	W�G��/[��R��K6���g�X�_$���hāPpa�����~��� ������d�uۄ��oT4rD�����T�j��ZY���Í[\L\8��}���v�X��,��Z*�X���l\����f�1�zK��V]�ԧ��M�Ȯ�n�p[ph�nLI���9d�%�~�(��kvt��y��XO��2�fhj��sOΕ�>��J� �t���T�ii�m�$^��U��+�ly��qw����O��C��}��X��@%*rU({f�P2ɳ�6o����c�)&jɺ9�U���;��j �X�_Y�G����"���ĝ�4����M돢n㌬�x�k6�D��V>���=	���x@Ѻ��Y �y�hAD~U�Js�e��wD1�M6*x�D¢�XϺ�^9���LXt^���q�ô?��+��B鵑��N�S9����I��]�?B6^�.+,[��
c|��Iͺ��YqdWI�>t�r|�C65H��?c!����I�=��)W�y�k�]�i�zLS��'o/����1���֧$�,�}_}�`�Qv���q�ޕ�!T�ڣ��V'9E��'�$��q�'�AO�%�D$,��h�G��_@�I0S�"ȤB�ˠ�����Yz���yk��7P�T�>��)��m�kΣQ��Y:5p���iL5D0_[���K���Y8H���|�#3^��9լq�C��I	�c@~-��m%��փ�ܲ��ȫc"k"�8�*3�}t%,�[��<�� �P���-��.����H{���W�v��m���$c1|����\挐�O;&C�eߠ��໐�H��iY�X����I���vo�u���cTx%���Y[�&�[�g� �_rV�P�8_WqMw����LRv,g��߹�׸������D���!""ya�2M��jofX��7P��UV��Y�8��(�~A{���� ;����$� ���!�u�٬� %����q������E��{�)���2�\R �ɺ�U=�֐���j����M���@q#�����8��� ���ĀV���#��0�%m�����ѳ.i�h@p`{��b�+�	���
š-����gc��vS!����1�D�#I�_�dFa��8̋"H=Gz����w�T���S�XqP�j�Ԍj�)��{ߌJơ�&����p�TdI]6w#a:��!϶�x�39��r����
�����5���b�~�2w�+�5ɪ{RS�MkW(v爫>����f�a�&�E�ݠ��NX�a��Kx�e��?]B�;M�� V�����X�?P������NJ�#)d��mo7���4���Zg}c5�K	~����N\�b��>pW�����jg���@xA*� _!�<~�����|������}
��W��%�"Ȅ���m�!Q��2���C�y|ڇ�|H#���L{٭���W@E��f ����K�XL(�H�W?V��wd� �<٠� ��6p	1s�nW�������shY���~Գ{̣9rQ�?��a�
���V�����ls>�J��j�8{;E�<(>�b��1��J5���Om[!Ǹ����_>�5�Vh:dZ^(����A/��F> P�A�f����%�8t�Eq��T+t�XPg4�H${�/aI�����1��2��s_������P�.�I[��>+��(7*����ʑ��:�K/:�Tk%��<:�e��ye����]�$�r�����EҌ*u���h�\\2��Jg�v �	�=r��ã���ܐ7<;��a>�}��v8=tg��i���bI+�c�K�G�ߋ����ڤCn{��U��>�X��D"� ��Q��8���n*ÜpӺ�g���(�%�։�a�;:{��%IHӜq�<�	��ʑ~�~�n�9�ecn�A��z����K�c]��h��Ry���O���A���x�AZ7�<����ԡ�[l�7C��l�ȥ�v#Ł>� _.7E@�J�I_)T�[F���Q�P�b���??F�4�����Զ|�u�=Qf��>�������sg��}���?p���%]��!�W�c�>���Z<��'ɣ'�hcn�Ә�����������뮧�qS�uۧF�UiT�.�N���t<�\p��5��$fr�x<�'�ޜ'�Z����.e!��ķ�Zc�4�j)�Ƨ�Sɹ����,��;�H8^�8;�_4F���K'��0�G�2�%Қ5��"]-u4Sh�Ư#����+�ܙ�S�=�_/i�ؠ1��1�}������Mځ�tIˮ{�� ���Ȉ�)�K�~�Ou�;Μ���|����+%��qw)V�8 MJpDy�i��&��(
񘺋��=�zm�r�DΝOULb*�Y��r�V�>?2�^�`ج�g^�R�CC�u�5��]!����u���1ǻg��P��δA-bVW�}چ7������\�A�ɕh.z�&���x�P�yP��^�����I�[�T#���6��ll)�K���u���h�YIp�כ7tR����|�t�)�5���u�6jy�N"�~����⒱��r��� N����yM���a�8�y�9&˩�D-:4�<�e��QyA I��hr���a�D{-�L$�N��t����0��v�E�<�������_v_��v�����u'j��[��]#�bx�H�B`dA��'����Pw����'�]�U4nƋ8����m��H�wt��]ʯ#�
�dP�	�{�׵�M��u��k���3��刌�з�xm_z_q5ti`��n3m�|��|,ץs�m۴��!I�kY�Y��� �Gb���Fx"Ͼ�p)���b^8�[��=[����r�G�Y���w0#�j�Z,[a��zh̏DX�P�^��� ����g�W�_t��J6��.�k+�7�iK��%���R�W��>g���֝���ۦ�n���)���������|�r�P��B����æ���: !�����v�#%@��Bub\P��:�����ۨ���.�
�K}�m�b���%�4i��� Q��:?e��N�2���ܖ>V����7{�4T�����[�,P�7�̪@����K�@P6(W��.�����;:6^D��\�� ,��˰n�qL�}ɬH����6+��
	4�����EHΜ�Z�XK���&��b�
Y[�N	�0�{
-�a�^�pL�(���9B ��H`G�P�%�"�4�ٰOZ'��ڠ_�3�\J��SW[j�P>��?!3ψ7
Z];:8�f��V�𤁏�g���-��<���ǵbW�S�y�5��4�[=�r�GX��r�a��bd�A����%Ѡ� �(s/,5��4%�;.�2�t�����$捻��cL3�6�� K�!a�	��&����U�����oϝ�1�j��JF~���C�޸��6K��q��� c7���������&���)d�(��X�ܞI�zC��|!�q�2�� w��l�D�\gC�����ɐ�9]���r%�Ĺ0Í1��>����J���s�z[Xa�`�c�����bw�h
�����I�v�D������I�g�)��!��t:�w�Ԣ�r���' 2B��ۄ4J��F$�"�IAh-�K�����>tJ�/^p)����t���?�E��q�D��k���֓�v8`���I���"���*�`,��9�E%?0l�Lי:˾��>j���篇n�F4�;\@�pk�C\_V��r|��qmta*$ �t>�~�"�����n�UԔ�_�z��z}(-�M��\����x��.�ֺ� �훝�aj��ŷ�p��V~��ѧ֟O���Pk�=��BVF/m�P;1�z*�\�tg�s�O#����{��F�Sqt��MT7b촣A����ǃ�R���/�W��C��
]�ⴰJ���L�2h��e"Hr?����'S���}C;�B�6su0z���#P�pB[��,N.�̀^��Z�~aF�-�^Q�����d��7ʞs�<���L#��] R��@ll��b���$����s��G�K�X�C�l_+L���C+�z7!x�}$�Tg
��Pޞ|��&3��������EviB|�e^� ����s���an��6%:I�<P0�8�X�בܜ���s���4V9�j��PC%�Bn��:7SnX�Ngf�k4�?E�<"�:#�'ڃ��B�46�D��I8V[����s�R�v�D���a�~8��ųߞ0�yU��#S>.�=�,`���@�wÑ��4C��FY��t	�U�Wٷ�1�M�7��!�V>�X�K�"׵�)�U��܄�X-\�}80��ݒ��L(��e�Z拤> �UC�ӽQuv�6��H� 2*#�ƧL����%�6��~�tuX���w�I8E|f{�b0l^*�"��s��H�zU�h�>��DdT�NL��`E��r�ݠ�r:8��d��z��JI��l*i=⊳�/t;�l�r����ɈPnšKC�]O�[EA�D��-?1F��j��� ��G@��
o�$^����#�=��C�B:�b��y�r�yKN4��a/;-;ʼ/�;bVM.ۂ���ˏߚ/�xp�^[�T�՗C7��[��Y�D�zv E�
���_�)qֈP��`���K3�������Y;�����yPq��==1�^�^f5F��)���,`��O��EQE�-OopÓ}�ۥ�"C�v�����e��I(M�K���ν�mfk�](e�ak����%.Gk�s�E٥ԟ�P�ej�����e�oj�:)�@�
Z`�(��2�=s���ͦV�&��슿�����ƭn#��t�ICK�&��"&<����NAи�D~�\e[e� ����i��/����Or(N�ɗ���
c��}�/L���CY�H�w��;�-`=e�;ch-���f��uph��9^/���Qt8\�F�%�F�& ,v-%�EC�.0h]Δ)ȉM�Ù�Q#���uDF��#g�� 7	�*R?�a��� 4��#��V.;�<��b9�^`h`��
IH�˨*y6p��$��׎C>��4��>��~>jǹ�ѱ��vT1��j�,� ��3�)xF0r��?��P2���t&�o[#ym���p(K�	��H_��V �r�J�$�%;�8�;`�ۼc���k���,2ܸP/_4/N���)�ܓ�@Ѷ����2v~�J�{��%����6�.Ch�W�w-�g�E�ٽ��XC�b#�{�'�VH=Z�g�̾��rC���+ߑ��w�u?w�J;�
7¨>�Y��^���Uqoq�^L�'L�1�Tt8-�g[�("?��'�`k��Y�D��]�
����KϚ���/3V��覎���l��H&�8��9�F=�c9���O��
�p�K'�#�S��#�^�ؖwn����