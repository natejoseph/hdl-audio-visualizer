��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��N(��)�A\ko�}R�����L��k���>��夦�$��Af,爋�s���� ��:�V�͕[ti%�cӪ0�|d�JCHsW.�u'���Pem׍���]W�LH�6�t�$ؑ��ǆ���≐�%�R����U6C�'K�=��Y���k���2Nx�2�����@2�X�AKS: or|�<�wN�Y��M1�O����J��	����\������W4ƕolL貞;� ���hrǓ	���[&xD(R�A�x?�F����kvK{4���}�@�73%����*�Do�&8���%&Y�"9HU�G�L�C%Rr����3/��݅p�����ܭ��Z�W��.�B���+�B.���5H�����v���U2�fW��2�I� �k�k�
�u�w� �d�خ�.�ē����kCCd���%�nJ�9�H�m���AE��������2=�PJ�$-�eH;��c߮��i��q�"/no�B=q��%�<:k,4�ō�'�v򀮚�m�y������4��A[�goz�'�x�6�da��KoX�̶8�߃�	�ȗ��_��Є����<g��=���q����76�B3@��\��͞�x�b�іFȓ:���H�����e���T@���G}�x_�4�k���i�8��\�-�gt(%g�B�ы�qˤWf�������/�&�+��J��Z��xF�����4v�Iuy��gSº��tf�Va���d�z�9�j�n�3Z�ߜ��u��rZ)�nFrA`��3ql�`���
��JF����2�(R4�A���͍D"/�帇��b7��L!`AY�l��=���mSv�­0�q8T-�]�2�������i`|��&���� �~�ֺ��8l��IX���,�v���eO���C�琠���KD��#�/D��($�mb,P��$��>۝�/�����'#B��u���Ԋw]o�"r�3�"���9�0I�0~T��!��Ą�w�<qF�PQ=3�.7Ǜ��E��n���'+�%K����+iT�￠*&�;:�ā�5|�%(����L��.�aO(��_\�c����� �Vm�q�y�atnzFkM��U{�#�"�{�]Կ	�$k.����>�xT�2C��y2�Q�ƺ�� $����#�SI#J�w�b�!l�&��K���j��5��e%���D�3�_�:�r�N�� t�݇��t~���j�.�MN��oTćD��H*~��.��}EBo���!nu0�Q�ɐ
�tN��p�+@����l!$d�8�gs�\딊�o�A@aY��lV�#�7����}��W.��������YOS-�1T��#��>{����~��&*����7S����U9��Å7ڥޏ|G���#�f��$WٵbauP���^?��8������b�-�|�WW���@K��l�*#����JC�	���/6�Ϥ�׆Xby�b�wF�\�x������@� h�b��b�#��ZY	J(�)��?����cB�&��� 1�VőW�]�����u����
�n,�)ͪ(*�

u�8L��M�����`n�lJ�v@�b� V�{���73�QzM����L��z��
d�]�{��}yM��W��I�X��ߨ�{gB�
����7p������AQ�'4�'�LԀ��ZqHv��C�N ����G�KQ��D/� �R��0Y̑#D��!��w$�1&P����Ƒ���#\:��ZO�V`�"U~�� ��G��N�Ay���LI`A�C�����J�e��f{jҋ'R�G�y����L��K1�b0�	���H�9��`*�$���|��Ւ�eB8�f�&3$�8���5a�7��%��D�TT0o�NcsVM0�!�h���ІM��	��n�n�!��Øt/�+lҦ �&��� �JT"�)$]��5
j�5��P8���<8D4�A�!4HX����3N�9�X��q��w�|t�P)�x���v��?Îd������.��~��o�N8s&���K�F���#S��C���qs;A'�hX����q_-�q=��Hնd�>)՚��k3%�>�=����ֳ�}�pGA�;#�&Qك��ME�X�D�E�����H_6̣?3(��uQ�_�ao����,kr��T+�~��.�w���H��
/!D��\�ʂI}��W�rE�B�`�.(�g[�	^�A�;�]S���a[����������lg���ᶕ�p��Ċ<�`Ξ@��98��Z�)�D�e�^F������D3� �&C>�R���yN��:���U���h*QV���h�T#�a�w���f˃�ه
X��F�^R�[E�&�e6	M��������}���Ϭ�[���7-�2y�x��֔�t5\m���@l4boX*`&
v���P�?O�����]��2�CPq�W��h��C��7t�d�����˸��|�&�$u�������;s9�M��Ɇ��%�U���ܶ�b#��\$>D���\����'�����t$£q�AX���H(a��TѶ�Aw�#ڮ�Q<�-�;�v_�z��^�"���s�:�
�:+Е"3;� �<l�^QA�n��i�d�� �Gay��J�S����m�3�ng�&x���RބS1Wf�c-�G�_L�� <�z��%��r�0a&7��;#�lP��0{t���N�������0èɍЕ��`�HjN�R9�c_Al+u45q�E}��Z ��Ԣw�Qs:gF�ȩF��@��"/�D$�7���u<�C-i0����p������z���U��Y���/�ݔ�P�#A���B�����)u �w�.���M�6kI����֧�Y��+n��Jp� �p*�yR�X�Z[_�������Y ��ͺ�� ��K���"r�s���ծ�Ó�ފ9�Bd�:��c6vH_+�,��,*WdTp����Y?�%N#1�]kը_��X�PM
��p�kjn��#%�����\4�kS���FY������3Ǔ�3���1U.+B�my�|��V����z^���W�ԄT����8��9������q����8�R�	�Qx{_1x1?�f���U���+9A�X��O����L4[-��z|b�7�$δ"O��7,�G��Z��	5U�F��"��X�!TC�m�-��b,�\��]�a��Yz2�5�u~���t��#�)u(��5V�Q�
���$n�s���Ś<���9�l�yv�_ŋMiЪ5wƝUf�iST$�(��G���-�7B�[p�g�H��r�(�D`�8;�u25j=X-�_�aU�G�%dL+`l��K x�Kw_�ұ�-���]e4�/f|W�X���}=Ez!������O"d�%��d)%*x����"UJ�a�-J%k��4a$�|���aٟFS����V�I8�����:���[[�7+h��d^8�z�+s��YD�����'�a6���Y�㮵�ڐ"�ͯL�毟~@�y$�"슯��mWx�c����B� -%�9/
�\i@j�Z{6�R�B��_��Aŵ�\ks�[��{H,=��K(#��1�3�r���x���k�(��5�VjE�-�|�H��.g�M�{�R�Ո}C��v��qGQW��~�rb��-�����!Nb�;6#�Q��y�Z+�@�с]��/@̝�'ʯ��K�k�nz��`(���������VX%�ӽ5�=(rg�8�r���je
�m��ج��2̷��mfj&46����/B�h��aq	�h���F
L�`������I�y�W:�Bg�4���)_��i�LT�K���l���m�c)���>�W��n��{�X�!�U�@��Z�qT�T���Z�#�>ѫo�n?�́s��K����ȋ�
��g$b�<#(� O��X
�ra� o����$��!t�G	;�dV�'�4�˳%�p� ��^=}��v��M~�\��_��>H��&8�Z]��$TI����~2�ZgȐ��]�f�}�2I+􋳎�3I�����r�d��.�@��k]�/�,&���r+���Y)M�X6�$x�N�vy�t��2��Z�>g���0R�D�3¼�����"���o�s�h�ޘ��:��>v!'�9V��n��\�pB:��0��-n�<P�:�<YTk��<�Y���;�W�r@"Y]H,�e�8T_o,>a�GF��JZF��:��W�M�Tv�s��%7��r;�7�,�9���D�V�~�F?��q`��>-��)�~���\pg= E٣���9ids��^�����_�`�<�cM��� E����_���b�%����Zgxf���i@��z�@;���]$4��e{��� 0N
�$���T���*w�C����dN�W�u�uM άSZ��I��$28����Wr{���� �(��K��Ν`ŉU)�د8&ͮ@�aLg Cj��~k�I#�BK�`����#�̻��F�S�R�G�"�o<)��Ċ�Z���[�B^�a�TF��00�KM(jS�UaLtO*/z�hu�b��	⽀�\bĔ����'Y�"r��ɧ)A���CH�n[K=��G y5�-e�9���1zKh�ݡ�Y�e�gA)�·sj5�)��>SkJ5���:�P�z�rwP��e����6ǹj#;�
��Zv�9˧�%e��?�����l��9�|�_V�s}�w,H���f`n5���M��E�u�%��։�7-d+���5��c�Kg^��p��p	���y�ʅ�����ǿסt[�}u����}\݌G[+ΟY�����_݄O� E&�����Mf&���IH�Lڂ�$:�����'��,���l���"�4k��N�D��~�"�p!\Z���N�W��_�$#�s����Y	�ޛpJ�1���L$���]��4�1���O�BGC�u��_�<K��G	)n��{\��)��j��U�8�ޗ�u#����\.�F���_l�c%�}i@ԫ��>
��u\r�5�6udB=�à�l��N_��sCb��l���A
�ISٰC��T�%����̼{�Z&9�n���L���a����5š(�~��zraЇ���7�%���喋b
���~2��?o��S~ ��B��I,��#��u������2��ڣ�KMM6*&t�-��p��䵡r�g����E"lvO77�� 0������%���}�5�g��2�#SsU�(d]��p����^�z}v��$���1�]��u��6�i?}yD�w�|�z	����-�T�Ϊɇ��\oF�� ���#Pv�7x}�?�%E��/:�O{�<�NA�{_j�}
Ik\3��h�-����.}���W�f5��.O��>����0����a'���%�j�$�/�->��l�ˬ�i�~��h*@>�[Mpx�irZ%�S�9��+���h?�9_�Ԃ=�Tz9��Չ'�%o	ꆪ,�#�����o%�����J�E��h	Rf�g���X�r)9P!�%�����]��pO��C�j����u���G�S�j6g���n��� �m�?���,�=���H��2�Dݟ�i����/�x�-9��?i�T��3�Ҏ,�����h����8Y� WO�,ѳ�5�R� �Q'.��H���a���4d����Q/=��dI���1��z�^�%%��2v�@��dH�Ň�R��b3-I�Iu��'�	���,�������5 �J�����xg�0�=��|����f��+~p�񜶵�M��q+W-X%�����tp�!�k͏�p��z��T�i�W�_<��y ����=��x�"p�A���w��T5�.O%I�i ���Qi�k���B,Ap6l���w�a�B�#�󷧍�A��7B�5VA[9H,�̩4k8+�v�"ʹ�Ix��~�k��/96����Wy����0����7 0@-�'���He�w!g|��%B5_z+ �/�_��w�_?��LF�¬vE���i�ƕ4ە��c��􃬚���z���S%ޔ˯0K�,���T!iYI.�^d�uc�V�?��K�y��p������%c4:��D��E_̋�던n���V�e;�~��d�=�_}۾�ӹ�*��6��m�\�9P��=!4|S�V_�D�coW�?4Ul �(��SiL��7��N;���g�|�M�m��Qf�ϑ�
��we�]�u��5����t��j�+$����˦� wY>�z�<{�w�M?�����B��������΃�1������^v@bnat0�1�O2䀄��f����R4Ǘ1����%�
�~�]�լ�a�5�T��UZ=@/\���=�� �G��~G%q�{��l��6�4�[�=aV!� �U2��u��P�n�!C��i�;A4j�[�RR�^�3�?��I��[��)���N�e���S$Kɲǲ��SՄ�<<1DY�DHP�(�GM(���#��vE{	��#r�t�T2dkO+^�Z�cP (W�?�%^s\:�.3u�kpCB�L��iJ����y��x�J��	�uӁn�$��}b�fj0��@�Wm ��U��a���c��2�2U�&���v��ާ��]Af$�u�$��2�9�J����_LhQeM��F�Sq���J���X��!������IT�C�D�[i�!�q�x^�mT����8�� �3���M8&�%l?-VKb���d6{�b�r����q��oS�n��,�&͗Q�g,s�G1�u8bX�Z���j�T����t�}~��`�G5�Ҥ�
�!H��&����$��Y&���\w/>� PID	�:z�l
q�.��o��������pr��1wEtZ��A��]��Ģ!qlNg|`m��3�b�N2��� �s����������-�zKZ�c�X���!��e�XD'�i5'Ccd	��Ur��L�lZ�韍�(�~j2af�\�3}������r�s�t�J@�镼o���2���m�@�q+|���.�������+DE+q��gF�_h 7e�# yߡ� ����Fzdf�-�'�N�"r�9� �u�R�6�SQ�� �4�uY>=��dr�K�;el�D����̜��t�J��\��fd�,kD��C��x%Cv �-<�s��Ap�-~cVD�h��\Bz:�v>?<n9:#>׆��G�g����^&(�.�l�u�ҟ�M$����`�`�P-��������Յ	d�0��h�X#��\w�H���g������|[��&�	�E��,}�8�d�»�vN��]ߍezm-�󱀹㊛u����K��_�O��Z��r\�5�Cl!*��@}��^�����A�I�A��?���G�RM���`����7�re�(�����h�Po��P��
������i�QN��؛��{�c_�{z���S�f��>Z�^���"�.Ι2}/s�HxT�{���|" +T} z�l�[�ᠸ+PF��������Q�*��7ءO�T�3i�T���u��b�=�"q	���]��)e�9S�@����|eѰo�U"`�>\�1i�Q�;k�m
����چM�[�'��ل ���u�����KZ�D=�+E�!fT?#RP�g�p�2�AA�`��M��Ʉl\���TP*����@�0�X1ò-���a����{����+͚	A�!x7��h���[3�N!�
on�OR|�B�<����ó�26#�[��	�����lb�D�T��`�8�.�V�����%,�Cv�GEV��hD�?R}9c�(O�f���(ſTO���-���`X���X[_k]��<e����&.�P6)� ��wE�n�{&�
]���\��?���:$���6��U���ȷw���R���Ҩ����d�����>F=%��s�nLd��)(�r��YZi���V&������UGdo�ͩM1M=����J��ʃ$��� W4��� ��a��a���7�vx���m&��+~���z`5`;P�\,�SO3�"�K�}J=�WY�6�l�ח
`#��҇�
�����#&��>c��F~��`���xr�����)V Tz�Hi�e��V�f��4��	��{xݯ��lp'�����Md�N��Bn�J��)H��F���u���MW�ĮY{�[�q2�,�� ���c�>7�T�1iS�.;����|Ź	<�d�#U�'M�����f��Ҍ�\�\�e��<����
f�q�\����`Vl�W{~_.�@�[�u��HzX�p5�9_�\�z�՜�	�0�V�Z������������!IꐊV��� �6.AW�u�!.�K�v��I����@5�y�CB�}�����[F?=�����B�*��d�^&��������
��,���X�����呧��:'��:�.�%�,_�߈���`/ԙa1�k�c�'
����0=:qU=�"_+ ��4x��U ���ރ��@�]>�'�:/b1�#B-�*�t
;�'��T���'�*#8S���5;���&'b�}|?H��̹���Eϭ�@mRI��Շ��x�)$�I��c�C{��{��I�h��X��kEy��!�(m���T �S�I܌I�:$ ���p*����.�BӮF�Q@(l�k�*���i3F��լ�V
k�����L���pq\�,8�sL!�c�:Ed�ܳ*�¿�� J�%���ˈ+B�/�ԧϲ�m��+�
��5=��ZJ�ͽ�¼��,�핬n�a1d=n5��5�Z����N~Ԙl&�p�fI���@���z)oyDC�om@ƻF4�Dט�p�.�B�䌦��΀�g�s���1t^"�=�J"��-ص��N��6y,  ������V!ʃÅ���O�`������hX��NtL^�n�6�9E�6�� *�ی^B�lj�'�P�{��~M\P�$%��&ȍt�%���^���+1�k������]n\{L�mߎN9�Hr�O���5�ci����3��1�33H�͊S���H4�g��M��x�<ڨ"�ִ�G&K$F�PE� fM{H�(������Q�>����r�a��ǭɌ(5�B��"a��V0$7O}ݣ�?���ڸxfV��o`~��:j��E���q��'5BNl�]1����]AR��Sύ{󍸻�{�Y���eKR~��%4�2�k?Q��)Ƚܘ�`����Ȋ�QM�c����6lU��-ף��&8����U^�M\q��V�ܪ3�Ժ�#�~���f�\w]�  -Qַ:��6�PuO��<��@4 0� ��qx5�!��^J��©t=����Xn���m;��+� F3�v��K�@m0�:����� <_�d�](VY�H��F���¦��gX�7�t��aʇ4�j���OZ^ʶ#�ߛf��4�ępR�T���k1�>���X�����Z�{R�n�ٚW�ɂ.�-��_up�Z�>+l��L?��	���g[y�V6��IC��1x[�*�Jn�I��\%C��i��g�R�~�N/��ir����>��e�{!�D����^V	@�?���T}/����W��o�@�o� ��(��=n��K���_��_$b
s���{��/��n�'�e�Ρ}�� �O��b��?U��dJ{�{�-u^�J�<��nNid�7oF�q���)��D޽ަ�V�O��#*�^�����7�^n�xpFϙ��� x�06 v��U�#W@�֝�z���䫈�?yz�a� e0�q��+����I�M��(�;7�� ���+��jզ���f��z��?ɗ�B���\�}�x=����#��x?P�Z_D��޳y��&��g���ʘy,�Jk��K�M�)�bتُZAq���Hd������W�3�	1��?luI<����k2���+�D0��,�9�&_��J�xui����̨V|��k �X��	�N�E7�_�+U.�h&�52"���fw�K���r�4G��|�dff�0KZ��V�rK��oZ'{�9kL�i���=8��r�A�ۨ>�R�G�ဟQ�}��C��Y�Y*�' ���+5�q.	���Wc�o�gI���d&�kz��[�@΁P��c��ЌCa]#tC����~�,jѷS���O	,I�01��[���xÄ&?j��?2�!�xp!��8��U	5����?a�C�鹐hR`�G�Q�zފ�c	�뫃�r����	��*�2�pW��}�h��
A��Ǫ@",���z���X�ON��VMs�(��B�Bڪpu鉨ʱړ��Y��`�����0Ks���Fi��!�b&D���>3N$9�U����gH�տ4c��9ETd�K�p��*�HGX��aX��m�@����7��l�\ �,���@�D��n�Mvq7���xecR��2�㛎�݃�%.�7��������&=�ǅA{.G���9�>�Dƅ�<#_�i)'5�K[�u��/X��O�#����Z��~u�`^\��q�~Bj��鯜Z�S[� �F�D����¬{_2�R�  \Sx��pS�Ț7��c��Sn5�Դ������p؆�����}�ܺ����;	����>��#��G��^˭��q�H)��\����3�3�{{�b��_b�����R�)�r\�/��<���: ��F]�6�~#w�H�k:T쩥crqO��"_Y�	|
��;P/������v.��#�'sH�a���e���e6��ɥ&�Y(�J{o�;㍽�:��Q8�\����-YW��[�:h|�M��Q�:~nJF��R^����î�O�~ȤaV�1���Ck�*e[_�Vm��A1	 ��eq�,�0tΩ�ҕ.	Þֱ�k��!D�,�c���L+�E*�5�x��t����|�(�q�c����!�u��2v��E����tF7�?�xC�MF4�@��|٦ЉA?��b�Ր��	$Q���� �N���xu�ٴߝf�N
�	��!�x���9؅�L�/���I�I��F�h���o
����ʡ���Y�2��/笀G�FSĴJlAO�?	b�s�|WF���q�3���t%kH�K��V��y���q�hZ�,ܚ��l�L"y�/�j F�(�i���Tg�+"Tp��+�uq�����丏�R���d����k�������H&,��R�K�-y�2��=
��6�����Ut��������ԩ�%3��}�ӕQ��u��@_-����^:���{m�|��Z!Ш4�_XLj9�/4���!��*���_����i��G��{��E���yy�ek�W��&�?��|)N�"��P�/y�.5_�β++��3�X	�v���(��y�nG�ղ��'o�i��!�l��eE��Uk��4_��r�{Fe����l�v1�<k��-��0iX
:(+&�&x�b��ܘ������[�wk�md���������9�Z�tų�Lu��s}�|� �H�%�CΗ�y��t��ݿVo�\/J�֨��7�_�E{�qՉ�4YzBs+q!���%�N����`��2�]J
9x�O΍�U��n�VN;D��w���l8e��Q�8-)�e�s�l�����"q8��(���X�D�Bؚwm��ƹ�Ϡ����?f��������[��*R���,c���'e��.4#d6f~ ���߂O=�}��L X��V�X)s(��]�-EG���X��Ё<�Q̜�RlG�r�¢;1kYVS��`WF���͝���;~+��ܺ�կ���n��k=����v!zDA-�7B��G�����@RL�����餞�Xե5y���8z^zSE�
�]�Ń�K2���)Vژ�?<�����At+���eJl�!Oˤ��Nf��R�?�]+LEBps����O)co�b��x�!�5�v8��/$���(q�����E[��\M�#���Q8wuQ��N��n�����Nˠ<�R,>��q�t;���PB{��X����$�Ϳ$J�x���_��/ķ?�R�0B�΀+���X�r��+2���ߏ{\��Ҍ�>��J��>sbyΡ�T�d����Q������o�E���V&��2��h	d�&�O�fwN�V	���u�8��q_S�M����! �XP���Al q��w�v�k.��|D���`�wD��&1�	Ϲ���'�/�;���B�ۈsM��ǝ:{��w���n��U���pr¼6��sL+3�ۚ� �:�:�'`�m|2�'g
]�?6�e��bZ���A��:|�d����{z���f㨶jya�&��O�x�HX_V?
<q�Q1l�3'�n��{������f}Rїǋ'M#�m�`z��0�w��7z�M@6DT\�Z���N��h�
����۽q|�&�IuY�Rzl�'WhS�{N�}9��^z*�����,�P�7�d�����wy�6�DΨ6�`�7Ϻ'Դ���X�$+��ޒ�y�%Ͳo����u�}�=�$�-���.��|�ni/G���1O{>�%��S��l�
-���P�a�d� ,��!-��9���#���H}��]0d��%��8&�-0����E���i%`�cڌ�]�p3�/�V�c����&�B�D�-���CG�!�)b���س��Q�O��bB_�Z%�d����Z/���U����gt�.BZ��ڲ��Y�R
Q���xF ϰ�C�~,�qPZ�79U|�#�w��"�K�h�T��r�0B�g}����B55ˡ)fo#QX�=1���y*W��t�V���X�]R?~��yͼ�
�Am|ђ��g���ʜ��k��y4����������y��Qe-mO����f�jҍ"z� �#������F���Hz�bبP�oyn��蕻VC#*��ċ����G����?<�u������mN�f�;NnC���h�z��J�8��]�����̶��--��Ya\��.$�m ��XŜ�����8�[V#�>]���F���Fb�z�זI]?Oa벧>�@C�U���vuJ����9%��ehj���	��C!#��ږ¤LV�%����/��6-L��ߝ�� �E�]��)��΀�D����8�I�KY�ߝְԬt��ZˣM@�(��ŸT,@SA�� r�Xf�I���F(���$����M
��u���t8"I��M��Fxý�2l�U��\@�M���GXxQ��oE��`��PL9OS2���<�gū�;��NG��ڡ�ZUȩ\��S�j%�Ӱ%��\t⾂��.k&��i�Nܶ8 g�o{a-ǉD���>�ftM0C�Z��c���i8����M�8b$�3�_�ZG0�������	Fȱ␆��%oO��'�h�F�ebd�`X�`}tE�]T�`����D�A+�h��FSy#,sOi��Q<������	�8������L��6NU�Z��l�'g��D�9��P��^k��M5���൉;�X^x�&��K�,�����tWu��Ԥ�~���Z���a���~n�4��Α�7�A�M�Y�2�^��Jh_��|Y�h��S���X�X ���"~��64Dv�ꋱy4�tFT�Bu�շ��;�mgb[�,ك��kQ���H{�2<�03��s>��)o���.x�*[o~�k#��%&텦Q����m�M�P��s�)����<���a����:���8���f9�L���jh����laV�کsD0�U��fQ�/Y������(Y�xy	a���s���Ed"�M��o��A���6'D�o�H�i���ۣ-j�k;	�.�h�ȧ�p�R!���MPw�O��4�Q̌��-���)i�N�����
j�rˋ4�$�[�M�����\x*���F`U�WK�����ř�8��T��sJ���	���4����~�:
�q�1��	�5���6Ws�.��XA�K��;+��F���lu�>C;��y�A�%-����D%`��&+�x�Z�K�p��1��.J�t�A���k5؊^��n��NB�0�FGi�Rm�Nk�����|�i[.|$m;ww�����0��mj)���*l��Ҙ]��k����ԃah����Y�T:�ߗw���I�tHjB�'��N�N���ػ��k�����X���D�h�ыϦ�T;O���a%�1�E���8�b�d���ߌ�s8ь]���l	�d܍y/�V،mD�������rzK�u�Ƴ�	��@,�e��s��	>n�Þ����Ćmr��)UJ&�� �S�^�tl,Y����*�T߭M)�o���Kb8e��	��?�f��`m^~k���:Wݜ�X�u�<�k�T�6�vÈ"u3�P��&
[3�E�/ 3�K���6��B����ye�����>$%Fq�O筫K����u�7���G��(��<w�}��)�&�%#�1>�i`��ɵVz���,7CnG� �ئy�i����+}=n�F�|CD�#҉��I�7��4;�.9�Ls傳1f�E^�:rm�R� .'�fτ1�Ĉ���i9N���o˙I`8H������`!��Fj+���h�4wc �)X�o�?�?�2�2�

�����악*vm�����_�Ptڛ�d�4�?G�
�-�E�U �{�����~x(*:j;������?��Թn"�:�gRn�s�-������o�=�wge��{9�oE�Jo��o��+�������@�~��&� ;���"�hܫ��c��	���,�_���*}J�O����Ӈ��s?[~-������ %0Q۶a�<L+e�]�3J�gB�
�13@
��:�֘����Q��!0α�dlܮ���-I ;�Z�dh�@�;}���uH��F+�lA����1�V�ќ|X�x����w��A� 
OcCZ��3�:��s�1��n?�0���aLZ��dD�SY�N� R��~R�)sk��˩�������y\�1��s�	[�G���̷�gx|�8b��O��H9�Ɣuv����Ih�u'W)FS粵f�<��&V�av(4g�=	���� CXAw�5aʹ�g��'5,�@��=D�.ڜ���9�A���=e���}��i���o��.���+�m�"�4@*l�i��<��vU��P��G�?�9�)�ΰ�x&�uj�
�F��;ɍA��z�($�i�ރ��k��{3�|N�ຖ�D�����Z��%�}��Q�=��[@zT�ОO���$�$�h<E�_�p�~�-��4N�)�7F��4+����i�1b���b8S�G��!l�toMO��iY���'�����KqB�����0\�O@Ą�VH��'���i*�fZB/�M[`���e��u}�����e��n򥬕ub���45K!��	,��fg��p�HU{�#|����w	�.�{:0v���� ���i%�h�
���~
'@"�������=9͗O���pX��Vv���l���FZLK�}�J�pX&�3�*C��o��o���?R1���W����m���5)����H�^R�ܖ�`"e�N�]�P��ĦC��D+�\G�OMBO�x'o����Q`�\����䉷���NN'���T.��Pf�wc.�u�Ң&s­ ��dn�J�X�
5����}^�<�j$�$�O4�s{O�=�/�_����͚k�Yw�nFz
	�1irYȂ��w�y2��NQ�Τ0k�W���geY:�=klX))M���<��u���Ce��jz�:�<��R<�ػ�gȨ�Yİ��T��u���Z]?W2'�Δ�Ow�-�5�K���*�)��~�#A̫j��m��}���C��ю�eJ����<u��%�5��,���c)b`�#O��s�K)���H�IGJ��\HΫ��E��x3�e��,
f�2#[��#�>�v��Sj�~�-bҭn��DI��G2?W��"��C��W۸,�*��;�M�'���U�4�7N��U�t��E��{:�Z������'��	O,U&"*R5c����|�Xض�}g�1(?z��Ι ��?g�D��P�x��%A��PÆ�A�K�Tj�:�Ʀ��Ao�db}=g���(�9+*�Cӯ���Ce�x˾�O�q�/W��F^��\݄��2�.p&ⱻ` �ý�;�Vb#�d��������$m_/��(&�k�x���&�9G��
��Mӯ��0���U���ҳ��X�sBTx'Hs��Rq�oR�mޙ�C�UC� pFٿԌ�\B�]��n�[^=��ɜ2�V�}HKAvԱ�tW"�>_})��!��c���R�h{O��s�դ;�C3V��CPe���	)��.�8r�cH~��KaM.ЭJQ�������L��l��8FK���K�R���y����-?u"�7D�~'�� [a3qD`X�MB�}��:x�m�k'������$�D�u�j��L�8"�8��1�od�&g�g[�w��$s��*�a�@Ck]y�a+㙉_��;v�ѭIT�32��=<����L�聻#l�V k��)'	�DH���^wUַF�zC��T�q?	@\���&	&2�E�������O��Rd����6{�M���<��������us��;����������x��$rX6ٯ���|r�����`�"�S�"и[�$����.R���� �"����� ��7Eh<&8�0�yTɳ�jm�	�N��S�������Jr�15�tt��؃Ѳ��j�!>��0�ϖ�1|%a��T�`A�2�?��AId�Wo��S�P�2��sЖ�����A�h����[����2��\N���M�s/Wmhl�53Neg�G�a>Y�5�R�����8Z5]����R4n��7}��y�Q����Y�܉�w4���mb�.�P�<%06k|gt�Bp��Qo�A�C��c��&l��d�v�{�	��5)`Է*�"(2<�`wt�!%����E� .c�lk�j���c�=��o�SF��D��:7���/tr��x�S |T��\��E����)*�?wG�Cg�1R(��p��MTM\�D��0�@&o�q\��p{o����5;����)�(�t\�Hc�H�	���<��F|-�Z�ᵘ��I�U�"j�iA�xEǙ|Z�#�V5��-�籹VH̸ha9��AGq�F�y���<ŅtF�rj�B
��i$jαb�;Y0n���\ۙnKPn���KE�,�~���ם-pqA��3���լE*�y��þ#d`m_,ƪ�<A��ɌM�ԓ\�0]�J*�L��^���1?:���z��{]FY���{�Š31VI�-��#��D�z�|��=��qVu2Y�S�`�:�:סgS;��nUXe�b���^D����f�o�i����8$?v��[/%�56�����)	R��M��3i�3�yAHچ�F���}�js34����No�ACm{�Т��|ō�z<}ܖ�@���.��F����ꡛ����>ʦ����)ܼ�I������ϝ�tY'�]���Y��4�L4�C�� �6�D�{@�ul�"��W&~[�����a�)�6��>@ƗxVp�B ���g��>'��A+F�C��	�����M�QG����ʍ�4/�%�+T���'�߾Ub��,��/L��wk4�M>�	��`�� �r0��I���t��ܶ���E�J+`��!\q��+��7���k�7&��������m���^)u/Lbo�5�#��%^#��s��aG|#^�'�l/)�I����x���&b��g9B�\�+�G&)�~0��3xTg)�~l4�||_�����r�tk��n��kT�l��Fu1W�;���x�/��	�`~��fʞ�F}��D6�e�P��ݳ��O�sX�W�2u?�%+�]����kM�{�%�F�{Xw�d��Q��\G�ŵ�G�b�(���a� �*�mv�=���L#S3,\��[w�O=H2�ɕ2�y��p��Jm)��`c�z u�[۵tHա���%��ĺ*��a�𒘾��&�v���l�a���R��*|5K��,'�+�%0��M����<8b�m�M�5��u��ޝ4��A����z��q����f$��~�>�.p�5���L%h�"@�QJv����d$�4ҵf|cR�T��
��c��+8N`������`0�z�(\�O sc8��������F�p��]�����8n�8�9�"���(�#A�ͦ	k���'���P��8c��c�h��Z5 ��f^ߏ���,
�5X	��AW{��A{:Ap�4;�8�˒I�	����n� �a�Ƽ����+�� H�[��ˑ��8�.�bfQY���¾I&w�c��Kl�L��؊�К*�߃���A������q!T�s��w���\ҵG&�������ތhԼM�k	��,s}&tsοF�]��с�)�,��iJ+�4��" �'�@`xB<����P	��J!����*.+�&��Ҵ�z�ΉƠ���<��8�ϫl<��98�W�7E{G!�W�_K��R�KRC�DA�6f��ZqT���3�S�.����Y�I����?���$��85D�k^�@<�`��N���u.��21�Z�c��Y=VV�}Į��<�������,��m�MdW^ǻ P��
�_V��iH�ɪE�|2��P�w&�� Ʉ�X���aa��ۚ�={ݦT�(�w?Ź[�1���Sz|l������<��O��^T�X��{�!& Dt�&]΄]���˓Y��lH�Vz������!:P:l��d3X?�e�쬎��nz�y�a�ҫ!�iNDײp�](	L{S�C��*fs�J�A��>�0R�Y#㠗 ��G����f{S�QΛ=����v^U  ��I�s�M�Ӣi�u�n��M�`�~#C�v�J���t�	��Txp��G�l<�zf���[�M�#�&�ˌ�j������P�T�y[�Lp�r\mUU�%���`�t�����l��Q3m�*�LX��?��P#W��oy�7�Nzr��Y�5n���nt/L��x��W"�����ifApT�F�Ejz�L�V�����Ч��g�dń}����Ϗ������?%Mir�W*�cZ��IpU�4�0��.��g�H�}�X:6��h�=���kgu����f�]F��?��5���,�n�We��RRpY�+�p�}��sn�R�3+��߬x�S+@