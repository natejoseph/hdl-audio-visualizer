��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��W��<�֯�M�8]m ��>j<��&j��E�$�Ƨ%��I�vп\��s��k������֟���$�4T�)W��"�W���j�؈A���R�~��0s��R�@��b�2�q%�݀@\��,���Ӵ $b�n	�r����{5_f���A~)V�������c��_�7ҖcIІ��T��7ج#jk.&��� �x�Ï����fnW�r+�:E�X���/^=@���9"x��"'E�^�n=�q	a�3����,���x	4N�|$h�a!�̳�e�Fl&�ޯ���9>g����3|�(�h�j�� �窅��0�oŜ�F���
��HM�V�� ����um�mʚ�WS�KJw���EĤ&�4v��_iϮ�#^AE�}���:�'MYP�d��3�c��p)k@�'�=҄W^̃�m"����τ>�
����
���n2����I�����$�t;1����S�N�1���7&�]�B�����3�a���U�����T�.
R��v�96��EO�snK}�v����"�3�����y'E���䞲��E뾘�}�X�}iL����^s��̤��)���T���t+򧃎Yվ��alm�B����~ctS�i�>*J��dK���z��
�g�=�-ԌuQ���w$zP�[Q�ο�&`��_�7E��)��t%k�S8VM�]Nm�o���?f�����8A �6�^�q��s���ׅZbj[zDd��p�,]���t��FOT�ɔ+�Р.���q]M��Y)���E��^�����tr 2$m�<�Lh�� G�C�d�D���p����-�U�<2C�f��0j�NZ�=92����ZY���!V!X�N}��Ůq�A�U�.�yZ?��0�V�G��	��8�[�� B�9x�MF��W�&U��M�������kq�x8`(1t$+�eh�mh�R��W���G�nmU/J7^B�����h�h;�|�G�RF̓�V�����Cpn����d8�Mi#�ꮪ&�w6�GA`��#�mU�O���!k ���Vs�4�:=M�\"u�,BǓFa�z}��槢 ;7E7z1����������X<��m\:���Z�Ȩ�U�q7�ļXK���V_c̡���+L�i�L$􎤫ܕ�0���\l��h$؏�/�o\=�����tNPPV���Q�aܽ�@�c}�>�nK�s����@��2}���3̳[8���yW�=�b��$�|�F������<-
-�N��b��^읉l�����L�M)�H4ɵd�]��Ä?���a��A|��|Jf��u&P
d>B�V�nA��{L7�2�~�Ǉ�li�G���N�<�n�40+�g�3�=K�P��ˌ��-��F���ky$�]=�H�/�Db9���E�D�fFJa�
I�?n�䎙OT�7�? š��Ϸ<  .O@���'K�9f�Nn�x1�M����A$�ߓ�m�P}B��&��+21+�0_���u`�U\�f�{߫(L�yDȺ^ Y�����h*2�5�}�	��Ψ� �Ţ�k�����`���j��n^���� �z@Ҝ8���43�X��zBJ�J�/��.�txg�0��?��Xw��DH���'�p�n͹Q��,-`uU�/�	�tB��A�hfY c�ث��#���s�Τ��=H��@�r�qĄ�˞:g�`�]�����-#����8�{-hD�B���`b��1\SB�ce�w!��9���AJ�,�"ѹ����E{��`֎��*��d��t��K�xY s�k���r��+�(̫'��=�-�%&S"$��H�>Vv�D��h	�pn�L����S`��ñ��Zf�pX��؞7,�ڛAI9VQv5�_�'�̿�;��(� �]r֝��x R�$�x4Wy����^�l��M�Wu���|pas�HJ�������C
��Y�z��%�3��[�!Š���j�ŀl�-X�!�*B`��#��<�֥�'χ����t��):���C���pNƢC�_�fy�-�� ˆ�HBw!�W)Ǭݳ�������j���<6�vn+��鬒!��o�#�!��3�K�3Ew����Ԗ����IWj�y�ve����\Ms�L�*�Lq����]��&6�ֻJy]���<�&NX�S�g�n���)=	u����_̌�x�eZo��VmDb��{�b��.��,IdMB���5yb5�-�Ns1`,��|��0����\��]�##�8��i��k��%)���ZcE(�ڄ4p-PK�ʅ�>{�6Q.�*0Ϣ�0I�z��}��N�"Z�̆���v�=��-I��X "�]m��!ڐYZx�mep�T�j�k���2��Gh�ʴ�Yw�\�3(sl���^�:[��m��[��"7y����>V�m(n.x�+�܇�6�:��L��y
`��	�S� #|��!7�X�O�p��[��*���]/9�����_`G��E�Z尔�z #��i����,�/͝��3�� "p ���qk,��M1�g>����j,�D�K���w���~�>��
�pX�4^F1�}�E��~I�������2W�E^�g1ZY@����{4���mKB$�e��Mk�,�f͢E�;��0*tuޓD��5J��7�#\�����߸�JꝠ�wUٱ/���\�����Q� �|Čk�@�T��C?��e*�@��"r;{��@l:��D�}�3᜘�� ���'㊯����`��Vg��=�oL���7��A��Õ���}�/��j'�x��C�?�ji�?�5��̢�=���a\*�TR��a�s>�<�D�|�{�D2T��[`%z���#ʄ�A��Z����P�ml	���$�Im-0l�A�GE�n���wr��-�Z�쏁{k���@�ǫ��(BI����QI������E9(����:�pǕ�6��
ag�x/��<�����m�j�t[D�QĎ	n9��X�t,x�z��|�Iܞ��B��c�g��7�l�zs%5�}K�X�y� �`�a')��`�6&��/���L
�>� ��< h�Q���S�Q`�D
- /�!�<dxS�$�p��3P�S���_+q�g3��	�^�_�n{�GJ4߁ZOsn�r��F<H�2�������7;��־�!uF�/�f��䑰@��aw����Aw�.��bC�4�%C��o�ޔ�?�Rk�j���+���Nc{	)��4�l�jؖg������a�d�+
f7A1t5��iV'0]�%
e����ѧ��F�D��_�6
V�a�[�s�T�^ �m=*���&S��^�nF�[�HsH%�GM�|���)���wmb���Ge4(�/c8�nC�gEp,j�@.r����9J�R�b��Y8f�?�h�w��<ۣ[]�W*3ng�JFG"X�I���IK/���{4�}��K(�WJ4K9��^$�`'����o���*�Q���5�ۆ2R^���[y�%��M��M����M�:�EZZP�\��'U���i߄5��J��lv]+���/T�u�T�$L*��k[
D�G�:��S�#�0G��C��&Ϲc���ݞ7߼=*�W��F�kt��>f���JR�x�D
��˖h�A�V��2�E5��I�]zJ�!<��xTx���p	�`��9������D3���p��`��&��^~E<�^'�`	gy��!�4�v��+Ji�E��Rzp��8�CcD�����kƈU1�ڸ������{�~�� ��	>8�\�рQ`-��1������s�p�����CU,���*XT���yFr�4��P0l�t��rkk�'|K��ĕ7D��� ��o۟}�<P�8��b���}��A�~��j�.f��B��F\��/0�Z��47����x��H�5����o�_x�<>^�%��?��$f4�!1řc��7%����%�^r w�E^no�Z�袮c�1N�l6ս۹<��X,tz8��v��ZN�ds̔WSn_>a~���%��C�l��� �o�Id~�y�xs�
��9ΎY�J���'��2�b�!���;h�T�;�Ósd=�j��w���YhJRǻ�4X��������[�,l_���̲@�)d=���A�ه�y8�nmi?А�OR�ꗡ� ޾ha���<Ⱥ���Ѱ2��)�:e9�&3��`�ܑ�ڻ5O�Nn� 3p"8Ȉ�f?)��œ���P��
{�5�Q"6$:�eX�Pn�U�4?�~�dL�Z��*�O� Ő�;ls���x�^�y��F{=���E�Y �y�2
Я��)��k�>-��������Jk�-g���yf#9��u@��Bߡ�%��q�=V]��������)�_0=5򭠪w~�9 �
��oxk��q��.<�&���=!�ۢ�D���Yb���8g�.�b	�����O�S����o(�A=�ң|E%_�ci�q���*=�WS�U�R>���e P���iy$�vL��_#7�uj@
aNy���̈́Ti���Ij�6�`��.�k6��2��>�[ɣ�ϰ�3�b�ԅ�;�?� {�]۾�oUl�@���D$��0��61͒'���4>�թ�>
Gc\>O���{\����!�"ԓd��!���_ffftA-��kh��sؗ'��8�cV!��Cn�?I-�/�SHMc ?�9�R2�o�=n`�s|�/�.�
��m>��i-�5��� �r@V�9�_[�˵�9)��m�X���U��� P�wv`��i�����*z��$�sS>a�Yq`�P�ƃ=&x���RL��{��X~_��uut/�+A���|8m'C�X���4�)vZ�,	�7�k���'�vu�I�,{�R�+ N3o�kJ�Xd���ŧ]�iLⰲ��~��f�
hm�<N,u�K��4��c��@"`X�i��/o��(���}	L���-�of%h>�)(�Սx,�e��\j$#b/��g�	��-G00ޚf�@��H<���q���B��]j=��qk�H�͜��a�Sŷ���|�tB��K�\����$���	ra�M<���>o�X�>�*���]����0�D�0n��������@�����t�'��l�Q�v���exB�̞i��N�����ψߦޒ�qز|����@lWa�)�1��hi�H�x�v[#�p%xi��\����my\����r��I����y�&��Lg}�ɲ-�*��;���Du����#t� `���C�L��S�d���R�l	���� Yĉp�G�I�lu$���X��-Wu����3 �!� }9uZX$�LC>,�ׇ�K�5��#����,��|0����?���"dFR&��㍟p|�hfo�&�VH}(EFE,y�]�j�Kac\켟0~�V���#�� ���:5�H�of���ux
��Ͱ��)6�n��)[��6�wD*���/f�p��m�Ě�3�}$�����U"�Bg��	��#	��Q�5/��E��s)����Η,g�2=|��'�}5�*o�H��FNvKj���%�yù��0�P�I����Q�=�T�	����q����@@��݋��)�C>�@023:�@��Jcۏ�j>�#�Va��h��'�g�6��"z�:�0�zA�X�[�B==S$h�?�t��"�p���m�[reDգ���q<���I�(~��e����Nx~)i�-�Z �)���#���!�U�{�{O�Ԓ��C�qȳ'D��jJ_�S�D��Z�ɬ>J@��^�Ұ�<�`P'�ߕ��w�^vғMRK��y���~����+M�)R��S�gF�c: ��C�_��,l��F���3���_ׅSA"�#L�������xz�c	@��2HUV��#D$�+��֮���T��NGcs.�-��@tu��$O�#Hi��c!)>b�_Z��Z?Ԣ��޹���s�]u���	�6V�H�Hm�a�@�� �MHB1ƙ�]��5�E��+�=3h3�S�K�]���i}&��j-�7�w)�0�4x�PS@��GTN���`�kz��N�ej������GE /B}��5�C�|��6��o�\�&ɓG�Ek�OVB��1<�0��v�lu�t9n]�ΚI��=�� 2����&ZbAn�����"KT���b�3N��xx��%�ܛ�ӼR	q0�G�6�?��\ٗk�ظ0����6E}�%{T��q���eʅ����I��̰E��?4��?����ԋ�$�M����Y�C��Fa-EM�Ar���v�b9�,��#O�goH"��V�е
,9�$��G���`#�.�'j@����\d�Z��*��Th�٪�ڟ	g�H����T�	�-j'���I)`���mk�v��J{�`CB�9M�o�%���<����^�in:��r����R��������b&�`W��7�y���|�l��t٬E%�v(,�rթq�:3S��Jqi{�*�3O�t:�Ϥ9ɚ�2u ����QG���d��3(�FǨ?՜�8�F�]�>��#�tU��X?��`��(��x�ih+#^�,�}�� M^)X8�Y�O#��c*T`����a����W�J��p�~�?Fkt|����m�k�#/{��6�_��D�a���NG$I�?��Te�u�F.'�A?dY�Ѕ=P�c��b����Ž%"�5H]f\S��NF�ѐ
v�Al�
#�n���� � (����Qm�Y����`���#L��<�<����̽�:U�dC�}Y�ҳX�]z���`��܁(�<��9�Ǐ��(�|��ܬ�����>��&��1�ӫ^6`�d��/�;K��lEK2�
B'hB��Su�F��i����8{�ɜU����"��X7���$<G&t{��]�EՅ,]���QV�1eH��N�Y����y���aY�P�%����P׉Vո	�5�]�؎��'9� �Ғg>���sO,�A:%�����.0����>@%Re�tۃ��[ ˍ�L[k��yk��!AA�?*��ȷW�*�HR[4c7��ae���Um�]c����>E`������a�3�ME��eTБw��-��/�8�Ń�(,�܃{~�^�jY�3���D�c?�1�h%"X�[�䂍z�/����v��
 :��E6�:"{%���)���؎� �N� ��O	��P�n��M,��"-s���Cw�?�{Î�֪,�A�m�$~d�d��g�@;�Z��^�����]0�6M��YfAE�?/�F������9e���sXV
��n��Q���{�T�n�nd!�y���W/ غہ�Ɲ���.٦y�^�*��M�c��e�Pr�I�0zI�^:A�˚��?*�]�^����W�ubr��<�Y%�	����m�k,��0R�����揊�X�/�&σ�n�ĉ���
���n@���� ��~- ���4�tc]/���F!u��Ǝdۥ��!
!1\�V�:SY�9�������q`v�zw��-� �$d9���Q����9���ъ%�N�s��r̤_�k0Qt:��k\*�ͨ �����+VD��M~���"5r����[T���g����j�c�W�h۠CҐ��3ˈ��WaK���������4�P����� ��J�4�m�~t�`���h���ԁ*8em�<�Ԃ;�}	@���p�3Y�����Z��5�'.ڪ�:Q�������l�2ĵ�B݌�=�kC���q��>ɍ�5���S!�;�*���V��e�R�xAu�zHCȷ��k�Ə�CN=Q������%\�4��o��-<�|-��0E*]��H��Tl7���cȔ^�u�9h�iՄ*ς��Pk1Y�iE$�=�Cs����P�('N�5(����+��ɮC���V����J�@��Gmr8���6n�� ���;پ�nc�&Y�w��QBЋJ�����y�:��֩���O�=R��;�[���+������B�w��m�e"�4�!��70'�m\�Ӈ�i��5���X�N>=!N���/���E�6��w��f��ԭ�}ՋO	� �2��Ty�mA}iTm����OW=b,n��m����󆂕����~rٶ���Ó�H���2��s��A��K�MD�2U�,��񾢇��A)$�豹R,���&ǋ���J�=�����no!
�o0 VU����dKL_v��|Q3�����&~`�HfC����R-��#}�k���L�����7&[-q��+���0'Ѣ�{�������a/k,�2���̢rВ�j2v��2q�qKw�!�q1~�AU�v]���W84s�c��*�x�˂��d?
ZS$D^Z�8�`&�ۛ̩Ij7�����V�BN�|NzI�|�HH����M�A���~�X�tQ���t\{>��v�&U�Ҫ�w �9�G#/��!�O�ݛ��:���%�E���г禼���j��ûb���{��_�Z�i;�D��I�g��� ��<'�kޠ*�hJ1)"'��d3�=���8iU�Ϫ x|�'�JH<�Y[*����yԈ�27U��E��#̡2��'�Rk�䴰(�'�ыK�	�����wr�hzQ���
�G�������[�C�]���nM�	K��d����~4��g�P8��s.nI�i�(d^�ǘ�L��5c���(=��5�T!�L�f? rk;��'� ������iE�H�t�:�t�l�ڷ:L���Iw���< ���%:��jGy����7q�Gj+-\�2�?.#>�H�b�=��KzƗ�wB҉��j��cK�aΏe8�} �p�~ނ�H�D7�d� �S�M��D�k)Њ�v��b&���F~i-���Mv��Lzoer��Ʀ�Q8��`T<c��P0��k��2UJ@RR@�ݍ^CG8Ib)[�g3zu�u�H-���%�������[Ϯ9�Y&,QC�F�V�*,<A�s��M��0pj��/���7q��*�����Yqh�J~��LK�!i�J>i
���[B\o� ��K�q ,#�VC�R(�,�	�L��M�	�V�4��р�H�U5=H��֌�R4$T����Kl�T�����UJ������bȳ��Ӳ'k\t�{]�;���Z�K�n?�x��|��ߝxө,�� ���O���^IS+̐��Ƨ$j���ڭ�p�������'��� ���C���3NGҔ��bԲ�S�#H�?sIdB�6��~�a�o�%M�*�Ga�9����	��?�7�)��9q��7��<��4�5Nq٥q� ����.s���>��p��ԋ-�>�E�vi��r0��-��qb��x�-[x�:�wl�5�9�~��I��2�x(�v��L�tuL�?�}�L?C�pK<�ZW���^m�f261<j���FL}�� ���T�1��Mqt5vؽ���MI���ʲ��+�4������7�M���uAE���1Qr���"O��ژÞ6���X&J�^��l}��E�8VmN����CUXes��E?�ӈ�+�b"�+�a��|��5�?������/1��#����w鮆�y��?pz�]��Ⴕ$�L{V֔�g�	\�f����5��V�����8LMȿ]�7$7��?<����n�I)�=VM�$ur�ޭE�bZ�`����Y'�3Ev]��*ۀ�����K�$�wA�']��Nd�wח�~�UF�R ��u��1J	�?S�ɴ:�TTA���m�߰�e�?a�'g�[6k��&E���Z2>���iKW�7�Z�h/љ��M�5�3�>�ſ����6�u�äw�u��'Q� H��@W�u�h:~�O�0�"O%4��-��O���L�@��F1J��ت�w���/�03>�tq����f����/i�OwF�/��g��\�Y)`�K;��s:ȗ^���/)&*�\\D�A�X�!UAbg��������n
�7,=ҲPzG�l�1�&�,`ը�2@�D?ls�
�M��#=��X"��	j���^Y~$5@���]oH�1R�e�'��C9m�e;hE�M�ɷv[V�e�����d�����U]f��jV�Ӏ0�˝�ѹ牨u�Y�x�@�ꊁPm|�
scb5���0�!��?~�wVq�,��?�'�G=0[�órl��,��8Ѥ:���c�m�e�6�dW
�s4�61��)zʘ|�^���w�n���;��]�:��%���Â?1�������'�:��o��%��w�5<�K%>4.��֪��2X�0���f�ߦ�o�ƶ�QSa�ˣLՄh�iS5�A��5ݘ*�5"�2n���U<qd=usq+��#tImx� �".�����I�q׹������B�(������p�:�(��
��HM��؂ʒ��ec3z`N��-���ޑ*<��[��"Ǿ�\Ҫ�y�����줴����Z})��f7���I97/�ŋ�6�ze��`;�aP�<D`$\D&)_R���Кj5� ��j_!v2F�K�;qk�8���ݝ̸J�⹟.V�Ò��.�{����D�]]��F�u���a�d4i����!��/`*��J�uj13Ѡ��Gk���1c;R�RFge�����ןٕ�Z�� ��B��fԇ��Lki5�z�9���j�Y�|t�v;� ���6"+�s��u㐰���!����5>�!!�FL�fKNVy��=ȧS�l^��X0�+w��R��f��m]��k�'���K�*�2�$�&�z����F�0Cp'n���ǆ���wl\᳕3ݟY]�E]OL7���<W∦�4V2HN#��W�7����yS34���L����i;���`��h�(��]2jp�^���u>5���=��P0NWjW�ʗq?O{:O��?ң-��;��ؐOv�Zon�G 4@�шX�y�mB���g���o���QMG���"9G������x;�P�+p��hӔ�OR�:pL����ٯ�+��̉oi3��p& E�O`�/j&����r��Z:�f���~�L����q��YF�Em��<��q],��^2��Y�	7ׅ~lS^L���Ь��J�LY!g����5������~Ƞ��$~��r���� �bS>���T�k���y�,�|�@�n�Q����
uC�f,-KJ@��!Y�Aj�"�z��'KA=��f�ώ2����[':�$���kvg�g��`������{��L�ױ��XiT)��g	f�^h�e�	w��ouH�5V�x���!�4#�9���c��UPf�߮,��GK�Ӳ����;�V[����k	�R�} HՏm�&��gjzQG'��2]���0��6��#zWW��;Kb	�>L�����x�K����+M$�����/&���H:��=|�Ds�xU�$9����;��YkQ�W����Q����MED�n��_�M��(��K�M������GV�F�����	1Y�u酤+����RQl#�U�`��A�<��3u9�	���62��|�Tf��r�?�fԥ�+��
b���6���h�V�WʏA��T�u���Q�+F���F5�bq/�$l_C�0ۤ�/��l�GGa,A,ǳ�_Rd���vq�[4l�P^��g�e��J�5��(�$T�?���mNnT��;�(mGC�����t�=�r��Y�O��$�E���{�z�I�c�\~ ]B�Q� ��p ����){��苭\��I_vv��a���s1��.~�tK)3��5������1���Bsxحp�?q��H��R?��5\�PY�+�炐U�w���t�t�̈́8q+Ay2-���u�a��赌�,�J57r�!Xh�[d�F	��<�5k�5S��4%҃�u]7�yXɎ*��yD��>��Ď���!կ�㻦��þ0�Hǵ*N�{��«{Q�5;�+�A)��q��.������(�:�썑]�Q=Ȝq���6�8��3��و16w�ꨕ�kH�!v���
h}�rx,s�fb��cV_usp��Fo�a�D�M���N\H����J����f�E�ƨ�+H%Ta��1��sz�����s�"|��%1��\����ٸh���kp�Yh�p?�x���5��C.4���v�-I�8k�|�d��"`.�i�%��>���C�@�SMǅ���A����G���O�=�d�����n1١
+�T�
ʫ��E]�ΐ�(,Ԇ%�7��;J�'��!!�ŋF����s^d�e:Xs���}O�L���l�r�l��sxtl���ˤ�T��T�)4ÿN>W�(�s��く���(���r�����z�`ݟ��t��=����*a�:�S챼?��~��L���9�'}S��:@SK����ba����l���J�I��3[�-�R{�Jz	���$ ��6D��h9)���Ķ�U:Uk$�ފ�Ml�G��PgcR:�Z���B���tg �ej��|a/�%\�,A<r�0aJ�~y��V�fZ.�!��ؓ��
�0@��MFs7��&Fj�-x3p�`���Y�G������q{�4D��W��!����K����k����m��ڴ�7�0l��C8Ō�3��W[���4�5�.���裁�_� ��"����|�2�Jx^5LCu=$�0s�d?�R�mH�����,j�V�����f�ΕxO d����4��>������/BH]*���W�y֪	š���ۡOadYDD�P[F8��
Q�h�19_]>:���ozlC�����o�l��6�(�\綎��Pa{�M�BQ�ۿg�����xp��f�|O�x�L��<��?�{9֣]r����\Eɒ/��+�*vy�tQw���� �e-8�BM�Ų��K^���4i_���sx���*����>�����V�[�*�
��=s�c6z𣾉Df*�n.�[�~�rm"��WQz���mw7�P��E6����ut-P	Q��5 $�3��bag�06Ѹ�.|����<�����G��GZo��A$W��e�[9�[����5�kHk��}��R�Է��7�2[��X���"#�e�P�Bl,�}�5�4>��n���d��;��+>��3?R�:��}r����=0��(��e� ����u��s��_ɽRp"+#�ť����е*B�L�.��Z�M���-^�j��-�1>���v�B#3��u{_��q�~A�3�q�s�1�=���\�Sy��ɛJ�<�1�UX0���|>r����.g����,�$F�s���W��ʇD{a�,��W�X�?/K�;�����`"	
����M�,�0�"�N_�)K{TIA*u��m��'��f!���*���=Ч�$t6��:����jvf��;�	ķ�'߇t�s;��I�]$f�o8� B�(\�u�� &�����`��&QŸ0���i�)�teXF��B?�ِ�>Y˗þ)2���d�=�NZ8L	�+و�h����᫂I�9�n��J���Ǐ ��r�4W��z2X��W{�H'����tN��&��בֿ�)�g.�"��۟GhW�f�i
K4L���f\w~�"�P�K`4��:��=#^ⵤRW�-�Ó��3Y7���M�Q�;���=ߧ;��^N}.6�hq���SJK;v�I�2�G���J]Cʏ�՗�GJʃ�d�����d�2#zZ��9��ҙ���F����ǋ�D×����ӌh���2���t���ԝ�,���\,|e�jw����,��W/U�
��ض�:�"-=׹"ɴF/�
!�k�+�YϏh�l�1<8oT�M�*/�����'�]�����/� �3�LeEz�P6i��L�/�²#I]���eA�����b�7����ϊI���,�21+,g?<���Ո�6���A�[�:j ��x8����visXn��7'�RFj�E�*vcd:���J�_��7�H��k����0��׾�6_U����.�����{�gX�R���6��2ɆI�-�Tx��o��)m&S^GKF˒?���rK9�2��Hĳ�7/Y.z ���H!C6|�Q���D�z��Y?\5
G9+�x�T,�ggpVkx�b�Xc��rR�����Bʱ)�����0�b.Ɣ���%9�Et�6�.\�wZ��\*�ۺK�v,p��r,�"����
����v�Fop��P2�b�x6��N%��6�apL�N�7q��p�x^��q��t�>�$�S�|��x��6 �9�Gk՟$�`:���[A+Hݼ�}��њ������U�:�X��n��\wB"H4�D����]N��*ID����ˡ|;����_�IzT킃g-��/�����,~�"�S~���o��	z7?g&��c�����򺆾��"t�F�_��4L�k���FT�(#��J���[��C��y�M��{�9�c���y�uD�O��V�t~�k�Tc�u�a��Ŝ��ӈI��D�q��	��
��HJ�N�R
@��~���9k������XGfj&�����ch����&����a�ک3�r�IB"d�؅5���7�Գ�c E�`qV��q�M���*U+�V��½c^�@*����#��S�ނ}~X�� �kFſ"!�Q��v2��T8F�j�-��A^�r�ʿ)Ëx�é��� ����!11�i �4��6���kv�gN��m��Z��<˞j�X�y:@��@�R�O�F� �LV���YDs����>�z���E�6Ї�@�M5�����s�
��^�/��3�~:������Z������,a��̞���v�����r�pƌ�V*0�l<lǑ��|��L���`
}�wSd_��xi^	
�H@s
]�q�&뷱C�l: @KN�=��7�-1ܒ�z���G$c�VJ��h"�{o~����Z@|]�$��W3랤���胃�OZ����G� ��jb����Wr�s�-���q�I���~j�ޥOE�\501��ҁ�I9��h�a>�:@�%�gKt�^��H�zl��.6ҟA*��Q�H|�/_Rl̶&�:m.&�|^��[�v}��W���'./9�ke��@(&��l�m��iGZ���,�陸��Z�9Næ,fN\W��b���30C^� <�[��2n\�C�`l������F�i�1�=����.�U���E�f�Jоst���?(tǳ3��(~�"t���~�����I��������r9"� ��Ws�-���M��Ҏ�$�5zX��� 0w�ߧ(�1m�l��_���G7u,��@gƚ�VE�^|"tx:X��a�	�?�d-�iJ6��Ьk����f��ç>U75mU��L�W���z#B�	��Z&��v�6 <�A�g�#,�����:�ϻ�[�i�Ϯ;D� �c�|�/��ٞps3�]uٺt�"G��2W$�nB�.�Eg�����3��Ҝ$P��QeD����A�h�k������J�B#^��d�V�l�On�yQJ���P]�-�c�5I��Ƒt������ d����9((!���o�$S���`��W;��Vނ_��HT��<$�p�i�w(�!rG��29{O��^�M�r)��Bai�L�͑!b�Y����
����/���_;L/ˀbE�iLNR&vH��� <G�z´�Mw��O,��� ��yP�p)P?KIk�j�2{�H^��U=��Q57س_�M���;�Y"tg2)�V�����<l�,?����}曡��B��"Ys-���ZT=�'�~�e�.��^N�,a6�џ�[]�{>,�Cx���Jn|�ע��������so�9֮�ÿz��	�3��O���Fo�5�JV���B�������D��5��A��:��r�}���!�d���6[�r�WD>=|L��1�M?��$H����#�fwڶ*y�>�b�T�b`H1��u��TeE�&�`�2�b�Ys�XJJْ5G%򥚾@ tOy���P&.���-}t�"����&w*�۝��H�j���~�|��y��Hd�5��F�U�۠���}x�4��y��uV�qZ߉�7	V	Ƅ. ~�p]��t��%��\�m�~3�Q�y������[?uk�v8�R �=!>���ceN�k�Ht"/4�Ϙ�G(G��w6a�ǁ��YϪ���J�f2	���M){��!5��4<�uP@,'��m�Y6H\qnr6�����b���Ǟ�9]�e��H��K��a�n6ٍb�8�ݮI8Ҁ8��=LyNRNs���ղ��>�a�_
�b��C�5Y�t�����+�Yd�@Z���1�0fn��MnX�������)���n<

D�.�sF�c�d1냆'k �݇�G�ݧ����U��v"Қ�J1�_�ui0���
&�����W=����ȫ����!!��j,콓VIz%��.�b�Vm�a�_�O٣Ӗ���;RC{�*����gM�c����<��Tw�� �4�5$��h�/<�G��I�[aONِ3��1�91�4�)�k�����Kԟ2�~w*��R����)�5�H<�������y�{R�7���K/X��E����$pQ ;Y�B�zT{�~:�͏3��^}�g�s������K��;�C��s������o
�+��Y�m؟�]��"`�پK#���6���-ɖ�4��g�Pb~����/j|�Q�)�J�<l�V���f���"\X��h�P���?5�2Ё�cFb�c�b�����M���D���ԛ��.k�]ݍ4���Ձ?�d�0���ڰ�H�Y���������
H�M��v��H��@a��V�ȟ�K���y�� o��8���ѽ�s��S�eW�H>zГ!����t9�Ñ2)��;�6ZJ����U��9���	{=��#Z�J��aDY}��~�9*1|�O�T@�����
r�����G�߼%׎�_�,�2�U�K��a�?czSР/�D���\ڊ�vܱG��R�������
���e�DO���<�9�*b�����c3�z�,k�LUs����<d!8�N�#���_�n^�FunB/!��#3�� ��%���%�����r����  �w7�Dy����V�*�
0��땥��n�b�r�f!���s2!~i�>g.�U��ݖ�Ԟŵ�����97��L��#}�
�$��9IUa@cLH�ײ�ǝ��;(����Z� @f٨�ʧ%sv���v�T0�-s�R�M���g;)):��5R��4�^ �g'A��"`��ˡH1*c���t��Q���`�b�~8�L�(�[�<��4�E7Z��^�h��٩u B%~�jE�#�箜�6pW�MGU�)#��E?ˀFz�C'���Z`�� Ʀw�}�鯟!:&
�	�=1Aɺ������Q3�h���˼'�X-��������l{W�r��
6ձ����Ǉvl�O�Mr���S�ݢ���.E)+�? >U�v-9;M�oa��M�п�m�4z� ����_#�8a��n�&TD�񔃀��c�+�"�h��b$X��o<{Ĥ�G�h/�Wf)I4gXCc��ޚj������_c�X?H�mV#�/�"�Y���q��#�R�F:<J�	}�
5{cJ�£Í�������,h�����ܵ��Ʌ��̀�b;����`O%�:˪��1%�6���R�	�>��ĉi�����}�}����?�o�<r���.�p�ކ#�wx[	�.���>A�	���}���G����n��'f�B���������ԇSѼ�!�_��h-(�ٔ��cB��}&�h5�`��@�TL��J,�g�f���v��XQ�.^4��UP���|17a�9k�:zV<��Oe�4;�FR�M����T����ϒ*���L��}b�CC�2>���_���xZ����
�(�Dz���r�E�N���	�όO�x�u��_gc��}�0b�il�2�ZC?b��k��<Z�U��L�qCeT���p�DCF�Y=)�d�t���Me�z�_�м����_��M��?���D����9�����J��7���>����|���-Ko���j)�v���
��(��)�t);�B'#�M�BM�ÖCy��tUu?~�����!���¨���HCO��J�7FG���^B���|���2N�fP3��xm�@�x��i?CW�ͺ�kE�v�Ѓ���"n����ܦ1��2�{j)hB���)\Ɛq��3w�<����:��Wzfx�oh��� j������ٝ�\E�t(Ia�6�@�Sl\�E�v��_]�&gGIcY��H�9C�vRg���iu8'�(V\M�,Pʛ�i�O��a�8�5�Uz=0�Щ�ߝ��;CA�Jp���	p�~Os�1r��!�_��sM����+%Q5%�Z"��@L��4�h�W�����(��?
˺g�R�s�A_��4�S�B�*���!��|�i!Ŭ��k�N��T��*���߯�\	 \�}WT��T&S�YGrw��[tK�#
6ש�״��#g��N`��&�w�OMZc�.�����!���iׂ
��b�g�:[t�E���@�:A6Fھ,1�u������f��{�$�$�AO"���3��9IC!�9<�LՉ���;��"�r�R����� �>�NI�g=K�Ig�Ve�e���x��y�"r�}ٙ�.e����n��!07�G�
��i�V}"	���R?� ���l�d����!���&����ŵ�y�:��
+��+��?��Sk�c���lz��^hV�%���_�B{�ik�~U��x]E����� x@�d�b�՞k����s�%��t��?N�ݥk���CS����/꺟�F+�(�@�͐q��m/,;0��K؉��PKO�7wǾ�]k�B���x�����L�w�\\��+-���޻8B�%�>�����>J$�+�k�Kh'f���L!�?<��d�v�Y�$nʆ��$�3҃�C����s�K5��jTԲ0QdwHD�� ��.�op|�J�ߞd��)}#tl�ZW�^3�ӳ�b�����͡��`Q���W`���uP��]�Du3�	�Ț=�T�l���ÉQ���+O5�����;�V��s^��˶
ޗx%��5��"5�b��fI"���v(��q�֨�vץ����?ñT���J�����85[ma��A��.����2&�+����54�	W�r�/7��"�h�����V4E�)|��ݵK.wb��-���%�P�5�����m4kl'�� ��%'uޠ�D9T7f>�Q�5#�]��&`�5��8(�B�	�#�/�>��u��+(䪉O��K�� �����`�m��B���u��TOrs��~,HW̋����Y�%f'gL��q���/C;�ͨ_����pn!�a����IZrOu�!����0������X�gc~m����7V;����]<��+�O"�<�/��|e�x��N�+�Y{C�sw��CX~0nx�5Ǹ{�\H�Ed�B�j�g��v����l�K~��b�׷L��a�w�?j�1�H ]c��G�y��wW�Nӊ�.��e���.?��D��`�
�%i~x̷7T����>��_JM�#rK8���aP0=����0���%��q\�4*�(����[b˫6�̙sk�����U�CwhԑSr��;�����iP� ��WH�Jp��E�[��Q0)G%�5~AuDe�+���_�K��g�$�I�f%�Vt)�4SS]Gu躁��� ��?�Y�$�~@�ǈ7��٨�t���"�GP�
�YO.J��Taut׈#[�������p��e���]��G4	����*y0����N+�'m�u�|��I�~��Ns�  Z_���C��`��m�<����~�k��ZC�7���75�*�r�����`윣��ء}��eT��㬚G2�U���CnA�'k|L��]}��5GX"?߱��j���(+-B�R"���2�H#q���W�8�}o�}M=���Y
������q��D#��$ܵ(��-��B�$+C2n��OL���ͻ�[��=W��.9b��T��C��b�I�BQBj_��*Y#Vj�����2��1��H��<n���dA�8���q������8~J�ki6� ��/a��J�^� �}�}�'Z5�{IC7�z���?5H�j����d�v}�/')�4��y��"�[֮7�{h�Ĺ��k:����v��i�
���Ӛ1�쐔g������A*��Ϊ�ؚ+/�\��'4�W��7��X2�$���cC��5��G!U/�P9�����&��*��������k���g����>�$��DAp�/k�5@�jnJaŒUF|�hw{o*W!Dƍ�xT�]�.(�e�>�	���ɸ�އ0�8_+̶&�
h���a�*q_dMħ?����I�AـQVb����I,1��(��f�o��dB���?+
�Cq�:��.DC��}�͂�/>�7��D�yNM�}������"y���_�܂��p �D:���_,����s�f�d�@�Z����\Z��! ��ԫL�\���SC��`��E�[��T!������!���<�WϪuG=U��St�VU6�ov��r[+2/{�Ŏ�/�g�V�p��f�W`�m�6�:ݣw$V)�a�����7�ݲ7��R���,0.�	�p���ؠ�Ę�Q�u�Z��[q?�`���jgeQ<�rW���lF��-�^�Z�8Л��G2n����=�&����^�3��O�r��J�Q�Q�\	g�����Bå&z��KBU&ڮv���>����+�o�
��%�Qd�x'<kԟGE=�7#�0�~:��_cY��1	�,Ke�u+�x�	Q:����!k�lPx����%��y 
G���ۜ�Y.�;u:d`�G�y��=r��7�jz��f����+�S�q�|^&���VE��ݎok<�Kp��M�2�^`����8���E�j�{�٦�wO��B�D�M1�H��J�G�����XmI�=1�זwT�(i�/4�*d�#1����i`��t_��;^��h����}:�ԃ�Wc�!�"q�UYy�#+TM݄=��J�O�ܙ�K�f��׈�z3I�Uy".��	Y��z�X���H����Q��R�5�Tf}�3E�;���ϰ�iD\�s�N�3)}+�9�<��]�B���d2 ѺX���ͭ��j�>�hǎ�
.��1y�fb|�G;���[!��.o� ��(����.r�]�����r<��sw��)�	����PX��"4 6��.!_���L�3���U!7�����}<�^p��S���E��m��V�ځ����A�`�WW]��e=G� �Y ��o��9D�Aui��d6g��(4LCdg����QѼ���ֽ4$2�.#��;�:�Y���y<$0HW�T<�Pa0�2�)Mq�%<��ǣg����_-���AɅ�p9��]�n�Uq:H�˯0�g�E��c�%4o�_�6l���7pG���4@�} y�Z��g�� %�s9��Ǝ� ۚ5]���f��e'w�̖E&�x���7���.�먋E5��I�ݍ�����;�'������ħ�ş=
��
�J�u�*�3����vY��֙�zK�F���ê��gۙ��j������k��b��h��6 haz��'bBE��QG=h�?��FZ[¿O�4��M!��{���=�(J�'���z�0�����e,����x�z/݊,J��"w����w��TQ=B`FǄ�i�~[�0�Y��d��fsQ(���}�n!kL��8���Ka�xy�����I~��4�����}0K��$l.���">�̃���{�J��i�]�n�q�	`�=c�������v��2a�k��]K�7�Ў����Ց�e�{��s	�d~����	��F<��p��qZ�T0�	��i���2uf3<��W�S�%[iZ�D��Us�y����;j���âe�L̜��*F�?{�UW�(�,�*r:+����lA��*G�K�jK�5��:�̊�Q��o��{N(~X�l��_��SZv�����*FH��3�S+N0�/�?�rYj�3�I�����t��!D��e�N$VR���&b��M�P0���A &������������9.63�������cu^�of��������C��+s�r�a�"����b,����_oAL��:�m� �	z3�b��#V���N���]�������!�&��(���=Ǘ1E�H���9��!����W� �m������n��֚Tᾫ�z�c���z���H�^7��*(��Jé�9�(|c9����՛(��àC1���8W��4��\�y�nUcc>ۗ҄`5 ���:��i�f�Eh�.(�M���%Ro.�;��?N�~�Z��p�ς�~��Z��c�v���\i�����w{)$�D���r~&��aȞ%r�)�v�$�� ���I3>\{?�M^�)�4ѥk�S{��j��A��~ƥ��X�;�z?4t�����V]1EF�4{�Ḱ�롳/ھ�U�,4_k��ed
�Wl�$�a��sƃ�u�NvB� n��>\181z3&�۫7�ll5{y�8����{���+����U6�stc�D���S!���i~�)�QZ��23�
�w��P�nL��uVjT�¸���n)�����Y��[A�rCs��{(�����|2
��yI��%���b�5��~uhFh�M������Xr��B^��u 	��-F��p�;���4����}���ò���z>�R8tԢ>��s,1l���NIn��'`a{������\��`����t���F/�rt�����WxP��Oc���<V��D��� R�z��w=+��ؠ�ĆC ��+�U��c(����hՙ-bWp��;��C����a��kwiF�S��L�Å±�,���`|�%��[��(�(��J���{��@�W6�c,4�~��������m���/X���9itj���i�UQ���h�p�0v���f�"N�K�di�a�)T�J��Y���MZ���iތY�����#�|���,~)MAY�s3�� 7X�O�41�բWD�5|Ƹ	x�0���ݷ�a�j�c�?��MZ�
���2�������d�4K̆r�b4�X��`b�-���ii�ms��������� � >�ԍ	D%F{E���)6T|��sZ�i�3#�U�[����u�<����r}�	����\�yz���
���c2c���k����~0�k����?	g�����<L�u�;KϺPր�;n/��e��N7)��_�F]Ӂ.�]�OH-?�j��s�I�
��-��]�F�p;Ъ�HP�}�ZC��dW�\z��;�4��c81{ա�=�a-�����	����ao��錂	ZM�#3�G�S&�2�\&���v�h���A����B��I�'ګ�D����փ��d����"s��1����0��r?�����ěh���Ӊ��l�n��e�N��RPVbgc�nA1q3��k��SJ�k�\ C䆡9�N���XW���NFy�~
}�u)X�yP����1��Ζ<��@��#�R�p)b��m)����=7���E7�-��[��������u,���%����S���i2]{��{y)}�R{�f�m��B3�:��(�l��_3Јe�*t�6�jc#���2�S	�z���?�v�b�.N�L��?#J�G~��5�w�)DV��6f��|?	W�1��1M~�v���v��"`�}�
$�۱1B���O��ωZ����فFv��$�S�L�9�_0b^A��d��}�/�
8��z8�82��R*�<��K2�O�~Rs�U�Ƌ��V�91�����J�I%I��5��w�Av^K���f>�Y�R�����g����z�97K0�y��=�Ml���D�|uC�2�%�h��G�Z�>��U�e��0xZ�E>O(|=�;�5���v����@��Yገ�_�J��G�}�(�k�Q �I�a*.@kĨ4��qW�3å�yٕM��I�$X�g����mN%E�D��Z�	Z��^dS:ט;vk���Ǫ�[> cͣeZ�Q�u�������̓d�
ݼuK�)�~�mtpe6 O��*�H�P]�� d��t4v歂�?�D��;�e����
�������΂fu�n,�|b02m/Î�5�¾�?������H�J�`������#F�%+k�΃+�0�����VHq��q������7Yy�4�l��~B�#؞[űt7:�n�h���Í%1I>��3�󏒩�
j2�e���_�@��?��Z'�)*��s;������ӆ���բ{q{�DJ5�|�bb�<r���E�X;�M�P�
��������H�v:������Mxϓ�\"ۣ"�.-�j�lv�+@�4W8�9b� <$�jzR�!��B/f�E��Gf*��f�~��5�y�$-���X�~mg����
H�2'�j+���`FT����V26�^��$�
�5WW��N=�~m!\�� ��׬��>6�����6��5�eŠKx�4X
YjrA鎪�{��o�:�����8��I������ݏ���|^�� ��pܽ�R[Ԁ0����O�C�hD��C��$oH;��"j�5Fk2YA:nO�W�ip��h+��Q�(��pNR7���%W|h���R��X1
^�7İG������C'/J���\BU[�_��2E�nyx�V�v�T*Gі�c#g%Ǿ`��ĞZy�ޗ˱}�c�F=x��i�߆TL�)(#���ʻ=�� J^�)�(	�+[�0��Л`��7�O�9��b�z�\�J���`���F�T�c���^A�O�_�P�(�~��u�]&ɕ9��(R����(W�.���'��"�����7����oG��-�yU����|�O~������حJ�>�9o�����$���b��m;*��W��*&Kf��4����1��.0E)�P5���h���z���F��>-�!0c[�L╧
��K��������i�	���o��y[���iVoR�^s]ЙP�ZK��j���k��c�O)��)	����+�U�F��W�y�"pí�#m���0��{����nC�a�A���s3�0��T�ExC��t�����i�B���]>*��&f�V�p
��H6,4�F�f���Ţ��W�5}h$Z��Nf����.��]a��xd���b�"��>~6(Ӓ;�ee>dSO�i���.��=�@��]6�b�����S�$�B)S�Х�ݨ��8�k6>���K��bB�Y�r��p}����N��d.�՚��)P~'��'H?2ŀ��fk��y�� �i�#nK�+Ph���җP!�/`FO/�pc��0������TPP��Y����o�_-�Jz����옪c��X�knV��T�︃��DoK��U*�E�m�N��RՂ��9�� ΃�p��4��v15MgNc�����;��G:�B���:�!C�=��#,#�[\5aY�Ey��=��p8a��ǃ*�\�q��4U��(Z�l,b�T��7٥p
�,.���c�=z�r���ٓ�<��?lRa�Av�>A�6ҟ�n�i�yD};��]�4�����h����t�q�^�U����Vf��!4��"s��h&̇`�E��\U-�ě�k����)]�2TPq�p�H����Ǫ0mT�º'u�44�=�Of3�/ �z�y���S0��{W�_���I�c՝G<�]�Q�����E��&�׵;��zV8#t�-?�5��h-6�&��o Q ��rȈٌOt�ϲ���hR1/�P�Ua�9�Q��|��2(uT�W�$֗U#�&9��`�yoQ0�|pɋ(^�a��z
�:�1�A[�.
<��V�Ȃ���&��)R!�c���1��, ?;�ߴ�SF��}���<��X����CÝY��rq3F�G:d,��m�L1�mD�!�i�!9�e�xLӭ�y���>U�:Re��S�Ȯ�
L�҉א1�5�x��k��Ϥ�^�o�(�����EDu8\�!�&��S��k���N�.����B���kx7lh�`��W@��=�:���כEӜ�<GB5T��?X(ZD�Zػ�U���_W�� �m���lf~}�d����Ʉ�5+kIϞ`���/m2E��W�J�CչG���mݽPZ��}���ea��u�~�F��%�e�|Oм�����n�f���x�ry�����˄�o���1����P})�%v��f�5�\��Rqs'e5�Gp��'���.��$����ϣP���]�;�#a
g�s�7�Q��+tI�Y���KU��K�$�����(AX�Ey�������:��q�	]�����h��Sǅ�ϩ{��gZ����:���G����;���*������l���b;�6|C4��pa�1����������:���'��魳�6�i�y7{OA�g��D�3��jF��&�=l��u&I���"A�m�]���Xg7���9���2��DZ��jW�3U֐�}���-���T��tÛ:,}�i$N��272��_7.���'.tm�CX�Ï<���>h����\��4�ZjTxp�彌��6	�d����(P��c%�Ã����z����k`RîqP^$NGˀO{7R���b^xv�dJө#��_$�6txRZ����#4_@-P�,L0sh��$���ܪ��كI�z�(1�������&e�W[��Q��US)���ZX�=�Q�(�����}�_K�BRk��B�g�G��}B�Nc�r�#��h���w���-��`r�<�u�Qg4�W��e߅9���f�	�èY��u�<�;�<���; �ѳM��tn㈤X�/^`�c� 2MI��E�h9<����OG]����Ӽ}��q,ײy1BT$�j��1����]=Yc�5.ӏ���g��"pS�;h���T���L��!8.�&�h�Z�i`p�|Ԣ�cy@c���x���ǭ�#dg��n�I���"�Q��F8v��GHk�@F	G����i�Ż���Dd�Ǒ�����I�b�g�aZ��)�=��|q����F�@�wJ6Vڧ�:-��k Bp4ǕKXf
���!�u؋w�� ߒ-G<.6���( ���j�gJ��ڷIn��e�L]�x_Xy�';ъOd�=����#Ã�qU0���A�$+�ɬ*��
��=(�kԚI�����.����o�K@�v�r�w�b��zGA��9ܮЖ�S�����v�Z��?���yla�<�o(�cXx��6N��țV��%/�QB�'f"�ȧ}�,/$	s���
~�)� �LNv�������y�4�+R�ۮ�b��>̈���`ڦ^�&D5fbG�g'�ڡ��zj$��`��)�aY���EQQLo�l hL�@��k�}j_�#oy��O�v��e#���ŧ�H$��hK�A��e���ㅛ.R'uc�k���ngK$u�O��E ;�X'm��͗����N��yb��G˩�WZ���B�l~��6������`
�p�2���aӻ!����)D��E�3*-.�k��'��Ƿ�y!G��y	o:{֐W�L)�^���x乮J���(�Z�t��u�<bض��ʫ�p>q �PC7c2��8�ĭ8`��l�η��$�+d����z)Y۬`u���x�شj,��#�2#A��r]���ڒm�Bz���)� 4�	���~t�tlz+=����~/��˚e��լ6������4AT�6���@O�����t_߸,j�d뗪�1p��Ա����wL�ԣ�A�빁�y��z>R�΋9Իr��xx��[�{�q��d�DuЉ�oo/[��k�c��|�!�@�4�9�9��)V��mP�l�(Z	�	AV���:y��:1�tR��-M�k]V��d>fV��;I��\_lm�GG/k�����)]c���AΤ���kQ ijw�Yx��7��np S����T�b��.�F�͈TN��$� ��X���}���8��Ao��.�S����
��LCnR���/���+� Z�v��4�Rˏ������AN�>g1�X�P>�)�H5s?xۤ�����Ժ���oӑ��N�)�����29�S7��.&�R�Z����1�ڟ�0���:9p��[�d�F'�T�IL2�G���])C�}�u�u�����PY�h�w��.�
C�q��C���;eL4���K�ˡ���{2DA7yHM���Q}%oM�o]�0xP��O:Z�w�Hj�p^�:�4��M�{��o���`Ġբ����F@�vn���wJd����-�]L�������a�,�#��:�?�o8��*[Yh,u�]�N��!Eg��ɩ$�v�Ϗ���,[�ܝ[beZ��Z���)ϭ`��I��|��?�]O�jy4��)	S���{������ �	�4���N�@�~���1{���k�8Gz"I���db�h��/�������{��x���z ,��(��\��%�@ʦ��݀�dҠ�4K�?���_�Tr+}j ��F�E8��"G�����G� �V�Y6z�A��.�V��
B}�rg�j]Z�B�Սr��~=�%�l,m��B�v��L|���&��9��aSL��ސ\w II�kN��4� [+s��ٙw8�ؑP�#�Z7:WNv�S ��p�,*/1���e�m���(�S�]mp|�-�*Ӛ��s���C#vG����}&1G��t9�}�Q�^z9�F�3�7M渞�G,X�XO+��U6Dtk�{�c%�۴� ��
��)��IѲL2�����񽫹d�S�O癭���"�g�^g�`�q�fFD�i��;�& �����Gtl<y��d��W���J���ucu��D�~WF�R!��H^Qj� ��9`s� a��c=*:��y}z�&P!���4�����"�ZCS�pNe¸�A��ދ�v6��M[i�IZ�MY�T�&i{7�~�}�b)��{��I��}E��f%��̏)g%s�Z�pL��u�0�T�UF����i���O�d��J	���`Z��4n�?�]�{H�o��| �4��ᛞ��푤�+������~.I*����ֺx�〄���c��~W�X��AOP@)���*�j�S�����_��(��	BC�" �:/�b��"�<F��"�ᏂU.�Ȧ��(�`�U��J'�ߟ���\��L���^�2����r���qiruF-�����,?[m;�g%D��!�j�W�#fK�o)���s0����'i]sИ��sc�v�A�g�`=.r�ʋ�*��l�c<J��Ɇ�����ݱ)I�@�1M�F>���9&ZLӒq����h��h\���#��N
��/��0�L��]���.��ۗ�l	��|-P(��d�t��@��É�S�?�� ����Fe���6��<e�+�9P~85�ÏPGA�ת�J��jԫ�{����W��wԜ��"_�w1��S�rs����P@��-7���Jؔ0��mI����E@�.�>�n~C��D��A>�9�a�w�hǕ��_@к�J]dd{�N&�w=��$�>xn��(:��M#1��� �`EG:�'~/��ꇺ�O�|���G��Y�
صE���ھ�m�@hy1�h�9�u�m-\ 5+$�4aPՄ��\*e��ƤoN#���ߌw���\N�A��1�2����CwM��FOȳթS�`��k���T�d,�����H!~o�r��{@Ɍ��@�����$<��b!.��@���g��'���S������W���aX�c�K�p��w�����ʿ>�M$�av�wN���c:Uǂ����θ\���u!�a�GS�s�AZ��1&����x��xN1D��A�x��en����
�ٲ	D[9����혹'�o��`�����O8�7^�������ϛ���
"�	-U�L��RE�[���Xێ���m�`�`K�wgō���)_�7�%�I71��j�z��y�gagn�TUw���W��MY�rK�I�\�+a��^)�M�|��+0G��<#���0:���=�O�M�㏝z��g~�;-a�:��}�wW E�'h�HB��+J�q�qr��Z �<!��h0.s�\�2X�D�ƅv,��}�$��\B�ß�������W��1����?n� �5���g@C3��V���`�g����U)����I�'�EY�����F��sI�~䀨}��Lbu�w�	7�f�m��a����5���3�O{s C� �}�&m�a~fq�#x��'�Lw��s04�p���Ya�ܜ��]�>r�[��!ߺYu 3����ʹ	'�d�L�ȳn��w�PEK�\l�ޱMa��U��Lp��G�J�@��.ţz���˥�	E���_�-5=����b�<M���1+f�an�__Hn�*��(��$_���aA&r�%�/�W��T���s�Jn��t�|n�(?�;�/��6���h�C�	"]��PQ�3l�K��4Qx�.���"��;`����S���$�XDm}]� ��#���	�������`��2˟������m�*��J�"W������;\cNM��)�D>���L�g�*���h���%�<��BY`�3�� ��:��`�kX���a��F��6�Y�{���ZeH�!���T���etË�^L�Tsð�hrmjgτ����g���vuF����[����\_Y�~ۤ��0����Ug����u�����t��6`=Dو�Z�8�ԿM{�0U����i�m����BlaZ���x�j���چWˍY)i�چ��O¼7��^����Ͼ����TLbQ�����_D�tN������?�ٚDI��Kɲ�����^���]�J9%�!��GC�`��}\�Q�ٳ� �,��n���y9(���PΜ�����R!��h����5��?WV'�i�}X.O�J^��N�I�e�4�1��x�T"����,����H�͑�C\k�y"�z�ţ�]��:C=�>���F���Imb���X470�����R�e�4\�	@�Io3�7�v��E�4�Ι{e��]�9&�����SU�wO��ߊ�)YH>�|j.!�9t��k>�6�[�8q���Q�6�n��n*�*������6��iG����=Q~e��fz	AK�l�'`al��bw�l����2��\e��H9�^�dHyrH���g��C2]����a)��N��P*"�hQuCP��+C�Yv��\����2�f�Pv���\�{U2`��)�w�e3Y�|tE��5yߝ�w�{��V���p�*��HA��$�[��Tq�
Cg�F�\B�S�͝����S��g`�l +�Y��y��N��W�0vV0��U\�r�~�T_�@��2�9�;�����V����Q׶�y��e��$K¬L�����j�f�qH%*��?�O�̳�p���&�ZwM&n�f�R?�Z<��h�a{�Y^�4�a���4k�YR.!C����+	_�˧�)��'[?��h��� y~�[lN#��e�'���V0�/����}���T���4��+@�,�l���k�Q��[�*�[c|ˮx�;���W�W*��x�j���H�N�`�����k��KK:b�6#�T�Je��L��ψ���`�>uv	�?Ҫ.p�m�b�ӄ�Űh���[�m�����II�}-x�4��U�`�<�!�Z���we�����!��*]T7J]�]�!��͕?��3�o���n��8O�U F�L�V8�����`o���^p��o��Ix, X�.�4��Fϣ1�ߢPѐ��is��#b>�T����"�X�`7�i[���~Q����,�z��
%��x���H��u� "����'n�cW'����t�l� �g��k�Տ�ls�z4(M\�T����o� �ה-n���9�4Y.@K ve� :Bj~nf�⋟PJ��~�3.� <�8i%���B��3���@��J���鬬o$�g�1ÚI����,^;��%-��\&#)�vκ�.����<'C��������e��D`�mW���,�$X���,ùwJ��BG3#�K��=风XH,�����W륚� ̳��p��u���g�^����-��C��z鑦�[�I��4�3ܴ�2T�k:�ל#�( (��F�����v"�;��3E#-ۜYߟ�j��E�1�Sy��U��{�w`��G����o�{K�U��0,+u�� ɯ}]�c��.�B��TYu-�d^ӻ���K���b4��+�GtM>�)�
ؘ�X�p���Ȗ��M�_Y�����!Y8fX���G�؉����vI^W"���(z'O�8�%*'�i.�n��9�Kk�ӂI����f�Ow#�Jެx-kq�@����=��'�!\����9Q���
M,��/4N�ϱ�9ߐN�ɭ��MA ��	���(ס/�R,!*;��"g޾�fZ�:;kɗ��Ҋ~υ����La�3����J<�1x�oBwc�^y<��Kn��~S�_6,q��S����TC��p��^�c�5�Z*fx��⩗]�
��c>���s_�=���;Vڲv�9T#�J�~�5(x�����܈g�-�
�ެ�Xe��2��5ebd�R�A�hᔥWHH���W�K��
�ep�Sۘs<��6�Ѐ=
��4�=�S�����l��DS�x��h
G��{qYl��]c�?����XQ��T��K�<�V���k��Մ^����Ң6�T���P?Eԉt#J����;;0�C��X��$�U��;!�~=��� 7��$��&~����|��&ɞ�������Odq��/F>P�s	P��Q���=��VEn�*̆/�A;�����^­Vu��4��q��ԣ+��ό��߻z�{y�"�*�_o2MQMp'"FǙ���O^����]��MQ��P����Q�:��>0|�'���#H�n�r-�L�H��f/��	���8�j��T�<fET�j�"k��J��}Ƌ��e�;�ڷ�O�F�=�Ы�Ct;�w"7�F�أ�
O��n�
|Aـ�K�*�l�� h��U��ݸc���$i�,��J���Z���u�3?�2�rt�dm��n"ո�l`z'(��h��H|���h��1󻙦��ʲ�ؐ j�_H�Nд�*ڪ|M�!�c���@n���^�B�M�+��\LF��gͶk�r{ӯ�`�x�W!E�W�i�
�t��T M�7�>���hհ�꓌%jN�e3`IC��uՇ!?�H�H�y�Pd-./q�e�B�^��?Q;螅��s�	�=E�H�3�Q��L��Ru$p��Z@��<���:+@yV6����	C7+'��t8v�l�D&��b@<�� ����r�"Ӎ8�����[fSCa
ѣr����M�d������o3���̘!�YK_������ƣ��+0�J��ȔR+��!.�t�lq4_{�[�K<�h5&�՛H`�_-7��;I�5����^����2E�6�1�T�fgҟ��݉
��lխ*�N.$��Խ��&�*v�OR� [�I���c �8�W�h����k�v܇�uy����
��G�! +6Ռa=�l�-��}�̅C9Ս�� ��D��XX�����}�0��Χ�!��a{h2BA�j8�aOu6yc7�ːBV��_�TR�3���+��88{�G�S��3Y����>S 򅦊��4W�(�'��Ay%0��7/���lq�5'� �1�4�+B��'��YXddK��A���FZ�,R�v{���ɉ�������a
�x�cu���s�I��8�v<�>fU e_w���w����4:m �D�/J(0��G~�"�E�ɋ��N�Ō�-��x�M�$BԼ��t��$5I�{^����6�*t�V��7�H9�6�x�xe�2x����S��DTzc�����̛��p�e���K�D��G�s��:�7�ҍ��j}�1H�鲑�x�]��#]�;�2*�rB_o��o�O���w}�LI���d�KI�I�𺊤���z!l���ʁ�8��.M�m�{pd���;�ѷ�,�Wp�xn�2:��Z�vП�D/ӌ��gnJ��n2Mvjֵ�"���R ����wP�Ϝ���d�L@���g�Ǐ����2���^D(�޿�#,a5^�q�5ڵ����v�c�):)��5�C�)桓;=b��sa�.����~O�^���H���1��g��l:�����h��iFza![ȳ�M���ߞ�d7���Kc��O�"2������� �QGE�?���4}~�`p>�AL�7��D$B5����0�9O���pYb8X���������`��2���.�Խ�R�N�}2�0ٱ�C�D�v)�7)����~^.�k�p[�?����7Ep�W�*uN��>[m�<i(�<DR";����ZNzҪ������d�����6�g��B����f��2��^�D��o3��g��]���Y�q2�qx�L�i����G������
����P������bU
��n�l7�5��P�྾r�w)�����������9{�����,�B�f��$o
?�CNۻ5R�Vz����>(/ #y�qX�C�͚p��r<BEn�/V�1 �}�|��O��/O��A�PփBʨ�u{��=���u���Ύ�؈T7O�45�\d��)/�O�V��C�����&"��I�RX熷 �A_�<��"^b��~�Q@pD=9����*e�� �����o�(����b�'_L��m�Q��N����^H���g�΄F�f���5`�h�Z�<ܞv[�P�SA@}3ڱٱ^�\��X.�oo���Gd���
�Q���~��n�aZ�d��ǽ3M��5�]q՘Jz��qK���0��_l%���އ�D�sjC���R@��;���HH�,�}�uF��I�7�gzXL7OM�9@�/����*��#=6�zXl�"��S��� PjG���b�^����;ݱ����b�ަPY���u�l��o90F��c-2�*�
h&,���IY�E��V2��P��<V��o�[�+�Gl���J#�%�T�o�L�!h*�ϥ�����=�wC��(!�4'���/l��A)(�pS��*!IoHdm�µ�`=4�L\9��"BLPG�r|��g�A@�a�a+�O���������&C��/�kȎ%�]�eUj�*o�7���D^�I��9���,*�1����@�	���9'�7�?~/�a�@Um������@�q�d�;�=I��G��N՟V��i���%8�GGd�,���7^�-�6�_���$�=�۾�V&?��u����T1�<��B^��D��X)1%� zn7��'�y�ڼ/�',1M��c��� R���M�	�m4�g�[sZ#�Ux[���Ԧ7OtK����w�X'Fm��u�}��[�w���?�̅���j��%܌*5�6���D?sLf'�#ʰ��j��!P�|�u��M5G�/��#Y?4i}0���:E���m[W��W�0�P#��xaܮ��mP�^m7v���8�'={O��HHkΗ�I��A��4�z��^�l�o��Nw�]ކ���|.����&A�݇C9�̏{!Le�kށ�;'���/�]F�������)�7�N+{��
�^��C�y$�[�Dn0�
�I�"�xC��N�!���)�}������(��.+����7�{9r�E&.���؎��$��$�JS�����k8�@���`#�\#�L�k��|,y?Y���ĥ~��37U�\������d:��o��F��fF'�i���I��U�r����V'�aw�_q�pث{��3z�1'�b6 EB��pB�yT�d����^��.��( ���D��WM���E�D�����Ov����))L�6!�[ǭH��&��u(�G|T{T���4�
���%��`���z6:��D9��8��8�jK�Vpo�L%,\�_r��!����0聨���i9����=A�c~����3��:@�g�r<��`)�k�ꬂ���et�L�L/A6��ԧ�������D�4�-��ZC��Y2�a�>�,��u3FX��O��5�-P3���_��@H��e��Ȧ�x�w)^��F��"\[�6�ŏk��,�O���jGo�NH;���]���|�1U�6�^f?�����#���D	P-Ňki�Jʚ�v��Ȑ�m�O�WM�$��x�,���/�eԨ.�t5�{bGs˧�eT5;Q�%35�{�KF!�`��Z�����7{��$,N��9������<�m����Յ倁^o��1?�r��<�HaFB���=��Ie?��"�(6�K[�^�G�BGo���.xb	�7����]b��o����{D��M��.�c���ìz����Ѽi�s�'�G�����Q�"�U�Yc���+�;��2X��Y�f�e�������O�mv�tT�-8 >�j։��X,`=��S?4�����!/�`�n�y��>CE�����Va��K�����hy'i�� �hnq7�(�Mn*��mKf��_6f@�H�7��	2h���]Lz��gb��Q�7
q(l(�]���۔���B6���x6;R�T#��@��9��'�}��j!���wnɪ���=���@J�w�v���X�W�x���zW)j�#��n��H��_�2��>C�E<����-��ٚ��^Τ�� �z�7��R��1�2o���͐�pAw�'��J�A8h���6�՟s^J��a�ːĕ�,��}7	���e��U����(�����<Y�.�s֐۴��Q�����n<��+������Xԓ6+����\�8��X5O��=d�`��<�Խ�ǚ�21o��ڤn�g���IXc��0g6B���W,��lc�=��$m"?������kq�u9�飼'��my�j�Y����( Ui��%7׺�y���+e�	wK�����f.�(����ﲈ��O{�ǳ�㈒E���&;�� uz��*���M�m��2=��x�y8�s�����0%r]0�ǅ�ى6(��zh|�<���SPX���x!#�m�]WG:[�y,~H��I�xNC���K���k� �T|($�BɌ�KV���=���e���� �8r���|�4�9�ﹰ�>�tS��zt�f�R08F�����ah�:��n8Ί:os��`��h�w��	�zzWlIP#����^��V����` �0i���Q�=^��j56뾦[,��W��ؤ3n�[[�FO�,���N�D�O����l��GD.ܟ;Ϫ��iL��wV���Di�u�(����H�w��<�(C��_�MNSQ�^{���I�=4�V��Gt���uI�4��L��T���oȯ�>��A��#=� Ъe�����m��i@QV��q+����!�>�f+ �X�_"��m��"�B�\��?�w��/�,e6�n ��꾘4���m��ǅظ~Uy=3��,~�/��#���}*�PQ.�0F���q �o��?�밢#��X�3P�YƷ����f���i�=7�=ZT��gI ,�%��Ms�2Z�9�R�	�;*;���p�W��c�`�O/5��3�a:���A6>��&λ�� iE�ҿ�����7�jh�(T~��b��[$5!�"�;�׾���q���/�P�`��W������/v�~v?�d��6m΄�C���.Q]ay��Hf�;��E2��;Hp��ԏ7�%�2+hV/�pί��qV�p��a��_}NԞ��r�i�9r�i���UW����'+�t)�_h*�$����
�d����&߿����}E�Y5��_�ը�ή!���]D�7JC�O�5��r������s��:ol~�q�D�ȭ��4l)�GKx�v9�@���y}1�ع�b[��V�w����^�1���Du�q?����4X��3�����2���Q�by �@Iǉā�3�%�)�(6�ܽ���j�����_R"}����-�|�hD�B�johK�f/�[?�9sګ`)��VP�H1����Mf𤴾ɖ��Z�4�~�&<���%$�M�p��B�x�#.�<v�d��sD���Y�݁�o��0��ߙ���"�%zER\�T���x4Cǟ�@�f=LFJ�?�������]l���G ���!QUHhd_���������LO��#�}�s����O�͏V�)Ӡ)�*[ \�΀������g�W�cM�]2��t1���$��2X��C��p�W�����tl��E��Ly*`V�CO�n%2�񥈇5�0yYl�%V�2i�:P'F;�X�R�r2�B�y�,`s�������;�y<��J����&����|~: ��ꢓ����:[Q~�<���W
2�I����/��2�P^;�h��#Ov��}}�`��Ӛ��H�_�%�c{��=���Vɪ\^�<�䮣�l���de�5�O���&g�Q��wE�T�e��'!��B�ۮ:�GpT5�����]d�G��d~��sl�ˊ��� ���H�R�j�>9("�Un%��I �����$�{y���{�Nެ�Ԏ�1s2P��6��7�i-���}�sЪ�}��D��&��is-�F�� 9�jr���~�N!��|��8������9�y�H��`C��Y�
|��9�o�Wj�vK�?E��
������4dW�_����]��a������k>���!�<�r����/K�X���%i��YF�΃d ��u�6UR1U=��U��8��Y�j�;j��ۤ�B�C��1�fv���rU>�_����=N���T=���iͻ"��hdwCCgQ��:���Zq��D�KL-Q��p<~�>��ތ���_}48߸�4�2JJb��� �gy�qAH]?���c�ެ�xvd�#sW�ތq�H��:�`���x��kO�n��;	�¤�KG v��S�[U�$,#W��Ƃ]����2ϻ]c>w��{�?�SZAޚV�Ӫjr�~�$��p�ܲ4�� x��$��в@��Z�e����M�K�u"���{�bG)�ŕi��瓯�4�W{�x3��3Eu��Ĺ�$��p/���ڹ �}$G���qq0GC�H�0>HRV�����=��msI�}��	2�����@��/^)r�.�'*з�*��F�?�
�0��X���=��������v1��Y��%+�z+�]p=^drSB��vUT:��&��`����@��!��4
ֳ�W����<"��nvEdbU���9��B|�C+�ֈ����A6�̆����)�D~4uﳀ=IM��D���\ٿ����5�h�(T��5{��t�K���X��T.�5���B<ܿ��-cQU��'X�s J�y��8� d���_T雓�rK�c<�)6���Ff!�W�q�?�jhඕ0_�f :��p?���	�Pb��V3y<Qm��}�K�dK� �0��ƀvwp�D�FaS��+<�lR ���X�)��/�J��;��G�R�R/3�y"�����_�)��*�=�����^���ȑQ�Y>-��ۥU������Q�I?�A�MwVB���
�h^0���p�>�ir-+u��E�.9� *��L�iw�K?\@
�W�����}O�Yt-cfsS���7�3t���� �k���t�T��)(�41��,���$��G�pByA�p���7yC�J�=49F�7uzYF�`-z	�o�:ܯ��2�������@��Η�������J�Qh��+�Ʈ�)������2��%V���� )�0�HX�ʜL&�^�6�д���C�u������fr�Q	�YK�k6�`w'���f!K�dEdsu����P@Y�!7�@�t�]�"З�����q�a8�)w�zˍ�ZEp����6��z}�Z-����3~��3Z�И�Ykf�x*����o�����	���I�V[��|�a$�|�=S�x�VG"Aؑ�ы:&��X��	��.Z�,����tb��_����\Cq֯���B�o��Ʒ	�M`Ξ��+�G�)y�r��B��0 �  ���4�Ұi E�m�S���, '�dz�6�[9⅒yW%�$/���!���� ���
�b���2��:�̚k����	#)�
�X1sv�!T�xPzg���1oM3�B�Z��
4V�\fP~u��P$�n"}?�I�K������o�nŃ����1ad���; ����;�izR�8��q`�E/�\R��ۖ�&�Z:#�'A���	#��Xq_�"t�%���zgo�8����+�Y���;���P���}>+z���6��c��k��>�n�$�1U#{�%��<�b�(<���/�d�Q=�/v%d֢w�0��S[/�o(���DB��q:I��R��l�'�eb�΁u���i�7<�r�Bv>���*<�o�p6��m�r%���0���k �ؐ`o,���Nz)����8�CC���A�v�pSV���mmJ�<Q��M ���j��C�1M'�R 1�C�������ʢ��vL���(��g��/�<���z^�>��*��en��S����:�V>Ht�c�����b���!�Q^4~�G��@.A(�z��.3'%�D���M�w��K����$/�/�ha�U��I(D��{��|�2�btF�>�/�<ȏ��F��D�n6���t��Aq��r3G�������E���fkܚY �'G!�v� �7,��D���f��%�*��C���n���.���G���6Jo�-�c54�h�S�/��*���!IUU��Co��v� �~U��*�.{�]�EQ(B<��3��3�������~�a�G7;�����ϐ�
����W�$��c�Sn  o���ζ�S��V��Aֵ Z:�`]A�=`	)֙��@���F�;��؆m�݇-�lyt�-i������BG�l���T�� 
�,�%��Y�l�ZG�}��ۋxLjv%=���rNM��6�[2�Ao�;S���Gz��W#ԛ�G�5�ڛGJJ�B�n�X���oY�$C�hq�4	���3x$�x\��:�<���ҁ�TF�;!hZ�?���"���3�:��|�K�?��2)NŸy��zX�����T?hVB&m}��J�s)��0t ^n��)�B�����B�S�·�Gt�În���"�C����6��L5���� :N�(Y `���<�b~�r��vnl�"��`���٤fM=�ӵ{�I$�;k�uS	���QD(��a�g�6��'�_��f'�jW�*�H%�m~����k����#@6�O<�#�eK��u� Vsb�?�C�D�4c��X"�2��N=(�#-�|���3\,-m=�^���rA'��0���k������G�K\�J�t�i��s�J.����
���.q=\��OkQ��E��Jʬ��y�j�jf
����N_b�����F9�*eؗ<�W�c�|���T�[���'_[�u��c�i�[g�璕1��	��H��$$��͎jѮ�>��/�5T�v&Z�����QVY�7��S=�C��MyҜ�%��"*�mz��أD�ÕI���T���n�,���6!�G:P$y
�rB4�[ ���-�6�������=�UNr榆��gQx6e�>VzWi8�U�;(V��%�h�h?�������4�Rt�_���a�y�ݙ8YYN	��#���cif�ߒ;�7�ݩ�mZS�6I���Ӽ�n�y�v@�^T����4�g�pL�)0�ʣO@�.���z�h0�A���X5Cbv��s�����g���e��B�
�rz���g�/H����V��Zm][Р���E�b�F���r���3����>_��>�^����s>�7|WUԟ�t8������"U�|�'�M|�b�{d���K��i�+F��{)X�6u���G�3��A�KHW�1��%.2�E�k�hv@����A3��<C|�L��>�^��c=9ܝ�E!�����7My���J��o�x�=�do��-]�c�%�=n���'���P���!\�U��cx�fP�b����ڡ��{Ǡq��3�n��L��F�º�4������Gt^�C���f;c������t\�O��L��X�h9Fe�|A�r���X����BE��"J���;+a�;�{`�!̷�]�	��I��?�+EV0���y԰.��� ���t�d�c�:���� a��y?[P�\��.x�o�_Íp�f��q�>DW��HB��w��¸*�u.!�Nw
�TҢi����a��@6QR$�6���iø��xc�/̐��p �ʺ�f�Kk�N�d�r�!�N�g۵UlAR7�ш���/5T���I��i�ef_ @d�Ѡj�E"��$#�C��]��A������k��b�p�]O̴�D�Ƞ��T�"�e4iT-Nx��-L>���[��\�~�S�_��%������3�%��hv�{���x�;ﻖ��Fh:^��D�(����)x�b�+4ㄒ�X���t��+�l�����/j��X�̷l���]���vl���ݦ��݀YF�8m�*��-��#/���lo���Ҡ�\��谤��U��q�1*�V�)2��v'1��P�o��v��%�LE�K`3ٌԞX���}Pv��ȼH�V��W�ǡ.ue����bӬ5����dl �YW>ΟD����fYc��&�q���RӉ�c��(*�C�Jd��tA|���q�Gl�x2RBM_���� ȷ�E�|�6Z��,(��,����(T2��t����4�	�|��p[�4"p�0d�v]��T��l��~#¹D��q.�L ����Y�w9���r<��FE�ޏ�ޱ���]�� f���z����mb�����uKy�G���=Ĝ��Zțw�\3��3�H5|���!��5O�A׃�ȽU��L-�����oA~1x�J729����A���̴�!kB ���0��|��Ep'J�!6�����)��.��ªK;�n�G5�j2������W��Ԣ:�/g  DD�Ʃ<�/w�s����hC�=o�h��E��7P�\��r8?�[��_���������j7�<�Чb`ߡ����,�I*��#߽ �����2�e�`����id�=�w=����4�� �c���A�8�Z�\5w�E�B�?�{K�M�(����:Ka`�ƒ>e0��EX�k>�z�rM,��pH V&�%�v�Q͒�̈�'E!���H�����B��O����s��<rj`����l%GN�ۧY�Q}f)}L�a�7t�_�;(uK��t�Si��T�?K��c� ���`�Dk��A��N�N��X�M�F&�3�NW9�t�G+^�r�Y�JVc�uH3���������`������]�#�`D�0$�4���ϭ���� �V5eT����}k`��0����@pie��oާ���I~�s��ΤS�խ��f 4m<��sT�U�C���� �6J�<(湍d^M�]�C�B)�ԟ�8T��(̆+��i"�s�](Slߞ8��2۪:��L:JjYb,F�E�1�:�@m�*�µM~���Lq�&<�A�v;gQv�r�ݖBH���9Y�������-a��g����+F�L?6�}Q����mک�n�'���OG���OZ����%2��V������ ;�u��݁��,�=�a|��k-�?��L��q3�s�X#c��SJב��������
��ݐ����ge�pk�Ya.& ������K�dJ���_Ў���E����i#,�"��[�D��S�� E86���]4�XF�_!�+��4��3�������d>�>�Op7���x�a{;�.ET��e����Q�Q�_͓Fl�V/2�d,���e]b�o:�g̴�N���=�f���z6:�cu���q�y䘺�~�gQ8�W����	�`���N�\k�Xs�:��Yc�qO��	�4�50x��xpLZ&H�a�9Y�5�ɘ-�Y�����'+�M�Ƅ祱��U��5jH�L~9C��^%5N`��I?W��P}�'�d�%K���q�ʻ7�����܆+�D }����j�l]`��Ư�$x�ַ�H���H��YIo4-=�m���T�f���uR��m�Gyu�&� d�Anj
�7��6P$��D$l�O��!4��\%�LϬ�bH"�9tD����(�Pྌ�]��7�(#�jk����T����s|���\T$�XS\�n��_�f�>��D.����1�yCa�s��P+��x�����Ƚ,P+����S�s6��O�K�ea�I��W"eEv"���j T�.�3<)�OVy+�>hS#��s�����BP�����b�K0��
y�vja���]7�ˀ��c.����q�`g���J?��z���,��v���U��o��Y/�z��.�˼���3"pd�P�ז�+���<�	d��Y�H+P�{����K8������ExRb�LuQ]�j�~lx��5#�] Ok�M�#�������4����6XU,���'-��M��I<�#|,��qiW�[tG����|�'yܐ��T#Ls��1Wiqc%�	�#���f�Tl*��%�������$셤{0��	2����J4F!�~i��?�c�ӝ�	D�U�3�%��rs�@\݊=IWb"�;�����٧vR6n����4mȌ%�w&�I�\{�"���k�w�`���Ȗ�qʽޔt?�l�!��Z����1c��n`���|���ƞtI������x�[���S��"*+Yo*�݃�S�"��^��v��2�ջ�O ����{&�6�<��MN�9SS)j���1g&L��W�����RW�ύl$�U ��2/���:n�ͬ��Nq��dݘJV��~ʡ�p��)8�Dw��x)/׽���gE�nr�t7���4:��Om׼%S��C\�q�F[`�kdK�� yb0��d� "���A�?v}�NR��oxz�:1�+�)	���gX�ǚ�	������`e�rL�؂h�Q��U�S�t�Ђ�ǤnFG	�p�
Z�֖��篃)��q��L[���)D]��nu�K����hc�-w���b	\L�gLٗ�t��X�|R;��L����#��:5B������o04a��,>�%	�l*1=��s7�s�X�ö��f~P���.U������@I��.��|��|X�ܶ����/�K�_�DkQruF5mݝL"�(s�P��''4*Bb�����f��3Ó����b�ziS5�
����Ex	�.D
�Q�`��� \D��.ߝ�{�h��� :%�*dظ�Ai��~]o=,��G|�Q�ȗ�ϳ,-(<U��0�ǢY�$!�ǳ�����h���O�C#��B}ѿG�.4/'�d���d�/5��o���R릸V�%�,��xre���0�(���@�u<�(nG�?%�p1+yBIC�ٸ�j�R��{����~-ͩ�54��|�HoL�$������A���(Qh��m���}Bb���$ȬS�11������?���֒XZ 	��E�1���Y������*�7W�	��u۷�����X� x�i��z�]���O�5�>�º��?:☮\��,�̥���o��A��ۙ����Z t�i3���Ng�>��.�Tqq��#$ғ��A{p*��K�7�7>ς��
� ��wPa�SoN�
lȷb˞�����¼s[*�11����,�+�=Zm��]L&�R���ɝ:��}sʹ��;��u���/����<�n6^ρ-��b ���x��R�{��XM�5��"�]6�E,a]z��|�����<�T9l����ץe����V���x*��?:�u�K��-M7Қil3���b7�1��Ҍ��5|F�U3�=o�${:�Ѡ�����q��6'\]��nsV�����6��*~{	�ݭ��~�)��R	la3滣� ؝��E+�����@��2���Ŋ1�>r�9����v����^��l�#qF�E��*����~��(R%	�&�]���k{���+\�~�|��re5?�¡K�ps� ��P���/��L�%4��(y��d'�T+�=T��8� �.I7�[tnk)p֛�ID��hXU����г
���;b���.�������&5Бh�_��Dp�"�+we% ��be_���%�+� �g��ƾ#�@��U۔��L>�W#�_�{w������y���i=�G@�2���XcA��&W���|%&��΢�X���*b�'�X�y��,�������b���No�w%�O��g�gs&8r�#�z�߻�Ee��Z����&D�q4M+!��:b���M/�,����! �������7� ���m>:�x޾F�H.%DIl�y�Ac�����xL�J��� 0��du��,�
�AZTN�-�~�%)���jd�$��LHkM\,���O�綘�<R>��c�N?Z3� �"��q��go�z(�9�\��w������Ǖ�I�	���7�T���r�q���u�s*�ǶAe�D�򭰗
�5\S�"l��ui�R�Fm�H�h�j(\e.��	��d�j�.��GG?9<�s;�����O! ����RHP�'�&�fp��y����A
ҳ85CU�nM��N��E�=��t~�>kG�Qvηk��Y�u��ZdYޕ0�ϯ����d�u���◷�Ζ��Q��9�@5�z	uH�oa�����M\ �U�ٿ�^�&
�.�qB�:�2�,"�-ZVl���%jIQh4h�s�L0jު�b^���%��q����	~�>�2{C�qG�uVdj�����u<�6QFT�[�{�	j������c��8��6�팂T��i�l]�#�MB$��x��[��A��^�E�K�ݭz�f*��/q��}�ziY���EUH33+��ݖo.M�O&�IT����c�(�OA<=�4�c匬���!��7��)q67}��ɠ�a�'��8`f�-��C;�������	�@�w�) ���̏KW�Y@�����s��X�Ԥ\=�
�1m��M┏���^�g�DS�o��!��/t#�'�6�:Up�#��' 
�Ah1NJ ��4��#�_�M�Z���+��d��8�
�{2��m��r*^�03�UUq�� @��͓��=�M��s8i���>��(�?��A�F�$q��4\x�B��.�����F 2鍄9X�\ha���M����o]�ZU8S���z�M� ���w�
"/'O�2&��\����uV޾F���/;\�ԛ��+��|n�ι��\%�]U��C��,]���x<���*~�-v�V.��f)�1DX���-W���d�3l6��\9�8�� Ų��k��\ʢf�Av 7h=����k�R3h
r�6�ϲ��?	�A��G����+�Zo��+B�������U��` �;���_��\��`A�)��Z���TF�����Fl�L��*RVW�qF�׋[3�>�Իe87a�;��X�>_Z1�J��uk�� �6Z�k����ZHhp��T��G��a+���ȫ���:��}�׉%վ+v�M���]�;�Z�=�Nbn ΙDh�g�]�&�+�YW���9��	ݻcB�(qE�\�x�X�!�9v���~��)�1G��/f%��<>$��F:�K����l����Ҩ�nz���\����v������g[��H��nCUQǊ�l��<���l��j���v%(��)�a	�KP�ν�ǆ���o�̡��uʮ`��� ��o����@�fzN&5t�����WDі���jl�t)@�L����;KQ��:PQ��B��A��k5H�TÍ���]T��-Ѿ�^H�,�3�d:�����B\4!���tv�	�[yѺ�)V�ў:9v�1/ j=3n�Yi3�-z��?�����C1���ra��xc2Z�������K��b+��j��w7�T�{���[�5e��oHf�Ȇ�E��wl�q��#>Ì����}P��SV��(��՘�S���'ǻ�؂�_#a=�,%t���!;�ľ��h�	�Dk�5nX�Fn^����D����	��	P���o.a��NY�~|w![�R�_.��)���%�o��1����?��Kw!��u�����A����ٗ�2.�����rd_��5
(8b�q̨�/�Oj3���4�mz�|�!s�B��R���ю�/J3�n	x�z�W�F$�]�8��N����A\��mxK�������-���H	��H�b�� Eo"p=pe���� E�L��*e&=�}����RaeQ����Ju9���s��@�$(1�j8_u���]8��1.�O�{���(w�I����5#ݓ��}D��Q������$m<ntl7u��_9R���6BJ��QC�V�Ae�(�]��J7�CQ��P5�l���ol;��n���q/i!m.o���b�2���F��ICtV�&�)��%���{W'[�2�_w(�7���:�`�۞1��]�YZ�'��j��P��+U�j:Vw�Ҥ>-~=BZ!�$5u�����%� ٫i_[���`�g2;�F�µj�� ��&��QeO��$�2��z�yVɤw�o�C��%�ed��6!g�����Zl�L0�f}E}F��A}��og`m8�������I�b��2W-���0ǚ�W��?Ӣk��A�L�yH�V�\�
FX'��,�"⡓�T�ĀO|�K�Hr�.����/e� Y�V�4L��;��-�%8��P�N�JS�%��J����|}<�Lu�* @������I���)MS���OOQ=�8�u+$�Ҭ�ɮ�3Y����- 2@n<��v���	`�I���A΍�Pe����Fqo�*���_���[ÿZ�1!֒u�������jwbI�w� 1�v oJ�?�j�t{���,j�u�M����9S��yX�P��R����kp%�� �ھ�����~�`cXf��.4�؛�A��}��r�-F\� ����vƳ\�c��j��[����cO\��{%�f�]4GOc���E\7�|P�
[`$\�D�g�͔@sA�(�{K�P���R�6��4ɨ�پ{���WU~k������{k��������z�<6A�gPp~;^·t�U�u46� Dg/9�&��2-�W��U���u?x.>�,��ٙ�Ǉd3�q�Y�uZ�$�R�+���E�!�I}�Q8�J���?�p�҃ac'n ��s��P���Ɖ�U`�F�i����ط!��P@w@Cﲙ�7A��8�`�pLb=ExD�����D˄0&0E=
���X[�^�$p��j�9�k������ul��1���,?�}"Jr��U�<���'ǏQ"�^^qs��X�b]$OV��MP�Wie�H�'z~'X{n#���kͪ��c�oS����H�HJ�1�%ؔU��!�	��_,�ȍ��I�<�5+���+����@�2��u%B��&?^�:�����Ԯv��EH�Սz����W1G�oh��n�Ϧ��Z��~fP|�j����z 	�����k�����`��gi��p[ 1ގ? �''*J�eG������ϖ5I���%��U��&�"�B󶤋�����sluϽJ�f���"��xA�N�z:&�,�eu���;�*&���J�,����z��º�|
��TPapP-*�����aR�=]��t�7���/7��'2�%�x�Xj�I�����}R���]��6'�(����z�>�\��ԛ�B��yv�	]I�q#�X�y� ����98��#3lO���H`N�C�(��Ʋ��Lk�u!��`�F���p"�V[%�6D^R��8l`�B����x�aqR��[��KZE���%bn��v�{�l}��)"���R��x����,�4൸��ѠG�HIW����d��rAho��zT�����H/w��5���-������ y� l�3M��
u*���x����jmIjx�ny�(��*�>���L4��!%�X,���J���OE{����#5&��˯�D~��ˆK�=2:�]!j�S[��f
�u�����Т��|��%��Β�S�"����.�5�I�0b�QX�L���X2u�K�*�o ��φ���1U������k�Ts:�z��ՊTӊ�bc���y1��~�4��/VU��*	�;�뇟J���T���p�|��էA�,�Iη�@��{��l�9�v�d�0�t���^B�VQPB~)�k�y�~��b���+T aw6bm	锜:Y��y�y�K���ȅ�Sݕ!��z�kh��/Q*��?�LX�׼��������-%��}�oS-�	(rNH1Ώ�p���]�"������bs7ϻ��\���L e �ϵ$�:63���:��n[�A��p�S���jBy��㳥?�Lk&�m�?�j=���LU�GO8�/')��;�~A�ЉA�'v\p�3ws~��k�;1.o��_�NV�b�L�d��Lx-ޭ]K��t��AK���m{�2T��d�����d�� �C����x+;T���g�W��y[��y^��2	J���uX��PM�^�>���Ҡ���T�L��zj��My�+ �,��3���_^C4���C�6�)�ɏ �Y�p
�^x)Y�b�,�y'6����$dv`��Z9W:Gžq�w89���]��P9�����Q����c�����&4��(E���?oZ�x�.,�k|���'�E7�;$[B�H�I�)o/Z�.üx�ܾ�$*���I�i-�T�8��Gܫ=E�/B໯I�@V$;%s��'��������g�e�T�<G�g����[[� @���r{���7j<�O��T��?�J�����!X�Ђ	f�y���ׅ�� i���5AhK�l[�k���}@+�qK�E$�G	R������ ��p%w2�������rU�c)<���@xZ=!�W��pZ���Tv������q�����*��1/�A���j>\�:=�;�M�骸l4�L�O�9�"��Q�s�s�c��D7tE�2�I�cc�eR�Ā$���m�mFz�?{W�:�_�#�C]��ΖF)-NV}�l��|b��>���>�.��{��p��C�ܔ��x_��H3�Ѽ(HU��Z���zۖ�fnՁ�)�
�� �ZF ��iܛ>�6>��"�1�p��C�UeJMЕ}E�"iˈ�j�6H��|O>��ڃ�@�ȡ�q��nC3��{�+o'y��|M
g�%NtN\Jl̵�ʧf�_�w\��a�ߍ�5ue�b��^�L��Z�Ln"�9��؊�x�@v�6���J�1�RX"�'��q%�p�덳^��W��_���Am����^1Ir�l�M�[4�F8����E� 镀�� ֩[�h*�*��X��*��֪z>s��*3�?7���r(=M�qL�NP!!"=���a@�e�W��
�>���:0r�;r.U��G��S"B(04g��X%�YNbg�B��Ѷ�20l7B�t_�+PD��g��y.-4/�������)	G��i��m���s:l
R����n~����	�s�98��Goj��		?Q�wJ��ம;�_���;Z�ʕ(!�2�Z����i�e!�TD�T����0�~�mr��TՍ�,���-��[���)9ʱ�TLJz�*�y���"5��y��]����Ņ���ɈU�~�<�D�X7�Q^�T�d�:}�8�+�&���f�������%�J�J$0��gQ�d���w�"��Thq]lw�I��#4��k�?냾�*�������fF��O�A�>��� v��}V��a\��\�Vhd��K4��5�7�v�u�J�Q	�Fs�|�D�;��Ou�!!fu-�L������rC���<��s����8*ר^����l!F��P7���?Y�K�<d�
��bI�}k�n�D�t.iYxŨb��9,ը�y%6+��R��С�%?bd�&ǖV���K�C{�����,"-���(	����W�(��?����!�}��v���"=]&�LOѴ����K�+�ǿ�r��Q.�O~9;�v�yX��1>�j����69�v��<J��-U�hŇ�����؍��2+��x�Rt=���	�&idS֪�K�o��iO|R�_z��%5<���O�φx��H�F�U��2�Y��U`>4��D��$z�!%o
���8�=v�J��`P�� �������"�޹l�	T�W7/��7��+`f�T#��'
�(���;�u7G����S���?Y��5����TO_H�3[$��=kx�J��O�qR�q)8���� H2(s�
*�$
n�510����?GWHS�fv�ߵO/��W�.����at&��w �bn�Úl����}�3�醏�C�U���c��wJ��L$ �������� l`6�a3��Ӹ�+Z���d)��CrM��F�?�*��?�����}N�7]��F��i�zZ��h�&�k�soDU���ۥ9̈� �Uז`��E���G��Qu6Ϩ�m�RB�`F���5t#^Z�����"�XȔ��~�5�i��E��ݬ@Ԇ0PCC��0,эq�(�AĤ��%c�W��A����	����sյ�\��8/G��A��}A Pr�^I+H�����^��b�s��E&u�\3I�Y�%bO�MǔP�y�y3�D�����6�#"N��+dMd�U)uXS~�ڏ�fF'�dE�(�zK����H���+�"Ϟ�:�΂o01���l�'ňc������o7\�|�����O�X��*��E1Q9(�������1p�D9F���$l�óڗ��e��[�KF�+��-�t8UYY���C�<:s{�{Na5ҩ՗���HǗb���������rd���:����y_[��^F�al$&X
g������7��է	�f�Ux޻=$��x��a"�?�� y��ș�=����JFKy��8�qx!Hz_�n����=�$v��Vz&��)�r��g��<�A���p��	���'���3t޿@�����+�l�A�K�5���I!�r�7p�����̱�t&1Eg�U �6���HwO��\���(=����D�̸cTR��� � �^Js&�� �3�a�}�[�j��\$ѷ�N
n���[�VF[0����*D�4��^����r'J���K���DS�iϊG�����5\�c~P�үl(^׏�*�,C�{��gM�9[��.°��Jn�׮�����^��Y0�QX��/783�Bf,f��72^H�x|w�f�{����@Tۨ�ݘ�E�D�G�#�K�,P��W�}�?e�#WRC�T�=��ò�^o&Ͳ�Ux�F�OlYOve��G�~�d�P�+Y^���bn^��^>-1�;A��F��>P�8����!2j7���=n�d(i�J���v�ц�° jDu*+����+��~����<qD���$Zy�Ûl��v]z)\�*V�Uϰ�o8��̻�h�ȗ32v�4���t$jgx���X���0	�����W}�5�xPxdl	;����R�f,^>�/�<f�=7'�6+�G�.;�KWV�����p�L<���V�;o�
mĂ�T{ѩs0����������8e�jal��o@���T�q~���ߖ��Z%��;�qV��%��������bmr���W��h��G���ǋjwgvH�6���e6q=�ƒj���se�����`C���
�Qo�v�^�.�_f�a��n���,x�#Lt[��b@α�<0S���\Kf��?T�j`Y0��g�-j���8m6,�b;�2ӧM|S�b���#`kd��7���f{��?gѴo?k�w4�)��H�̑��Є�[�S�\x��V�Gw�a|Dp:��xS�_��`:}�֍���n�B�[���PfGZO���Q�^�@.��ϩ�0ܛ�8�g�@����є�g2��D����A%Z�I�P+{��J��c��}յV�� r[Nz��p+���rA�첰-&�|B���3�Jُ���]& q��a9��#�P�ߜ���Q���ͬr)fEiV��%:)#��Y�����P1��o����Dl�H�_\(L�B[N�y�O����JcH�1����-8�U�ˣo�q�?ՈU�<˪�>S7%�:��f
f�w+<Iӓ����"�ʜ�0�u&{}e��\�]�)S!��s�s�/�΍�����V�{3R"!���"�e����a	�&P�>b��h>���Ѣl"�Q�7Bo�8�q��с��:�����`Ud�~SJ;бaA�Ǝ�J#���2����'
F,BM@���&�T1�JajGq;)&�L_3�^�@q����oA��G���0-l��8�%V���_�.�q*x?���^ֳA����q���|݉ή�_���-<�AM!?������?��g9k8Ƒ�>�� V�#���]�iu2u��:�2���h���l6�������}�F(=_�� ���j���t�Iw��-���\
��Wq��|Kg������{�)�zr8p՞!anB]��^R�k�lN1���<��6ÿ���:�!�W�{h_�\{J�ż� #]�+���R;�K�8�K�YK���&K�����:��N�1���@0fO��[����~y
#I\�2-*��3�ӯ�	���H�XH�:{Wb78U�N�z�>*{d8[#�)�	s�T)�j٠�.v �{��L%>W
��G�%�2��6U8�g��Z��f�v��ٻ7��lHڧJztzՖ>5ۼk/���*��a��9�e��^�����^�ʭ��r�����x������^��R
����FƑ���ŻX�$�]y�.�L�l!Ѧ�����b�a%{�u��n�G��{�=}+Z����	5g�b����w6q�8�j��ͦ�z��n����AL�Ϟe��/.]V���*VK��6�6�s�!K���?�YZ:<��@ j͸�1�/������1�cߨU��4�{S9����髾��NLO�U�4�W�k{�_�5_]���n�\CR�G�t2&��+�<p]4.D=b�	���S־�g+veU�Vcs��~=&j
x��� ��W��
��A��q'|�g k�I�KU� *�Ll�Y���-&���ˀw&|\�k35uՉ#@cur� C����>��T=M'lZ,P�r�l�=	�.趻	νŀ.�GB��=�z�2��^_�+%��r{
�̙�"��Op��l�6��%~&��C����@�7��U��:�Jh쪺�!�!����A��V+��>n��v���G�H�2�A/A����=v�n�v*N���y��fK�ֻ߲�
��:���Ľ�#x�͂�l�y(�fegq:/DI� �s!iq�_��i��/��(Se(]S͘|�!.bbظa�#��`�E�`�VJ�=�e3^�pTu9��������︀l��bN��Z�-�pj�Yz��i:���#1zFk�֮m(ci���O���w0��p�IЁ�r��v�\#�Z�B�gD����t& ��i�t�]��K4�g�SnŲޜr��R|��_�ʂ�w��d�;^vYL��0'5�i�W�}�\�l�q�2�T(;e��t`B}�|h����������n�f���j���}}C���	��gbEa��;qT�}R����P	6���u\�M_rC���{M!_G����W���TC�T��1�*�W%H�
���<��_y��#o�rM�4�V��]�3�0�~|q�wR=W���V,��N����M}W���w�%�ڈx:(ܯ�-��T����6�Μ�e0�T���R�q��P��]�5"ڳ��J�(7֗���-u��_�x�\�t}W4�
&[;���p���ѣAӔؿ�S��5�OĹ%����={�>SkW�=>��tW_w\����y�$�9 ��X�t|��-?��b=&��㪪�����;�zK[�.�q�4����*<��F,{lTB �$�/eE&?L�zX+��"�	ǣ���߻��	OQt>�tA�	��D����(�[ WT�JVR�Q����W̆��s�e>�����ڨ_e�B=�ܓ5�[]��+&�B�>����/`\H�J���I.�y���r��.�.j��5!�2q���%��#�>H���~�q�YO�j�ET�����z1�Z����I/uU��*U��}�Xd�j�������������q-�[Cu��O�QB?HgQ;K��ķ���e3��� -�����x7�$.fZҚ,�8ݧ2��$�8/����kG�
���Ԇ��쯿}0G[���	8+�$Ѝh ������ҷ���q)� �__hL:��T擦%�R|�����}��˝�2<��c����BK:F�`+f�xv0B � &^~�"��2�Ы^����*�6���(���y�'���i���K�^L��I�ơȣI���m����-�A��x9���m���r�-hٲ�v����@b�ҽ-x,kngp��$��B '�TU�}��w���X��ǔ��P�4�;��h3����e��F�:=r4uJ�A��+}$m7M�~U�m����-���*	R��`݇�>��z����wx���Յ��V�0�V�<��MN�Q�H��s��7�{;�/���}.��=����Ѵ�7c��� ��i}��M�Wϒ��?��W0�f�,���3�c(v��~�]_J�U��u����U=�kۄ:��޿�x�S5�L���h����s=�\�n�,5�Rʪ?��J6���Σz�����9�r,|��gVA�PmQ��=r������O/R8�|��._H�6�7rr�P����'cm�n���QHZ	�z�-���+�q��aj\}�b�M�}+9�����ܶ��#->����du�0N��Z
D
9��zr�WT��º�f{�]���x���2��$0������I"�|��-�u��u�4>�>+,_����)_+��:�� �©Jq�S?��첗J��8���uա�;�����&��8_�:j�4N�6qp.)�n^�dO�84�Gr�U�_=T��M1�M�������z�.(�&1�&�����?'��&w�?D����'��2-xK�����ؖƓ�z¤�K#%��{
��B������������]7Q�CEH�U�"�eK�|��Y� W���|j�fU-�"�zc�����yK��7��;Y{�l�w�<�7�n1���<�Zt�r�u�1Ia�rE�/9��w�pO��Xlbr8T��}&���.�z�����&��"j�(
�~~D��A��`}�&�I�z	y���_�<6m<�R<�j?Tl��w��6��0v�:��Ѽ�J�KN�� �m1�q�
,۰-dD��e��nJlG>�v9�A�;-�dr���m��$(h�]&`�4բ����WP�z>�כƦ���KHuPT���o*9ce�����0��'Y��>?1���2�4�s�q���*Y�3�g8~[�'�^�2g�e��{u�������.��{���E-�����e{�5ϣvڑ�3���vp����Wf���@�V��k�M�֕��C�S�i��,��^�J�����0@��V�6�����;�{�z�^9����3a��]�*W͝n�Q�b
юm��)У��^P+LU�械�.vYa�k�q�K�%*{O�dNJ�e�\����@(T����W�5��,�"Q�֯3���w"<��O}�	�So�b�C�CA'�H���-�z$Q6�z�Q\�n���bغ����QE"G� 9IS��ZZa ��t��b�HJg�^F�4���?<�n�Tq�m����l�o�dd�	>�Mn�IknG�H�u�s����JKŅ�����g>�	rG8�X9�ms���O(���d+}{<g�|ytH�H�K�ŰN�\q�`��v��GYa�D��Ԓ�rN#$xA80���+�.đ���
��R�1 X�~-
��].�5<��`�2i�$�AJ����cyXG(�AlcOh��A[ȴ��w �^t8?�Y���3�p����1�
�YPϐ�#H�.4k��Vk���p�p�r�+
R�L#̳�ô�:m^��������_��ڂO����!�*O�1��j��\|A��!�햏9n�kc�0j�׶�¥P${QS$2��x�<^`�+���v�_�ػ�2�l���,jb�8��l�wF�԰X6�j�eҔz��*E_r�������A�얃7�� qc�ie���v�7��k�*c���eW��WK���-nB���Lie����#���Z0IE���b6T4&����!��l���z��W'�rL!:~:��f�[P�?Ԩ�v����&����)[舑�"�Ɩ(���'V����ɴ>���5��HK�	o(�<(ƏH��F��=g	��C4����7�H���!�b�KSZNL^啇�Z�r�̩�rq��a/D�|Z�y3�_!�Դǽҷ�
^��X�]�N�3�Sy�)Y�Y�q��/�+jx��W�7��]^?˂x�ޡ	���h�~��~�����E��`v]q�7s�`0rK��i���\6��8Xp�9��N�&�J���vT� �`�����Y@����;8�;j�=�VGBj�mk8�'b���D��ON�3D@�M��{�R�pp��7F�qkn3�"�דiΥ�KBN��MGV��3`��6���r�� �ew��Н���6�f��~V�ki� ��Դ�g��^�9A�J������qJ�QE�_n��ᘺ���V�y�Φ~���U�e2;u`��ð	m�m���p�h28TT-ímΡ;�:^�z�q�3���)�_JH��oÐ���`�j����wOi�w�}�?���#!����x�Ύ�ؑ�.�y� �w+>G6�	��>%N�y�n��\q���|K\�D/%H��j��Rd���"���]i:Aw�>צ�<Ȑ�t�� ��꽔6���)O��Ls,�=|�8�٤V(�.*�`�Y?Z�� T�����6��G7X�Ñ1���+#��A���H�����o&Ti���>A�b$|*	���*8��lthf����#����gT�%屛ka&9��)�O�j�8�~
�<�O7X��&n^�6����W�Bu������V��dC�)C�a#�-��yW~{�t�RP�KH58��*8��®��R���s<��ܲ�%���aބ�l�k���Y�Q�L���Fb�<���]�,<��Xz��V9�¾�����g�S�s�e��D�0
�Q &l��Z�ݚp��b��P�E�(�IP4kaD��#<Z��j�|�aY�[���A�����B�17ɦY�X�<���K��-�Kt��-X�{d�'�7�A�H�
���D���=qB�K��,sQ�2-�������)հ��2#�����A���UMj�R�U���9�����ƞ��Μ|�:2�^�{�
�ꄖ��o4��Ǝ�����1Q�6x�9Z=��̒8�Ǵ��7?�X�C{����0�ٹЊ,
7��IJM������a���fr0K��b����$��u�L� v�^"C&�?�嶬b���BΧk�d��X��[B2�j�ӣ�?��0��Jm�y=��&��ln�=�;c2�l����\��2�Y,V��{]�MEa�O=b-� H�ƶ��r_n$�
4�{<se��l�vC ��m��O��]*H��h.��<
�u%QK��J��� �=���c2�A��N]M�:H���sC�V�c��ܲ9���O!���pk�U�Ώ/ J�ӊ���a_�������Ϲh�*����4�Blo������s ���V���#J�ɜ��I��e:��u_�Im aCݙ�+����]g`I��H@�i�ri��n-�no�@�hƱҴ�ɭB�8���"E=̩Ԗ1��P�G�aH΄���}qX��Ӈ|E����w'�ps�^x��l���]���R4��D�-O�8~�f�LĕӨ���i+�@��Sv��^J",��8��=Xt_����P�B���O��I�{1%���.`FE�v'�d�B��6�dGUp?Ғ�T#�sWd @ �fq�q�R����#�W��1O��OaܮQ�јwB��¼x���uL,������ΰ�j�UdƢ�ΫaHf��Mk�8E����w��Su�-Q��c#�S�,7[�H�=`e�_�#o���Q��<�ԧ8�|j���*`�v��^������&��h%M@o"�L��6���O8qK���YR4>Jc��Q4%�V�J;`������C:����q����N�R������B�n<َ����,�D���[�8��&U��y��,>��8�r�Jv!�]�5�b4DW6�6&���bcg\��<��FY�5�l|��2K�r)�*�I��u�f�{�A%�N��R{:F�`�ƣ@g�w^{�#>��1��`��ȹ[��^y��t|�)w��n��?Ǚ�|�|�$8���^iMO7i��,��1���.����;Cxz{�LbR��7�\7��O?<Dо�P�~���oj��nx@��V�9i����-u\9���!>�$<���Y����Mx�,�*�u��S���rk0������A:߻�`3�5K ���	-��%��RK+�zc��=9$TO���1-�c����eKؐ��Gӳ��QĉCTc޼�/�K�c@���L��Y�+��/�y������0�w��W���r:�nH5��rj#Й��<@���*.��V����|#��.@Qf�~�_Xi�q�<��ǁ�PX�Fz��挦�j^5�x���1� ���� m

�ߩ	J��_e@�z��t�Ж��q��>7%��C/���H�	�>���`ě�Z�3��f��������_j�Nyz��u� �����>F=��0��\����Zw��A0��Wn���Ճ@��� e]��.Wg{��J�*���NcQ3��s�{x�T,bU�x���;�Om;�E�b)��`"N�5��\�"X��b؀�]@�K�|ԏ�-�&���H5 @W{k�x�M�E �o0j��`uN��J��	uH�ZV�V�[��J�g�ī�O��j?��� �����W���}~P����K�r�=-�޻(�@Fw�eݞ���kR�tǌ�q��J��Ա �95�d`��۰y`*X�.��!��r�+`����z�,�;͈��@daa^�A�M�:FxDGB��Ƨ#˗7#�B���y��~��V�ò�����G�P�����!4�/2�L�f��8��'����}�~ꆷQ{zD�ճ�o#�MV��^��	�H8C
��[~.�R�j����b���V%{��Q�l�p���K�;D�؇R�����
�D�J���PVp*��9�cL�t��>/%��C�@ܾ!&Q�9�`7�˚	�^����#�C%>��Mt�>�i����(e 
w| t��=�Q:��Kh��i!�糤���)��i�tn��=�Vq`��2h�Sw�p�U;uF�Ӛ��>��-U���2�n�^v��q	�������Z8�\޳���kr�2L����9���rug5	�������b�"�xT&��ﳛ]ѷ�!�x�������~d����7a59���e��c2$�I�;Q�B��>�ɴ�^Q�U W�4DӐ�[.Dd�u&m/0Ջgj��1��P�X��6L��d�c���r��'� ���.M"�N�y�%Mo���8*���f�U#W]O���.��3���ɖ�gG¸eT�o|{���%�6���xO'8��WPƠ��bT�a�����lp�\O���;#_A���]!���y��m5�i]�%�y���Ep�qKa>���!��Π��g��+�(	�VA	qg^�bK��1�wc���b���n�L)�cx%:�,� �:&�B�n!��!��c��)'0k�����B\��&i���`+[.�����L��d6�����}�$D�\ᄀ�[��,1��0S)vt���.s`Y_���F�;&ۜ��S�ķw�^���gH��5��	�XhnS!�$�,7x^�r�|�OB]3�j�6�6H?R��(e��J�X���׽`5�,R}��ӫNi�~�
S$�]����)��B�ͣ��{�~�CN���K��H��»!�%a�ϴF"p���YI�#�	��*��u�׶�ņsO6����D�cڜ3�b��J�=ɩ���Bd�uq �M�pIH�qjx���N��sP���
�邌��;͋{exd$n�q9�9�Q�π�&i�|w�uu�����.��.�[��Rhɮ�;tc��̩���'���c���D��u�Gm����s�j����m* 2<ؔm������>{������;>���`N���ExdHv���E�C�(z_��%�6����X=@'�H�G�!����I�t���wD�k�6|%���m\��a�����������V� 䔢�i+�٩�?C6���W_[ �A	��G���yT�eJyd�N�j�9�	�$��P �\����[<������K8��p����.G���atth��%�m���=��ySO�w�	�L�D�Z;�gh�=� D��^�^����c��P�M����O�I�,��y���3W��_���O2�w E�^ǋ	ʭ}�����Q�Q��'�ڀ��8�O��Jd�6��ĩA � ��Sd�I2�ٺH#΀��~����=�c;FP[	�]* ����6�d�5a�sq@z��&����O��e$�u��`nrN���.����f�~p�<�KCd;��=���na�",Ϋ�b��R���.n��`5GM�؊.�_v�Fb&{�e{�JP�d�!�.1�5��,��C��h7B}o�ҐqC��F-f��?�.���m�V"��+�o�K�_�=d���u��5Yq��H44q=*k=\s�^�z�;��Az��	1VZ��HIOiq�b��ܐ�}YD�Y����[�s��ٗAݾ ��X.Ў���oaxO!X��`�����Ơ�#A�ع���[�j[�%�֡����>�#��{��4r(��XMti�^�]E�k�EN���*]"�M*��T��u�l�C����ĝ$��?-+�	8�`�!�ݺ>i�a�}h�H-s�T� !��
yG`#�'����O�T����_�S'p��@�����`����vF��f��4�+�a��{B�M{vi�U��c�sh����˅wz���=�\m[�%����2��H,��rw����8T�H�3A��i$b�X�w���9�K�F��v.X��~��6�g��s~*�l2�RP�}��[�ħ$����?ثR����f$�f#HO��#�H_&3�r�_w���>L#b���S��@���ó�F�%)�g6�Yx.��]�lT�I��N�r�"����]���%f���L0�5B��Z��hw��<{�hGK@m�A�ːˈ��`��JB�`d䧴���o����'B�gy�~z%M�M~�e O����c.0G~��*���GD�Hk�6R�#��xi����yjZх��6�P���Ts+�s[�B�Y��'0�m}O;e����;a^��M(e^�_��#}��'��˽�!WW̎�6�4�"�y�dF����~-4��\��� ��:�1Ʒ6��
"f�+�:C�W���|����Ƭ+8�:fn&�q�A&�N�5��E������C�6[��W V�R�HP�n(�؄�<#�R̭0��1�®����X�.��pj�#Ԕ�o��2��}G"|��W�"�4]x����P������ٳgW{�"Z|�Z���}*6�����V��<��9�p��"��oaܲ	�a����ҥ��&6��b�>q�� e��8=���5��XYj�[bW���3BQa)*�孑J���[��� �G`w�h��p�Fa�!*�=�SqU���O8B�xA�n^*=�7� �0���HE����ՁQ�;
�׉̎bI������Zz+��׿�u�m̑�M����~�J�9^,' w���1��c��j�s�%��5R���0���<��uB��;����'�`{wU�B��o��i3�Y��8t��_ʣ湆�k�iS�H]M�Q�xCD�� a�x)���s儝��T��	�aV <������b��n��VS%��x�s�m̗r�t��8T�puK�8�,��n���J\�F�i	��;݋��!.;A]��dkM�3�t"�|p Y���� hX�`+�G0��&Oǥxg���o��~�y��Kg~�r�눷T�����k,;Dq0��]?^�԰T{�$1����XC�g��h���f�R*2��o���s�LĜͲ�	f���� q���
gœ�' "��S���/�\?c��B��
-������Z(�h�-Rk�kZ@��QͪY�C�k�MV�<�<ic-��&�5�j`�6�אQ�i��B��E++A��W�X�����TX�ա8�V�QF%ǧh�9��h$%?К0��A���N��H癧22���G��JUe>��!(̺2�G �y"�y<+`��-z��^�g(HWt�D�H9�����1q�U�ap}�a=� ����C���Y��mG)�GI�dcq��u���QZ*�y:~˂G ��A�ˣ�ޢ�n�|:�~~'J즞B��fҫ���4��2>���x��8�M��A�l�g�m=�`f�A^�����"ΫQa���jT)�^� �:�]�4�F� 9R^���F81�aS�Mr�,�ϵ��p�!GYm�,���P03QZ'�3=8���
��ѠTO���>��).�.ύa5���w�����B��NvG�7�`Nò�\��2C1o�b��[�rs� g��pg�jgRY1.X+]/,%��E��w/z���l��NCK�"r9-X&��=H!n#]
���f��BKMCцf�x�R+� ��>D�$��tY|DJ�Q,2=�Y-���6�>��pWt	31�Ky���	�m#�"@*xwA4Fj�"�ϫ�/=��i=:�[>�H��a}��09��;�ȏ�u�nz?��������^�4��cF���׌b�9�b06�<)�Ļ(cLʀ�9����	��|���\&UG�F�]�=�2Z��s0"ݘ*��Z'���o@�6Jt�	.�.W�)�\�>��	}މ���g��3��Rd^NNP�[�ߊQ���V�bN���A�(~ɜG�c�x�R>�5f��#6p�]���3�sʊ+}��
^�_\;C�	���F�+ �N�oo��I���¹Q����g4�&��o�꧿s����gm�<�T���w���1"��xc�o�>+)BP�Pu�����t��bafNZ�R�g2�D\��t�ޤ|��x�!P� g�| �F��=�)<a��]�p�b�������B�⸖A�h#��Վ=�}B%6����j/���
po��j�;&L������$91E���uᛉ�f� '⬗VP7�MF��M#-,��ۑۛ^N�s�6���ς��ν�L�/�f'w�8����V������+���q�j���ϯ6�T8��C@[=}o��yH�m�����L{g ��GuY�B�Ԕ�	ZNq����~ԯN���T#�PT��fo\��ВM��k��ajRz�䎀WZ���dIߐÓo����0���VH��- �|z��3���޼T�P���PjJ8
T�{h�.65�S.��[8����O�&a�І��I������r��*�v"4$<yEZ-[����{ɰh��>��t\�}iM�!,:��$�}��L����f��?�\#��jċ�Z�n0<�i<�*K�Ȓ��"n{8[��ɪA��#�d5mm ���"���<��N��*@l�ckK��$��;�d$��2�r����A�%t��9-(��c)/ϻAb�҂{!vnݴJ�%L�	\<���j����=�v ��ٌ]��0P�+O]j9
֙�@��t�?����I_� :��{�`%`�븵�#Y����ܜ���jo)_W
��i�� [ܫ	��G"�m	c()�57��N3/g^�p�I{�ÞuKG���n�r��wze|H �"	�`4,)!�~0���U���D@6�������T�g챖�0_�4#t��;�A�J �1�/�B�
�̛3��VYG8���������]�a�E��U�����6�������yj�����Fg�dV2�]r���U�T�дObfڃ�e�����>ݳ<��nF���,�� �1�*O��f8ɋQ�y툈�{3�w*����O�q ���-b_�����3�t>ƿ�<���.�[�on��?*E����e�ڜ�)aJf�0��&Y]�M���S�५Av���uR)ohn��aCN- l FLg�A���J�.�:ƀt
���X�i�n֌΋��"�y�s�0J���G�l��(�"�!�E��^|�	�#���M�3���W�� N�n�[
�fN&���ί鶴�����7�n���g�tT�^�6r�:�ǆ=Np��9�:���^@k6���m
Z�P1�R� Fݤ�f�L�e}a��n ��itL6��(ٴd�z
�\h{lV�8b��8��{���)��8k7go�X0��	�et"��76VxRp�m�tx߳�W��%�k/\\:q��W4��qU��~h�!�h�f_]�v��<��l���}:�ԳK���J8������w��ky��L��Ֆ'��c�F�N��P���🕟k1��-�iRP�Yb���H�G�k�gv`ҙΫǨ�����8ȳ�\��4Mi�*9�,�뫱�e��q<��`^&N��~�6X��Z@J�7�1"�0_�;�q�?�,P~�T=O�
?��o���P��i'��ӑ����VU�CvH�	��*M0��B5B��G���pM^0�!i&�/����,�����j�`Y�݁-�;ZC7���+�4)���B m�đƘm�'C'v�#��RؽƀL=U�XF=@@�.:��R�'}�fڽ����8�����?��Q�'3�Hag��n�H+"B����G��-n�\G/ơb��{Zv��4��<��m}�<�a|��wФ3��G����.?�s9�$;u����'����cb�"����~ȿ�;��c��q�d������1����)��x6pPJ�Hɽ��	9r�LV��s��,�G\�������e�|!�L�|4�ӗ�Ln�����pߣ�LrO�o��M�������:��0������@4���n=�Fk�6?�K�Z)������8��	(�̇��B[6� ?[��vT��T��L;�N��
,r�Gב���LZTv���x�L��n�G/erB�~��k)��P��d�-�h\ɪ�7R��D�&�.�k9� �,��vO�Q(Ӿ3N�::^������7�Ⱦ(���o{=1d�Bu9�Iq��3Jo��m��"lƲ�V�<���{c�8���ƚ��-w�!X�l�\}��R{af�U$3�I~� 8�m�Lbc�����[)�d��S����|��Qr����M��χ��5)VȆ�P� 0��otK;������٨i��6��ɦ�C��.��RKُcj�:�W~YZ6�>4x�	#�5Fۧ��1���mЮ}X�J��Q�jk��r�'�g��;d'
лپ�$�z��8�)�l��L%X���4i3�eO�~���`�=
��q������!�e�\nw�KF�����E�f��(P}b��ein�pdM1���±�"K�(T�����(�� {���Ɛj�?d%�c/��Gְ�v��?�,��Xb�ĂI�S�="a��(����2B�5�Ob"\ë��A�$�0���z!�B��w�05)2 ̢�����Ň�!a~�D2:K���-��=%�����z��"̻�H@�i!{$G�uQ�R<��t�Z�p��ĝ���{���^�@<���|΢EN%�����5:�����@{9�f�5	���=�!N~\q��?ϢՅ�w�o�Dk٫(�31����A�����i���Y��\Gγ�L���XSXd�>�*�� ��ʐ��ކ�lA,���7rF�&�k������A��%�ϧ�ֿ��=�߃��o؞��l�B^w���e�#��o���s��۷�*qr:D(i�p��;7op�.���}�>��Ul��@���0F�X��g��`�Z@`���՜2a4�E��"lJ�rJ0E�o�!TIo�t�$�!J�9)�Q��d?�]  f�?<'K��X�eH��1�g���wO�W��E�e�R~T��|��Pv�
w��A�S����JD��Sڬ6�E�%�O 
@�/&����cr�>�$?u����3������}<u��d����`[%d��#�V�.�>3���0x�jn������;���AARo"��ZNyY���n��(�'���W��Ż�4v��y׻�����t�>�м�t��B;�]�/ܯ�t�-��ƫi�J�Y�7�杢L������l���hV�#������XH���i��/>k@�9A:!��Yi�L�C�����a.����7<���3�t�<��a	��iѺE	�[���O ��CIqi}؉K7b��NVv���^�L�.q2��� w���x�{JjN��{�d����C���	@Q��Ypa��Ԙo�U]w1�̗	�T�?7��q2���Ib�H��6=u��\Nk�)�U mװi<d�ح��>��FGK�%&QV$��Y�$���24�o���׬�����1��g�Н"�Oe�=���k<�}�P�~� ���
�(k�5���z��$��6��-���eB�s�wOR������� ��Uq\,��)�πq<sY��'��v�ϻt%�%,���ܻ������W5��7�&�.�#���Z�����4Q�g@ ��t$�xc�y�޽'�Rg�}qߝ����B���"`P�}r��v��9��.v[c���1�u�x1+ЈC*�Qw�4�x�RÑ��I��ܶ5���t�h����*<|\���]nB!��D.Oٳ��w#lk����*����c����c��r��Z ^��٥r�L`��<'O�lV�%��Zټ5���曑�kǲI

C�[�E��O��Em�@��K���˂���(I��'[7�Ԙt��;2���T%��<{i��@H���Q�?۞T��� �>c��iN�$�<��cp>���Tu�����J�`~#<V�a�Mf���Ȃv�L#1}\G�Ό��� �0��I���"�cg����JT�ĎփN������T�$2b�8V��������iŁ.!�6�n��W����8	y7,������:B5���q���s;�k��J�tQ\�UЩi١�`�7�[m(�lAPy���"��߫Q�j�	�೩}�Xe��	^��
i��`{�-���]��2p�M[}Hv�n�����}��a�U��M�*!�}(ZY�*� ��7���E`c9���n�����G����Yf8Ժ1��%����	�;}�9dW��K��0l[��(�p��_��Pvb�*�ޖf��v���l�j���i��C#>D�����Y'�kK���6�؆��"����yGɌiz{5�Ao�5e%ើ#ѣ/͆�.�ⁿ����l,�ĭ	�Nk�����?�f���xx�au۲�8�u��B:�#Q�'�ӝ,���]zPQ�cC&`,c�L֢�k�T�����TD���!����O2�B��k�&��H�:��@����⸘�����JN�u��uf���;p��D�}��e�_��:�s�^�!�`�s���|r�|�-����7G -�|��dr��i�P�����i��r�(gӓe���_�򒴞��˶6���Xu��Uc��=��!����}=�I�F��{!�����ѩ�(�Ty^�EY�ݳ�����ߚ0�YH_���ߕ�X0���x(8MNT4Ǒ��W�M~���ꡋ8���av42�]�tE�ź`)v�J5��EB���c�`���^����.�t�:$�gX��Ч��D��v���~5��z��@ի�sܟ>}�2��[1S	^�v�uV�:Ǵ�@>�f��p�K5(E��os	/��y�/�`�'����M�[�� �j9��E��iC���x��tjHO��MQ�D�B����\ċ��3D��]g�8m�[D(;+���B���� �Ӷ��>���5�.��*Wz'FII���������e��3ma�<� ���h�e���rŗ4����^�3"�3�o�SL��(�4#��i��L�W)�}Ǡb�
�kL���x��k,?��R<�~�C���M��u��Ua�)�
� `��i��E��ue*�7���H{�:a�Ȏ�s=lIx����������CX�h 3*�4�]c��M�S��
�8�a��_T��V��A���[��b���Ddb�rjk@���jh@':fHJ)�ڱl1�vG��[�\�dԡ�;���ؖq���#��+KU@ *ͬ;n���H�Y��h��@��w��c����D���[b����������X�H�w-�H�/��&�g�$�J6�S��bUy���䉉L�!��t�����Z�4�{+�de7�vvRJ¡�̋,51�(�R���SH��u��ғ6wx!�GZ`y�Eh��/)��#�L��myc ��Y�L�l~�3�!���J-ƭ��nf���DU��8I����Z��.>Й:�2��b=��UA��Ƽm ��޲!�"����_yf*_�i���ѷ�5Ev�/-��ם�gP�}��3䥢��[���}��);D8��b���*W��=��~S�<�[X��U��=þ��k7RVXB��_�W}H�~H��<��Ψ��Zϝr�fV�%�HrR�w'Xd�ܽ�ϵl�U	M���fB�q`F�q/5�����FP	�K�5?w=w1w(j��� g2 �uo�8S�&c�M�xZG��!�y�L�-��#e-�g��1{t���I>DKGɒd��j17�1���˦����VzG���#� ��G���|��*Q�3d,�VH�^J�u�t���\�I�D�P !rܢ@��p�.=���˟��:|�n7�כ��)K ���M�U�B�2�g{��h�Z�1DvU<uY!!3�����=��	xq�qp�=p��])��+d����C/��qPx�>��(_f�s��2��uA�T�z`+�L��v
��;��Y*��.W��Aj���S���; ���������i^ߺ�-����c����x�%&ㅽV��k:7j�7�@rE�s噱2R�fqm:u{\h��a-�-4�g�����8�yW퐱P:� ���E��d�h����
�n�Ϳe��K�N��P�٘�p� ����1�e2���wNj,�Z��A[!~b�����ݕ\�I�\�&��8㙟Uk
J6�� ��+�!"�K�_���3/��y����:��EK�y�B�H�������և�B���q�������0Q�g�An��4j���i�� S��ƾ7s�,��9Q��|͑O��i)]�+��:�u?�G�,3�K�r�Lz�v�����~3f��]oշԹ���8d���B&ǦM��yÿ���F�e�źM,�0SC6�C?M�J.9�y�S���m����K�|?은(��f�9��[�1��P$i���a��^��l����:j�/��݅"��]hC0`�.������-�"p�l�ӕM�d!�Mkk\y+�����u��%���� s����J�B�=	1zbp�܏�::V��5ݵj��G/w�(�6�mPϦ�7|���*�&a�L�o�(�#��.�1`
k�ӛ<���Gt��48n^����4PB[����9��|��A�
~�M��L6"u{k�;R��N��oH�R�����ZC,��j~�
2�]c�7�\��3��d)ǒ��3B��j��!c7/�z�.���TXy֞�� ��{W�k�pke�bm�Q( :m�RmT{���%��`��2�C])DL6�i鮾�S�k�l4@���f7�-1``7�8�Y�X>'��Ї�9�P��;�����@�uh��_CV@8�x�@�J:�:(��I�sb�H1�i��~
| %)�qG��f?��0���r�z<93����'q�n��_1� L��$?��C

Z���M�P�-�!>{�<��$��zhGȧOy��kh�V_�_���,0�3���{��,2	\3��/����з�j3�#��`��<5c�w�%�Z�����u�9�9u�����N0SM��L����"��
��J��61+��㨧��^���+u�A�.�H�w��&=��ĳ�t�W��Y>3��N%�j�4��絑��BH�I���3Ph��/~ ��Ư���[G*6@HX������+#�@��fN�iΉ��?�1�2��3�,��/2��k:T���f������˧�ЭԲ~8�
����=�H@tza�$1�("0rq8i�� B0��A.Y���e� :�9e(�4{c0��/�5T�kx^�:�x�n5a-��N���:�r�a����� '����FR12�S�=1:4'i4�K�����X���룠��!�l��Z��Xb:��_n�A^�����d,����7 ?�<����h)dT���d�O��` �]ݍK� ��샥%xeWh�`x����)a�"��ĺ���H��Z�x���A_eW���_ӏ�0X���X����s�d�;������	�H�᛿"bh�f�NO9���1��
�~<c�W�]���S*;���D��G�B��NH2���üe�k�琝X�1���+��@��Λ�Bl@L6�Su�8-8笚�Ax��]�<4k��?���C� �[�>4WCuzÛ,�g�u���� ��xX���-+N[4$��[h��io����#0�ۧws�*�A<<��`��eM˕���TL=uᣚ%��"駱I��D���9��Aue���B�9�.6'�PZ�Y/���] ?G@��]�e2���{���mٗ����R��
� 	L��S��U��i�<�Y��X�IC�d�LL�K\��g�d����L����A�K�H�Y{)�l���ec[�����{]��fY��z�S뺟��{�Ug�,��~}���_�G�����q�ޕ�u��)|�]BN*��b�����wl�Q'n�ȩ�R`��(����6#��t����ZW�,����S�?��0�
zk�28|�/)�㉓4�4HGޙ��;�Dq�anV�� W��Ӓ��L�ua����9�+%ڒAQk�z��&9v8�O���,�x3r��v��o3�9�T|�^2"�e�P#�C!��� P��3�.��f��b��3U|�!vh�a�k����F�7��R2�����>
�Nt n�5+�b��k1<,<m��X�1�ry�H\�\����FA;��5K�,�����t��i-?�P��Jxv$�j����v�o	j5�M8��K�Y4��5 e�R��j���="0����e8���':o�E���xd,l����W}pC������\�?p[���g��8�f�f��M�>$��+UD~Y�fkUr���i��'Sp��
��T;�,s"l�<��8�Ф�h9M0�VZe�l��T�/�v��j�^���ƣ�~>]n�L�0e�M�gpb���*�q�5�QsRmy�
�_�(�}���������8e��3Ч@7dE[����	^��Q~�3�=X_d1ta�UFmd]���.fCHg�rf�;y�E�`�h]��V2/ڊ����"����^����Zm9�M�ՠH���΢$i����e�9&r�=�fn�T���$�t���]T������3G"�V+�67����m�$�M�� �9p{m�d��Y��.ԷI�T$t\`T���}v�gͨx�HV�s�QY�[5)� ٝ���5�T�b���~�rZSL��з�ҫ�_��W}�vIO597Jjr�c^x���Yʟ�F!�q���3y���.������o}P!�gG��p	
PS�����ڈy C-x_b�\��ZD�xtsJ�@�X`ӫ2�/�НFr��B'���x�s$�e��x��B+�*�֯�'��3ׂi�K[�[��w�cO��'P�͊����H%��#'h"!	�GD���g��v,3i�t��2Y�����#�����=�L���f���b�m��o3ޭх0����I����Ч�ޟ���疤7�p-���HD����Y��j��M][?��1Dk�s���#3 �v���vJ� Ai6e@����[:]�芜/�0��*Mi]�	�H�nq6�1�	/�M8�n�8C��m�,���/�r�B�����Zd/���P��M�F�Vq$UБ/0�>���:�j���ߜ\|�%՝��{�N;�BAO����w��WP�~�R.��o p*7�݆��h�"lg墡e�붛�+�,�Ιh:ot��� ����Z�/�d��sy4��C��;zavU�R�����NV���hG�R�%���$���*�:M�ldR�|y�J�䘖�-�LhL��|�32c�z~����p��e-�{�jE�N{�Jgw��~^Hh�l��ھy�0lJ_�|���n ��H����ȭi�w�",�Y���JE���2ȋD�y�7��]��֬� ��6B8���(�U��Z�ju����L�y͍�:��ٹrV����I$ݢK^���4�#�o2䁷�Z�}�/`��15d���ko�)Kܳ���S�£%�[�v� ^����e/#c�C�@p�툫"���{�Uu��\�g�no��ET�o�H<����O���������km;%��C7;�ʴ��U؅0Jƹ3
�$0�{R�|z��k�ځUw.xjh�פ��A�O�Hm�84	dkۮ�U+<��||�AV��Sw�� �g�^8,m]��a���[��@�	e���K�a��;��5����qU=ݐ�ܯ)����k�#��$2�Β/-�@ A)p����h)��N?�/�����g��(�	�a���t�뼻>QJ�C�GsG"�'�p�&��,ΖV���;�u�ۏ�,c�/���lL(a��IR��N�.
�:9�[���F��C����y8��zDjį�X�X2�.�"��&,���ޅPl���b��L�6�-�Ͽ}��0'��Η�5t~�uLsX�M��
7�.x����������	��	�z?�����8�`7�2���薻{%���/^�5��qNe��ꉧf�
8i�!��xy�U�O#P�ѧ�S�2\W�2  f�8���H��eS:c7XL�5s�Y�v�9҂^�=jl��=I9\s�-i��M��=h;i"Fb�~�?C�`�I,}�3��?=ۄ��v���(�I��yI}�K(�1^pB��w�_B)�2@�Űy�\T�@�K�P!H��
�������닊��0n�.�F٠�'�{�֔UL^����.����ty�Y�DD��.��K�ꯧ����N�D�s�U$��
/��0i֤�D�Ef�����	�jk���T�-&6�,����R��6[20G"Gk�+���W[>	��3�~o!t&7/h�?�b}>Q6-QG	�V����:�_�c-r�s"�\��VU�6!z	���h���=+�~Nd�B�h����Z�h� ����mYP�Kx�bC��!pG�KM�ߏ�[ ��}9�ml���2��0GH�����^��kju��G~�dB^�DZ��,!�
�]��|�Ț�������$�gmվ+0(V��`�T]��k�m��72Z���Ӳ����^���E	�}����^�P�7�U{	��� X@}���\9�Ԗ .}�LMµٱ�2�}�CWlAW ڽ�`�@C�t��qlO[nXɿ�<+- �KX�y�H��{���f!��f/hֱO6��BA�]�3~Fz ��S��*�b�I��8��j۫͐�g�}�+�rk�w}�pJ� ���:A���h�b*�o�.,�OA���V�z$�Yա��p��ಝ�57��'�������?�������3�ؙ���c�i�Cpҳ	��^��;ma��j0|��pq���80����Hl2F�TL|�7��|�%��a�J���zv	��+�"��HW���Gb�U���B*�@4o�`~�=��焇�@δf�"\"��:Š��ȶC*-)�����!n`�u)t6��m^������2Ԇ��[9u{l�[�٦�����O�b���d�+ϩ �
I"��o;D0K���hj��	���8�U��uB:#�"kz��u�ѡn�� ��'S獐LQ�F�x��,	��-~|�9K`-�L�|�鍾WE]��苴�rH ��_E��$V�p��y�Y$.��Br�l��3��������.�jV�6n���=�U��D#e��T��3���*�-����t{O�r-U�$���r0K5фP�窔W�<Ͼ���Ou�F#�jַ�LQ6.��g�㙎$�4=>�i�Q7$3�/��þ��I�@K��b�p���@�|��޾�,=Yz(���*v�Bye4�4A��y�mC����w�C�6NiU�����#�����Z+O�w�I�xd�B�)�K��r�V&��d�ˣU��6��c� �l���p��Up�86sN�;�?Qr�0�9�48d�.����f��f�������E�p�#����|輗ǚ�buLK�a��'Cك��A��yt���{�����C�'�Юܙ�����F=�ظ+?�z� ��SeQ�1�irj���	��w-�yQW	P�¸����"ɿ��L��MCO����d����UT�.PP��!sYL���cg�#��`9*��y��̶��_R�ÃɋRo+���F�ʅ E6g��[iN��������T����j�n��&y��?\�s��	ֶ�����y�lx�49Kkɬߵ�O:W����r���1�[�L��tMj�3v���$#�0_�����`m=��MSG�7�WB�[�~���Y��7�*��>:pMmU�z~ָ��33��aӣ�8SD�Գ�:F*��餣����g�`��2�r�g|5���2�ji�A����<����,��\�#Ħ_q*[Clo��<����W^bˈ�N���7�ů~�����S@�<�y��������(�^�[�o��D��R��(�|�W��\�@�*36���m@�]k��_��~5?�=�A=:,"oMd��Enp���/�7�3#�J!�����UW㌠�Ƴ�*MSsI�ǂ���j7&��kd�m�B^�?UI�AHe�$s��Nt�f�%&3��O~��O%L������v�)��7T8��`自o"�`��wr��>�����!�����M�	+E�����r�
���5�x: 
�U�:��gN�Q�:����x �<&$B^�U'�� -�����[���4�*�qy��yJJT�M6Aq��X����1�˸&��o����R����8��JQ�B��h/Xo0B�@fb�a�����%^���0��ekP�뉨K!E�����@�a��߳"�0�u�z�v|��"g��Ш���%�3Yp��I5�1b�vK%/�[QF8<�`S��ơ����]�`K*�v�z�q�K�5w ���L�iPY�se�wU���^�v5ͼ=��NNH3ᣛp!����'���E����o��a	��A�.'�B�J��k;N�b�d�Ij�/R/�s-��+�M
5 �m4�B��ur��v@�!��6]�!v�2ˌ/w���{KяlZ"4���v��n��cm k�����\TQa"zK.��k�7���}iq���׳
"Q�,A�\���+.B��,���V:�SL�2�H:<�z�e��eG�,�����`
��������T	|��]�b\�~�@$Gu�?��T�{���5m��C���(S,�4v�t�tyWZ�����EK�����Z2cH�	��<��<(#2�r=U��<�e�H΋i�h���	�{9D57+-9{ӏҺw��QMʎ�M�����H[�n��B%���S�ϜX�;I�@����u'�/w�����&�o�Yي�㹽"�����#�>�=)�2��݀����PW���͊�)�����U�/��6��+�{�4���3ld;<�G"�_��^��87uv�!�I��q�H�'��0P����,�� e�Y1�`���ߚts�)���!rN�ll�����'��H�*�݈"�(B�ٷ4+4�0���%gF{���սx3�b	�.f�(���î :�]�>j'�����^��r@�Ec��-��j��C���?��2�DI@xoJ�Z��=�7��� D���{�(O$����`h�W���z��Y�
1�Y:�/XZ��/�τ����xH
����*�BM�����	�»:[�X�bwE��5��fƫ�t�6w ��]��>�h���ET�����^��]״x�V��#�p(ٔ���TB�ϡI&l�J��$���^��}�� ��+�������f��-�x�\����/����2CɢC7��G�R6��-�%(Ƙ�mO�;l[��]f�s�KY]@��};���1A5U������o�Ξ�n�����;��}���2�����ƕSq(�]&��#g��|��� ��-�w��V�N=�	Q��[�Ro�K�*�vBW`u@6D��I;�b�4�9�[�Uz�7&<�>�c���!,(�.u�f״�$��7�R�␺qfb��	K$u���n(��
�`��Q���-�&��ݦ'����5�Z!��-�;��H�k�}� 1��.i�|<���v�M�h�A�Z��_3�5/�UZp��Q׋J�l7p�u��������x	U���a�CT5��*�r��0e�<ޞ�g���J�Z����;�\אBf���C����~!�/���=�w��P�RD;�����>nC�CĔ*��܅~�a��f�����u���8���İ|u5�C��;���0b�
��2�� դ��hu�5�>[�w#��U�d����G�ׁs��#w����Ra�w�cc�,c!X�ƪ��}�c$fR���"��
]��p���`5ԗ��N�n��kBOcE����x�e����A��H���Ǝ��WnZ���!���Z4<Qf����׉� �}	����R������ɐM���?�ͤ����1�C5���J!�_X���5����:y�6�@ܓKz@���0ł$O�@��ڶdu���c���¦H@�yx�U��Q��F�B�t}�l(�>�7�f6�bL!xW��Ha��I\�4včVP�C��lsW���
_J]�UgQ����<�*���k�~L��V=+Va�e��!�.$f�̖���nR���� �MCOkim~��Nl�PcΑMM}vX�%!h퐐���L���F�*���uN8渝A�&�A㫊cb�� �ˉ���,ˣw-��0�=���e������`1�5^ó(����;q$��	����E���ԁ���M^����<�ź�0��vq#�z��*�b��f��iiL�����SU6d���Bm��^M�Y���)7�!c��lT��.����z�C��c׋s8T��K�rR9d�k��&�y�$����YDr+���gVa�i�U�8�{�Rt���h�,RS�,�~�d=;�ܯ���̌�Q�dCvϞ����
=���N9��uݫ
^ΟnҮ>]��T%h��	�=�h�./�ū�1���N�oOUH��5$ ���U�|����\�!�&l[�F�24)A5��+>�ˇ��BڒN}��d\�7�2z��N�[P�2Ȕjq"�1�i�J�[:>��\s#� �3�x��1��^U�>9.x��+YncA;m�$���;΁�wߍ[�;�E%���f�?�A.��<�M�OA�� Qo@X$/�z���;'��L\��6��K^NlE��Ƒ���-�u�fF�%;��PSҿg����e}A��2����@�ѹ�z�������w��r�o(k���,��\w,բ��n?����>���@�7j��͒���Q�N�'᪮�>��цV�
�;���+�2�0�Li��g��j�hf�s�Q�%� ?�cs�W.�!�K���Y+�"�!��T�U<xO�x�/X�cw��+�v�Y��.��^����J#�b��8�Ȭe8�j��!��#k�u��'�U���?���5���'3����&� ��-_���f��f�g�R>im��\̔�B*�19��]-Df)Z����v�ܟ�G2Έ��^�loe4Z$�"�)g_j{Z����Y���bkQ�A�%����y5���زêԡ]�D�X��u���H#�#��#�4�b�8�
��8��
1.�`�"$ ��
RB�Z9�=?�V׀#_Tv�$<bLb�!ګ�/wQ�T��?��"9���Q.����K<5��U�~��댱�B4X#�[p�5RJ!���������>��wl~{��vDLfØ��2��B�2��ƅ;�l����3��W��*�v%��ReK�k�\m�$R����[}�f*��V���fS!�,�n�vlp(�[���hOM�t8"YTp�9Κ=dqs�r��[颓�y���DԶ�E�5�kK�^	��E�P�9���~��P��>�� �Jېd��(��oϊ�����A�d���+#"SU����|�ƃP�w�P캆8(nK��/�u�^�?m� 1��\��y�*1խ�"��t�2B�8��k�myn<�ݚ�g�O?5�v�/�Φq�xӼ/`��ʵߴ�
��ޤ��56������̯Ό��㪪g�˽��8r+�=��Kţ^<Xad�`
|7��B@�cf����'�^�!�P�@�[��B���_D4�ԢP�h�b�Tw�܋��`ܣ$�� ��ύzHhwx�ҐI\|(�H2��VeC���g�_r���zY��,	"a�����@&�=��s�2tHy,���D��Ԇ�Y�Sf���i�C��v���Rm~{�����IG�m��d�{�bs����:�Y!����6���L2)F1���r�[�^�,�����
[�P��B�������YX�B��č��U�0<��Kx\�o�*���~��" ���2>�I�iP��>����K�|O���`�,X��l(--nz��X���v�
����B\zvq�j���1 �y�Y"�z:��y%�`$h�P���e0�DtYT���x6�ֵ�����H��+�����@�連��9__ԧ=8�r�?�,p�ܠX�%���2>t�`�!��X9��X�K��M(-��z�
�u���4@�$Ð�6xvB���rs�W݁��C�/M�4����f*��w�>#��<R�&DE�UL��������c�9��͗M�%�-k��#$>� n/��n�}}�Ct~�O��3�+�6�%^��L�T��=��+?���eg�V�:�� 'NO���]�{��݌��m���a��;��� ��s�Vg��g.��ڏ�]O/�u@r|�5����,��ͻ�6����h�|	س��Y���l�֔Ϡ�[����9�U�A��n��VHT���##_���ѓ!&V��O�=o�m���6�[PDYu�e�k��wX-`$蕿��V}�H@1�d���� |�O�!��BR�/Heǽ�Ev��,8ܰ��~Ϫ�z��>�e7.���\��e	�zmu� ��˄P�q'8�����?,�	�����,(��,��u.�c��0��^�|k�V4��4q�A�g-�ќ�.ٜ����l���H�t��R���MWC�����1�l�Eˑ C�̫rf6~�_�a�g5�T&�X$z���D�u^��B���1������G��U�i�ѓZ�� 	�ț3>�H�}N��oFn�Z?�� Ǘ���D�I
��i�t�A5�t��}�tݰ��xC��"��%;�˫(�+���?��2�ø�K9���ߴ� q��q���)�L���rA�j/�������8SV����FA�v uP�c�bV�e��s���EKE��f��*?!5&Y�HQ[2���(YC2����@E��p���o�q��f_�^�ǧ���ii9���.e�荸�1+��\x��m��As��.ʅÔ#�.�5C=���DUn;:�.B�Z�{�G o��с1sF�Zˠ.)��ܳ*<�'-"n	�L�0��a��6E۫��)W^i��GM���w_�|�OM����T��c�A����CD�"/�����YÞQ%��
�a��<��w�t�p�����y軯�ݣ.��M�l4��ˍt]��gx|����
�8P�c�<��Q�M�>�W�=�Yv7���p����;�JIm$�.;9kM�� n�_�����7�%����gr$��#�'(�)�5�
|"w?�O�3����T��:�Da�N�������I3��1�u��rB������:�N�H���N�*ϋX���$���9DG+�9�u����CHnAe��g}F"l~NdS�K�u�n��h��Uj� >��9,�@E�q���-�aѭf���9��ּB),7���\��?G�"��Ҹ����t�-�
Ʀ�b]Π�hR���o�>��	�Jm;�uw6��ъgh��b�`��_�:��(�|������`��D+�'��Է���~b�;��ct�-\{6m#�G���L
PIįf`��g��zj��u}[�Ѯ�-���}����d���!=C~��E�z���ȞD���A��[4b~�%��C�8O8�O	�Ŗ�rUH��V��'���c������xC�X�pc�=����T��<0��`b&��\����so�	aiY܁6�$4��*��$��|�Z��
T3^�7�m�5�q`��/x�l��h�y��3�96aix�n��;Bd�`��4�ϸ�W���D��:a�Z�l[WZ�DHT��̅��X�_8j�(�������1���\��頱��s�J6�׊����ʂ�5�-��n�'K�A0���h�JZ�vL��/���F��q�"��W$���{U�LC��R퐰�����/7{LI1/��T H�l�]��-��_�gF�6���D��J��.*zj���d��ڠ��<��H�P�*-�^N|��N���~��2�X�������aF��&I�3pz9c���|@|�_
�Ġ<�Ϭ:9d�߆��z�ݣ���'Y
��uD��0p�2}��V�e��J2�1�� j#�؋�f�FF$O&&�&�;y�cu�*�Bу�,��Zq��镄�2@}e
7j�Rj��-�s��;,����b�Ơ�`������8gX����[�u���jE���E���Ӫ綀(��f:�e�+(F��ݱ�k؀�I+>��j�0�XCj!Hˤ�3X�pQԻ�~�Ͱ�j��#������g��܄}��sX�F�q��V(�k�Dk�=,����r�z.c~�I�����P��/D�쇐���N�Q+�;��(B�N�%���$I"���%_��2��~�v�_{���I##��@��f�~ڧ!���O���t��r�lL5C�7�'�
��s��SV���[4����A"4���${@|��;aڶ��j�
ߦ���� .{��ZC������ۅ�z#��,[�u���G!���R ���-�U|64~�$��� �o:�/.`���XIɰ���SZ*~�1z8���$��nĐ�HRdr9X�K�֋�-ε�|��B\�m����(�D�����0���5r���h���i��wr�+{B�B�ܧ����~<e$����J��a�q|��H}K�H�y�����ʻ?�h��=x�T8��AH�%�P���Ҫ�s10a�.���2wܖ�nA��@��@K5��l���CI��#&O�����*�7i�^��}�8�G��1�A�[�����׫���V�7r.7�_a/�겆oc���46:�%�P�C�w� ƚ£yoT���2:�����9�T�c��*J�i�,ozL��� D�V���k?;^��j~߂&d��Uka�3�"�n���r��1� Cj��	���C-$�㞮u��iFoX�y �O�!���u��%	��&�`��em웞�h �Vo���d%�#�m���%M��I����f��/�|+�?�4�=ͥ�M`�QPɐ��ſ��{�9���ssDv��r�׆!�ƌu�Wѣ�Hh�� v֫�['�F�q�_L�e[v4�-�R����pE|��a�����*�����V����K4����Cq~�c��l�B5�QV�l�Q8
=Hb����ůk^`{�C�d�ݥ-D>���5N�'!�mU/��#�;�5��7�U��
;:Fұ�C��nC���{��W 2����n�7Qhw*�1Fw�c(�=<��\��4$���2gQ�ؗ�j�$殯.�� Bg��ȭ�w�ғU+\����Y��[ �l��	�	���U^ҩ�h��eY-�7	�lmxg���9���g\+ȫ�?OJA�6�e���b�~T���Lv� �y�+ L!�x:~�r������*7 ��8�SB����Mm���ƍί*�d>Ĉ�][��Neu%],R�k���o��ƣ~���i���z�%Յ����*��19�iw�\��V=c����4Ѧ@�����j����Aޞ�jd��KqjOl1v��4�Z&"��!�-���j��f�4�Ҿ#����i6��i�3i�X�ڌ�;5�1��ͽ3xʅcҙr���rR�9��-c����v�jd�*(�T���j<���mA�]�̱R�1��O��.�<�����OD%�7�ej�5��d��U�I�R��t���=xo�����y�A|��o����ȬS�M�I�#��h�~�{�p�?��4��m>j�(<jNn����R��&����g��B����F����/��E������٥꣔�#�dw�C(��C���; �_�����jS.��!���O$?&Qؾ�ݣ��h�]��ޗ�s��s��9xA��8��5.y��;MO��e��C�/��･s�P5��9��H$�UӀ�+u�c�iu����������wi���Q=n��C|^�5A�ފ���L�_b�)E�s��#��1���h D��p�W
��/RN�d��:Y�Q����lCe�6�� ��:j�E}��!p�������8�(=�Lт��IB�V��n��=z�f{�yC%� �M	S�A�%d���NN��=�ca��rm$��<��%���,�b���̣Kika��/�+.V#�"��
��v���;���}�p+3�/���&��л-rP�Őa�s*^��a:V�lG&�{j7�(�փ��X��r�׭�=�R��f3�[�J(���ӂe�5MP8&�KE�"6�ذТ��{*�3�d�󓶏B�ٱ�ﯝ���F��!���ow���0[Pl�0���_��oس`���WQ�.@���3bmW�����_������^�!�)_�!�~��\7�,;>�7�Ӎ[�s�^q�����-%��N�8��>��o	"f�⊎�J�B\A�J��\�9$!o`��e�>c��[@H,�b�����8&�דl���uw0-�Ӎ� L���.T������0�8��.���\KNZ��}8� �:M��vڢE�)�U+��1��5��f"�Ã��}1��S$5�s�߉֊83��7.,��񦻖��MJ��c�cO�*㜧�S�J��*�`:��^����j��U<��0}w��>]�$���<�^�5"gW� B���_�rf5Z�
 y0�������4I���,�(4J�i!b��w���"g�>T߭W.��QR�}q��*%������`���^"���j���|?
#��-���y~聜��_>O�>�'F�Xt�������k&�b���TV��+�7�<Ƕ���	��#,d�d�
]��S��M��[����o�x�]4vMS:��?�\h�Y�Υ����+<�k#׉���o<��Jo�C<�ѧC2�&�%[�6'�44��m�6�L�K��������Ȫd	<����1���_
L=��&V^
פ�j�3���Ox-���Ţ�I�X`�mN�U���V37����>�?�76#-���i�@��nf?8�3Ϳ�oY�o�S|v�6��C׎�p�9�\������K�����!y����:��C�[_<g�R����~�w�6������Lm�Q�>r�0�t/V�\�J�ǀ���^�ֽ�>;��06����X:f���J],;�k��c-�wC<t{2"u�;W}$�?�_嗀�S���ȳ`�6�����4+�����	ɶu���dt��u���s�u�ym���==�ˡ�:��H����y�K�F�u�:��r�f�MR��JŬ]J�G�Od�'e��ˣ�i�//�~ ��h�@�)�{�HZt�b  �A�׳��)�u�s+Z�j��B�og���+�y�b�>'p�
q�X�A�9�b�"��jNQ)�
�=n_�C������,U ��*1�M��wC�����1��s�REH]2��
�W��fn`@��^���rq�J��6��W��T�e��]��mQo��*��H�����t�@Y#</U��m6K��̊|t��ao�m�@�r +[�61�ȦL��.�?�\�c���f7�_kVqs��3A�}$óO�o*�9�������c�M���������X��O�K�#�Ԍ�1M8MV x���\�u:�H1��K�5�#4�l��ѕ}���
����:�^z���OOeL��˶C�wDc+$t��]��}AOY�t��(�]�⏋�HLYj�S���$�yU�/�l���G�N��ʜa����� s ȏ��ڝ2�y&��/��o���� �Ӱ�L���]��s_��;��.�[�Gߥ�{�=�P�e����ᨓ��C��a��f�>��V���Ķ��s���Rv��:a��.��3��@d��)�Pѧ�ʇ���*}�-#�~��MFq�10HS;Z7QT\�R���$.�	�B��pР�����ӊpZ ��e�i��O��5�{��G�P]���52���t#�ؽ�����vP�I�� �����s|8�׻杊\c"5���g��j��p	�B;�{�8X�a����e,Ó�Z� 27�<�:�~TV�;w�/?,�/�
�����F�=����\�@ ~�_���Feۨ)H��ު���a[�����s�>_�F�������*Q�=��.�0�g~>F�[���w��`ס��*���<ⓤ���q��Xxq� �Ѣ������ި��04p�.4oq���n�ǜl%���.X��{ţ�;ۅL	�D���w��t?Lq��=���b8}�Hd�ڧ�U>#φX	��!4��;$���Z&��Vj-$Q���K��o��m���B����vd�=�\���jf0Fa���*�f���0�
ZQR9��<���C[:P���b^c���9�ێ�y�3�ǮRÞǻ�
j��C@�J�j�D�d5��
�(p�x��H�s�����\׵�[���Y(7	���+o↸��=Lʒ�|�"V8\�6⋿�]M�=�p#�7z��ܸ�x����#x�u�EK;���|��4��� $?t� ��^D��n�.�ܽET�����]ꄯ���@>�nW�[MΝКB�1�r%�"ee��_�JP_��i����������%��]+dx�~�@k���[�U±=��n���vڮl�Nu5��,Ro�K�$ߺ,��s �fM��5Ȁ[R^c����!\7��:G�%6�mu�)�����@��i2��NMR��:�}V
�������H��:3���G�=�KK�0Ö�GP�	���ͮ��F���S�5 4C���KЙ�D���1�u�h��U���ݠ�$�6`5z)�I$3�N3��ġg��n�[u����b��l���s|P�����~���ӊ� DvW\��T��te��/R��� ��Xr�t?Ex���8M:�����%1�l�>{t/<ٶ�L�����õ&�l-�?Ԧ�G�淰�`T�v�9�^[�����H���3d�������5k�n%�.4���t (�r�4���
^�DTZ1��<�?6ۅ7��QH^[���%�q���C�e����oX7qo9d��C��w��͏Y<�H���2�F@��*3Zf��Ay[����#��Fj+�$}��ғ�`/�r��#z����a�X
��a��J��eL<����ei���?zZ#u����e��Mv��Q#qB#"�QIv}��#�p*쉿coql���A��v|G�#.OpVA��QL�u������^�_�X��l�)狏1��pv�-���|Z��\��{i�޸$����c�m�v���K٧�AV�*�t�_�-�����ڻ�����$=�{�Mj�U�~A���V�H�^.u/j�cK�_-ZVl�%��a�v �!3�j��۫���A�Iپ�
;������������	�1�k�9hLԇV����;�`���JQ>{۶y��<%k���	M�)�H�����3���$=|t�"�[	�/j�\=ʩ�Vy�+ �h���o�KO|���w���𬺨�߂�S�p[:�5����*�k��i�uK�7#p-v�cY��J��v���7��w�Sn�
҄�g�\�_�v__q�k�$�Se�4�*�#Цa���m�D�����u��N3�qN!������)�b��c�w�eu�)}x�������ݜ-�Jm|{��x����,��Ԕ��q��\��ш���7N�TѽT�����D��a���"���d�=TΙ��S^��q�(F����!_�%���G��0CW��ӌA���#�~lK�Ř�i���)��h_��.s�b�Ř�7�mη�QyC�M�I��&7�t�Yurx&��f-*�1u�Ne��8WB@|C7�O�?��G=B�{���S@�k5�W�1UF͹t��Ӧ���9��#�#����}^�Nnx#�L��g	4�:��+��B��jʆ�b��K��q���T�`i��r�����&��8@fY�l�W���VG�;���������^���{���*�נʒ��2���8�=MY��u�7Y�0~Lh;�:r1yk�9�n�v�#�����#F۲b=0o>������0��%�,1G��u��x`��׻��Nj�> �A��X��Б�y=	Q�7�� �`(�;�e���)��l����B;LgⓁ��1k(�Bf%^*��\K;.�}T��V�w� zk@qFۨ�Ng���S"�"�~�n�Y�ϲ�����������cf5��"{=Iy��F�Sb@j��u5W�-�$�_��Ĺ����� ��;�D$��pX�4���,6Wq������^��%pKczN�C(�1����	����J�F��h8u����c��O��h�!�-���v6Ut���(�$̌v$��$��Z��!��M�
���n+��$o�0םpӕ4Y��uY�֥�52����I���Un󉣘d����>z��G���Nc�(��M��OI�����&���o��g�6�C:�u	�D]�L�R��T#��m��	V����������YL��ܮ���ї	�$�!��]���0X�rZNn4��	��47
l���=���tޜ��i�N��K[��n���,���#s�u�+��v��r�Ԡ����ʣ���1f%\�۝�{b,���?� �֡�����e�bWQ��&0�Wl�޹�S?$�Q��kD��esK"��:d\��g���.�m2�0����DԪۨa�fľ��6���:)`�
NT�"�O���|�̛�>}F� 
cJu�s��+���������o�����_�xu�z�r���u�=-��$�5:"��������B���� �d�`��*��a��Y�n�X�T����(�Mk����٬ �J�r[�A��� ����뉆�& |]H$Fxj�>��i�]��v�,KEf�s�c�\�ԕn����gjb��>ۊ��0�H��Q�I��\�n����L�����8�<��ߩ[����=�er~�F�m[m�j}~��������ExДm�A@sΤ�bXCfb-�M�y-U�|ED"��7��Y[���*����,׿�C�?g��L�ZRxJ��+�p��B�O���V���{H�7+��K$t�.�� !ݪ�6_|��hw}���<��^{�_��sB	�#]^���v\h��MЄ��4�U<���>���2a�G.�)��M���X;�6�u��g��sI�d�1��,�����T����h�Y��mB���
r�?3���G�x�͋(�}���T�A8(��pE���Ġ�f��[�8�Qo��iUN�I���t�f�L���0���ms<�e;�U�E��k^�����S�k(:�W�~�$*�H����/�ɝ�Y�S�� kY�P̖|�L9��*qJ�J����~�"�1�&��X�Ի�u�V�L�e�S%����!�PC��8�vy��kGkK�Svj��lv�f	x�m"ɸ�<\x&+�E�D�p
T��0�ȿ8��q�ӄ��(�� 3���5��"@�/��O���Wje!��	V�'l6)=Њ�(�J�U,��/�+�z4R��bBn�B8�g��3�K4���d��{��s3�ρ���z ����nY�i´ǟ�2%��Py���9�K�O���*8ze��=m�����;dhM��~c"�~� �3�[� W��kԕ7�c�z�n�$'+����9�����C׸�|���؂��KPl�u���E|e��8�M݃�V�
 ���t��ፒ�Kz��8B�F��+9s�R����q���{ҷe��^��Ӡ��qU+�,����4|~��2R31�h��)/$�s�CQ��h�~#V������H��n߂�K�&T��-�%��vi`��M��/W 7/K{mZ�+�K���4%8SCb�Y����'�W�ظ�Xg�C�=+�k�_�Mz���F$1�_�+c���.UӲ;,q�L������#y��I�������`�bӂPRT�Ƕ5��bzϐ10d��5S\j�2Rʘo:Zbv�Kԯ׆�.���u�L��#U�xg�Mp{Z~ǛK��4�*�3�����9�:�,�A�����;"&@�:�ӧ�7zn?���ߔh%�y4�jN�]�4���z'�]�|_�JGS���[�b�ǫ�B��V�N�d��Ӽ-�z��
�[�SƏ�h��f[�8���`Ӷf��\���=�y
�p����ϳ�R�Ns�ķ��N�^/8	�_�3:��ʙ���d$D�-|�H� UI�lz�<k�?�_��(q���M��@G�{��
�ŋ/�?�>X��s��Ɂ?<�r8�W�
ӯ��� t;YK[l}��Sk�5G^HR/��\�7(����-�ы�$o���0/�!���@���	�%�bY�y�����! ��u`�M~��W^�`��l���_C���mW����ω� �w��.��Z�ӡ�.�s!D���,^*�A/���9ס/��? ]#N�����x:�*ڀ�>'��(Mv�(c���R��E��*�F��U/rJo���wVc��.�Xa�d�88Y&�>tB6��Q��3r���R1c�����.8ME���+Q���H������W�.e'������� pi�e���̕���	�ִ�֫�ʍ$�+��i�R2+�y�c����+�(	�1�'��c��p#B�LyY@$k�l�����,h=���Ĩt�g�����V)�.}
�_�R� W���^�#(���:���v>k�����f�x�_D7飔�/��ʖ�lI�R����ybX����$s��+O��,��������O2��t=I��Y!��9V����HMG�/o�U�Ѳ�#�q'O��E��t�!=��PT�P?�
�^�-gi�#`�f�L�A(�[�X�r�)N �^$�Ŕ ,�{�	�*����X�B
�k׫��Z��>fg9�YW�������f�E��넋.�Mc�%�P���_䭫ꑼ�9�����M�D���OP0�j���)U���9+~!�!B>�5�� �4
@2�����1A���7������/�ӍM'�o�Ǔ�eΛNf_�q�Bv���b�����?�X�:+m!B掅zA����x��p��Z�t�L5]خ�Å4��[�
�d�ّ�y�Ae0-�1�o��L�S 03�@����n.�5����ú�CO���j��r�l8��Q:��S'��p��
r�YA��ߢD(���<��,+�V�ac��c@��2� }oR��ZA}_�܈ 'p��ҕ�
�\���ʂ}.�9��rrE�A	l_"��\�5k7�Q�w5(B���2,��_^n��h�&p'��tS��=��;ɸ�{��L�{W�{4�|c��<���m�ޢ��=)�$�� �F���JH���u��2�D@y���M����	,s�%}�����P&?tlY-k�QӒtYzaM�2-��=�IEy'���L"Ө D���+cF�����<����D�٬�?��.�o/_������I)�_oڴ/�B�<3j���5��gwBz�"�(Z���n�F��h(Y0j�@M�D�P"�V� ��%�E	�*	���=�f��l��������W�6
,�����F5�ҏ��#�;z��H�S����mb����0�F�j�U6���	P"��C�����n�ia��*���*MMr����??r/�Y�}7yY���r�O�eu�"�=K�?�oP(���[�����A:6�-���2���0Z�$��E��	3,"G�� ���V�
B���H��k��I�_߅�\�b���b�5�wU�15�q�]�w.����ˬG�U�ߕz��	߲��H���C�mE��$ŏ0���;�B���^2��|����.�C'[��ѐ��R=hc	`�C��}��SDwc�z�F8�?\��C�픲��l#��.���[���E��v�F�D��	"*��� �_�7��a���F��O�ܮ�96X~T�\�#��O�	*�$r�Dǃ�v�3���q��h���&./��"TW�A9`�e���i[�lb���J�(�+��-En�l��R�:�[�0tS2���X�@�H/�U4A�'Iܹ��A51�^��_��r���� ��G��iY]��:��hI��MO��y�J�RQ(���X�sef6�+�e��L�6��~���׳��q}$�4����Sl����7]S�#��N��Kp�]����#�0Ǚ�~�];�ܵ�B�W�*��!�j�&�<t��P��T�O�F�Ї�%\،�{�ӳ���C[��z��h�Y�b��溉�zI�#7,��v�ۆW�6��L�|�6-��$%/3�n|�9Z�K?���[ȟM��"��!ٶ\�|�٣�<+�W�w�M��3.DΥxʆ���dP�@�5����� g,Iɉ�8I}q��c|�c,u4
���R���m�	*�fg��l�� ���+����&��d.�������f�jC��'��l��:0ӯ=?߱�R}p�G�۰4i[��՝:��f�W# MK�K'8�����G.SrX�٣�����3��a���u�����\���s��T���=�"aVw��ن׭g��~֖(�s�zlZ!�`��D�c)�nhZMA�RG�@X����l��B"�
0�ߠ�"�d��^/{�<Ù�F`��$vv�ɂ��Pao�V�pq�S�Y �eǟ;`	�8I��w7���hP�0#�H8bXv�^>T���Ź^�I<��М"��o�������Lə�E�.�ђ��F�r��O&k`<mp����D�z�r�B��ؓ�7����Mi-G�w�Sp��Y����/`.R,f[�%5�6|x����)� +m�6�-��	�Qy/an�8��r�I�1��ϳ�(��,bU}g%�V�<�h��h�.߼ʾ���u؏F���J�މٕ\ :b�5$���^R����ˏ��}g��=����l�{�ً�׎��C�d���s�?8�jNw{qg��B��A���?�Z-|x.�p��t�l%� @م��Ç~��������[�Uga	�m�Z����F/$+w�y!��f�s�H���I��ǙS[�������R�m!-g(*a�Ozv�T"k��
>�}����ش��%���{>]�����x�9,�ut���(~ަ���6�i���w�@+(_:��7���u7/@!%<���ޭ�`C-x��F��M������
�Z�L�����ֽj�c{`���La��h�OHxp�B_�v���-��Z�P��^�_e��ւ���$^S���4,\C�+M��y\��ߋ���A��0��58|W)4֭�pɑ]>YAN��cXs/w*�����Kbd����f��h��7��s{ʞ���̯;�u��t'�D���f�/���#�=��� ���.�/٩;�r��I\9:�b,�fI�h�g�烙L`�q����1hCIe�nt93P�&�N� �L�MV�|��Vq�#eCj0t%������GR��݊���̒�핝{]�#2��J��;a0=b�H�ʀ�!5��y>���/����%$S�{R��lA�d�%������ ��.�L�H��"֥�z��F9P�����`s�,�|��:��`��5q}����,X����1�*��jW��(2�X ���.��������Y�l����\�b�]3"�3�	o�b��Mi�Lk��a4 ���+#�1���ҋJ\˲�d%:m�L��k��J�&~Q�A�m�<@��?lW�� W���!�	�b��%���ί)r׹"�k�3r�u�0U4v���w(����h�����i4�6˱��\�S�[�:wxFUN��TKe��7^뉺����薤Z]���r������Y�ߝ�
�Sn�gQ��������%U�{���Ֆ����(���D Z�S!/�,��'�a(mC�h��sSܾ�Nﬅ����k��#�!�����3���f$�%�P����c��c�+Ǖ��������[�
�v�!Qο]_�R۵I�oζ׏�;^\�~v5�s�G0�k�ا �1�d��0�jC#�Tn7��{pe?GR�R�i�o�Ą��2E�9"ͼnHYք��t���LK��sP6��x2��y��v*��봤ҁ�hF��0�����e�P���{_�T���s-�G��pu������:�7`����%�f|∑�IK��8T!��kK� ��j��VfoNk�o�(�w蔼F���^�z�;�C�oF��R��]�� �F*1}(���2���h�r��e�nm�e4��P>�NFQ���R-=*����T9D�2�/5�}b�G,��4(@�	���I�#7z��̛\�#wE����idX#'�,�0�.�C*{��R݇��Q��$a�hi߲V$|�y�Xˡ.B��#�,�j4�n�sl�f�@��s��A�<p��P�UC[�
���v�Q\�/�k,|��"�೷4c�ƈ*=@T9��'�R�YI=�y����r���˾}���w�#��hl0��z���x��h岦�( (�嶪�JP�F�G�7	�G��\J��\4r�L�C�XC�v�ў>�fٞ��^w6k�5�*��Rt�R<r�V-bN|%�;����!�5%ӏF�n��W���K�V�\HP9�cI�5k+�6.B��?�HqҀ���2����ۙ�=�t�8�mNqo>N᧹A/�n43��z��i&.��#�0��h���2�L��B�:w�`��(x�}�?0ܮ�ʵ2����i2F���#U�Y�89?F_q]+�rpV�{L�\�1��1)���_J!�t���K^�W}m�2GD؍���ya0�y��TER;V�� �A�gK�m6��bmX��U��o��(��]�;:�\�J�~�~�W�Z=��Ca���Oz�����W	�{�u�G�L\W��Jc�9�e"�
��̼����[����	����bzSM,,1��K��َ\�횘6_�y�/x��+zj�Y��:�pG�|�s;=�O;��\K!0a�q��4����G��M$ؖ�M�ٛ�Ze��B;Tf�=I������0֭�Ve���xV��k �k���{��)��b�^=���������^�%�c���Ye���=�yV�\f���i� �5�s{5�$�~I@&����;C�G�'�:7޳~���*�%&%^��s,�J��D���s�AҎŬ��T.y&�HN�ʧ]Q�À�(�i��~�SL�˗G�q�0Q�gA�V��y{�Bu�P�gG��9���]vT�Xx(�ֺǬ��z�D�i���:�Ad��Yn�L���&8���Ŭ�G4�3�Ī��׸�9������.U02 NJ�gc�� ��ai2
LRd܂��Q�u!��;�ua��_��ѬÑ��/��,}���&���wh{�BY��,���E�L V����מ3P��迅��(�?Ȼ�����5�Ӱ�}_ǎ�u����I��Z��p��,Kg��5��� �~�^�V���R�l�v��s@*C��^���%`Y2-)`GɟQ,sU!�X� 6�EΠ����1�I|I�2E�-ɰ�% �F"���ƕS�	�ڞ�𿘶�u(7��������V����N��T�k��L�2�4�l��^�@os���⽻� �;�eT����m�.��W��}�T�K=�XV\�P$���@O�I�l,Ήu���x4.Q\�r8���3HsN�stn�:;���S�&�z%R`s�÷!���:��^��͎�L�8@
��|���o���=���l��+�̛ĵ
��PU��'�'�W� )6*�p�+�M��]��7y�t��uS��XQE.c�	��l�� ���۝�^�w��[W�פ����D@��%3I�L��Wݳ���]����zY Q�C��������]]���/bt�7��^�6l������f6Z}_�k[�/�FG�S$���@g��%5$�u��COZ��A�Ski���a���Iњ������`	�������Wˉ����P�;����k ���~ˮ��Ŵp%Ә���Jp�����g���l�[띵��kŽ��KԳCӅ���'4�Y�0=�ӆ�#�;>�3�@��j/����}
��Mω-�"A�C�QͰ���E>�&{CT(�1x%�,77�]�G��o���Fu��.`����&��y��������Z=X��H�<�b1�Ƌ�u���D�{!
	b���O�l��M� "�J��k�=:p��#(���J�/q�����]B��Ϙ&��*�`������4U�a<�Q"����{i·�y(��P��
�g�9�V��m���"￶Yx��R0X�=
ݥfaC;{_��@R$f-�Z�œ���鹨C=���s	֎�� ��.E==�����.���N&.;K���7����Pjbsx��ʊ��W�8��%�W�>�p�vhY$J,�����,���8�7Vi��e6��0�cן�z	%��%��8���!��\�(��8]tLGm�e�#��7�ma�𶌯�>4k�����4���C����r������&=O�!�1|��!+��c_���8�-�iF��-�)�ˎ+@­0��S A8�gJ����㚋 ��i(��a�{�&�]{��y�vD��u����%��pxr�QC���h|�tm�����s��u�m�
^��ZB��j�e.D�3�*҅;8�A�&ZO�錌�'�IJ��&���_�u�ꨝ3;p}>P^�/o�
�o�f���ƌI|������,3�K$��D��2�kŦ|���_��i��ׄ��8�duv�FP4�4��é�]/���Ks4dܩ`e�A�j�"��L�m�L�������
��X���1�.G�]�(�}�Z@ؓ&W��(!|�t�nl�veĊX��z���a���2�;���F�y~}���E���g��<M�e"-���r&�Qb�'���Ui��:=D8�,㵛]fb�S�*���@�߲�L4FN��ᐁ�sqB[�3j���E���;^D�S2@�6��p�[�X�n�* �t�1C�{�_H]��d�^=�Z~�y�M�w�ށ�k�P���I��.�;"�^$�+���������6����B��υ-�W� fe្'����,xۀ�����'�i3����=�3�x�^aP��s9��v�%g��"!a��c�i[`"��DXG#b����X��O����j��5<���U�6;z4��N
���rWl�ae�کT��V�H�ȑ)����j�NJ�m[z��lL�Q��V��uvY�8q8�~r�g%��UUE�i;-Q��l��.^��V7IW���� ��j'"�R��;Z���޿��h�'��E�-A�v���Ca�!�f�������=g�4��S#q�ЌTV"4xN�U(�z	�Ŏ�sstpa�p6��W�Y����J'(�-O�f�T���}IҹJ���du�9�8�ĳy��F�j�;CW"�pLj�rle��-[	�9�H&r���<nW�fd`�I��Q/SA�ϗ7R��鈰.�s? �b�^U��4\�L� �T�XDE���%ňΆCG/&�KwUEEc΀�u=Ew��u�}٨u�SP��`V��1l����Xju�h�Rz��R&Sᯣ�&��9Dɳi���M̮*^,�\Q�L	C$�G~�8�~��e�4y)�ތm3Q���0{I~v�����b4kS*	�	�U ��a1_)��^��[���
ȟT�d+�T���Zg�U<�Z���r�e͉$~(�ęi �� v�"�&S�@ٿ��Fxhxy���A&1�m �l��]��
�Et���j��m/�t3��x��3�*a参��Pս���#i���Bj�`A��'<��>½{|<���X�\��}�T�������&�Z�a0K�s��v���*�x���߄ꑃ�t����M_+o�d�b�)e�\S�ixd(B�N�4!�C;a��]g�2`;���J�O��?F�ha�����i������N����H�	0~9XF�O qR1���W�M:ï,J컒o�v�<��'o���=�B�̵�;�L�fc�q�S�{�w��LM�O�`fJu���Ps���M���LPvQ�a�u�^d?u���u��0*z�T?s�D��;�'���DC|
#��炏߿�g�����>�8l�fF\܋з�ٻ�#0@&a�+�g:*�T}��B�BOy��F�� �M�3hh�+"��3���QD���:mW�)�"�m�ϫw�ʽW��
��R��Ѯ�F���D��R�Z���'I!��\R�$[�$�>^��I��5�rk���ˏ�	�?.Ǡ��U�(H��uԴ���DTz(߇3��5G�?����Ҡq�l��y�?�����AWa6�f$�-�X��p�����\ص�G���U'
?��HN��R�4�[���$Bu���?[=A}�e���?�����޷ۡDm�F�n�m�Քpg�L�e�7]�hyΘeTg�kB=������MMR����h��tzo⇫E�ʑ��fT(y��.0�-���ި�ψ�::���/�x��g��U��5*,�� �Įl���`��k����$�E�-'�N;ﲑcޓ����>�5����_J?6!oA���V�+��yj�/��v�l����I�p�fQ^;!�1K}��4�K�ǤJiAӚ"��Rҧ�N�D����A��vzNc��|*ԡn��5hY~s��0�-���͟bfm�u��uK��<� Z��ː9X+5І>�����&V�����lb�N¼��VRs�Jg�w�n�0\��Bf�1����|yŮ���ZW19Y�:Ee>o/���,�|{���׉dv_�`���r�xI���c�I��/�-���1F,4W\@�)g�W��-�##�v��9��£{�n��h�*�=�#�w�S3?`�L(�U�_>=L"u�D߯r��,N�a�l�n�g��<��TD��dU��F�Q����� ������ug��)=n1#S�?��`�N�"��q����іN������Zbҽ�<����F���Xz̘�͇Z�����2����h"b�jj�(F�S�^�%���M�"Ӟ��R����!ʸVQ(Vf-3��B�.�3?+��0�U:$����c��E���ښ�rE�9�w�����-#������EӬ�?��I&��u�q+8>��e�He��m�ܐi�S�1�?<n9��݆aψy~Ѹ+JDF]r�m��XuTU��׹ӆ~����W����;�Fj cg��\rʹ���\��|ժ��"$��|��3�!�VNI2����<bi4�F�g���L�i��f�d[(N�;(��-��V�!��M\�!m��Ƽ)�r�,tjw�_�c�ِ$�|:��=1��K�6~L�i7�YwV��w�#	��h[���GI����'�>���%� ����!��F�Ǿ .����[\-`�/�x%GH	*�e�"��~B']!��>0d��J��*�&��=-��k���Y���Ve��E�����aVe5�Ӧ^��X�Zv�Sr-#��V�0	�K,.��Pdv���򭻸�Ƈ_ξm7��L5��$�h�f�ѣʳFG,*+N;����G��q�U��u�6�b��6nh'(6�G(VA�U��zkL�H��-���檫P��Ӽ"���fș>��ޤ"7�}�c��b�<�=*+�px��1�1�v�i����ꈟ�1j�� ���
�S�g�Q8����cM�L�\E�x�ik�4!�4��b���ʡ�W�����.�":5�̎ ��b�d5Qc��ũ�l�Ч�Ľ�u���q���	,{Sx"�F���LFٓg9U8������<�&~S��>ŀ�i�^y�r��q�D�|�ێ<�-!7�\��MQII�%��fS�!�<S�'��*G�e����V�����OmP`�o�LY��.z��DF��Td��ߌ�����=R�:�H�^���|��G��X���}�Ej�AVm�s��e�z��_�N���mw6M(#��/�������1A�Z�A���I�a�3e�Xɸ��P�y� ����:�	-a^��P	6L� 8�����#L7#;`�7g�~Qh.��P~ӹQBq�u�r�7E��l�ş����0A�s�\PJ�!%h[�-�jEK�|aRŉx�Dsx�Q]i��#`
s`o��W�L��/w�^>���pD���=}��T��X,��s�Kb�nC�Ǔ���D�옝�b��2b�
��S�n�QE�$8�'i5��n�J�f���'�GR5�q�=|�0|���&5��^y47]��*K`NpO��Ix����Q��XJ0Uq<P��3�x��JN,�G-J��.:y��\E ��g�>K�A:���꾣2`� ,����{������/�Q�d�m��ڕ9O��u����Vm�� Yp뼚1Ivle0�tO�#x�!�L`\8�+C�pQ���x쫹1����D�+t)��g�N���z��-#?��r"`��	o�=6Br[�RЍ�?rW��N���g�"�'U�����=��h~��=���x;��o��z���E�n���7���]YG����v����c
jKS-u.�-5~�U��#�	��=6�������X)��k���#rAn/��� ����(����~��Vl��¸a�՛�1�\�u�4�୷����	@��#u�Y���L,9j�?����Qp�V��pPR��s��>��e�)�hp2�
�ş�t���Rْy<�/ф��x~��|v�G!6oT	�5,&G�Z�iS��&�����!�Mf��;�ϩn*�^������'h�ݓk�/_���C��SM�q!<����!閅Lj�LA�Í�����܌���T	s�0�<�tZ� �>iXxX��gʐ���3�Ik��|vWh�m:U�u-���!2��E�@~��v�ݎ�yz�iV��/�e�h����+�b�F/�z���Þ��@��R�H�%�n-�a���}߼�.Vdֽ��Ì*ڔ�8a')����:T�N�Fϝ=�#���5����1}��ը���;�WO�y���r��čx�\>���7�\`����@@.�M�wKO�tI��t%�~Wy�2���ei��&VF"�</�7տ_β�����̰�$�9����=��:�"y��:N��QS����Gh���T�n"�o��P�9*��>1�M��R.`2,���ʕ �����G
��p
u����r�<Uٟp��?w,<(/��W9ZQS�W�[81���SC��`+�s@p�P�����m(�< ��oq�Z�)>.�ϣgF���
Q()���%s����F�~�W	y��0�D\PϽ8a��7�ڎ��>՜��۷���Ҋ[��,=���W�L���#A܉����D�C��$$Y?��
̊��BYb�#ٰ�i6ԇY	�J���lD�T�"�I��iӞj��8�pdr����,��%5,d��=��c�AO��ՂFH�UmyUI�u�QLl��}lC�OW�w�z��!�����.��
����8Btt����>�ZN����t��
�ړ��A�1�0��ӠU����'�X����K̥a��a�aH7pF�M����6
`�+v���g�H�z�3{�p}ruB�R���j�<�%Y�!eȇ\
�A��j�^@I�j��d^=��w��&���`�m�sO�	�+��O�SS�&K����{��Ĥ.Y�VH�F��3�L�ih���O�S��{�S��Wɠob*P�|��dB�6����y����jr��E¡�p�p���@�"�M�M�\�r��pG��HD���{�aG�t4��Wb�"�0��:4�"�f6<ۨ9�
����^��Z�����nU}� ���U+�a}Rڣ:x"HR��7�WM O���aL��;��yx��� Fdډ��ak���ˋ��}�@�j��j��� (�ΞH4Q���l����Rѡ�l��i)ԅB	�����[e��ȆΘ�����;��7���)��4�� 㠷G5c-�]ˋ���6J�Rb�\��&]�~^'	�"ҍ{%�V�=����~s^��YK���RW�%�]$f�W�;��i¿��G�����z]y�4}A�\��^�K��p�*X�X�ND��8��V����O�j���t2O�=�z�k,���w�y�ܶ �c d�YJ}AEq�ʢ��=�Q>q'�Ga��٢%�Bw�>�O��b�3��=(]�/B�D�Z'����)h���H�DǑd{�PAb���e���9h DQ�~���0W0:��{�bB����5z�����=q��h� �_#W��6Z�|
�0�PΞ��F�K���|����ԵqT�?�z^�Hy�/߿���qG:\k[�=���V�$�I5��۞��Ꙅ֬���4-H� ��4vz5�ԝ���8��<o�R��B�e-4�)��0��	�V*�Rw���R�;�b
��a���?�)e�ԡ�ӥ�̴��HWk'߲dݱ%b����V�B���fZ��+�bk 8����$�H�XK�5P	�6�ܒ�����+�|bT�&Ds�.����'�B�v%Oa���Q�5EA�&���E��^h�}��5
[�C�H��a�E���i���-�t6��#�T�@;�#�KЉ��V�M�]B��,�>�S�3��À-?;���o������@ �C���w���@�f��´t�h�w�>�����K���г�f��_����a�"J��9;�C�c���������_��f�U������@�D��۳Cz n�D�����
s0���<�5��z�,���d��1���&�t��؇=#'�n�X���[E{8���u� �ozf)��D���Qw�.xWm�`1nO��{�-�.�4Ev��d\�Jޗ�U�8�6�����ʪ~��k�[�>����T_M��V{s�
$�����˘�PC1s��}�ꍁ��>[�k���ܖ���� ���ܖ���T�Gx0����=#b��N���F]~��O�*����!�#U_��`y�ʠ�ڂ��֗d�x-�9���Hմ�btd��IJ�C�ɿ���һ����b]y�|�@��Ԃ��\�*� t&B(�����N�RK�χ.��kGxv���σ�R��l�&���%�hv�w��噻z�J8
�� +T�A���E�V�&���͏{��j�!��|GM���f7��<	v�t��}.d�He�E��i���˾��2�J:N�݋�a����3��֤���a�{��.*)������G�֌����t�������I��Íܺ�u��_��+���G"�Z��-V��O�ǧ�R�&��FsJ���L��C�)�$�0-;�R��R�0��8=�v$y��6�"��v[�{��&e��Y>6�
����C����Oa�h~��1��I���A�Ӣ�M��଒o�8�"��#���R^څAvsK60�T ���'�>�mGs.�f�قvŮo+fY r�`�B?GuwD$Z�6�W�!�rL��`2�8�V�6k��P	�s�F�[�g�7����\x�$��0�.NYg��1�5�������tp�H�z�v|y�!�?<�Xa }�spʮ��MaɌ}�(P�:�\c�7r0,;�z������%z�)�(Yg!�������ZO���ow��yo,2Կ�B��"	KE(��?�6���^p�`�q�c�M5�#�J=�J���E1M�5ڙZ���/	��8���g ����Y�$������<��"t��|�R��'�0�Z�*�=a�;A�%�P�9��Q�`8��x6Hi��i�LR&��N��]kZ�5��^���Y��锽��$r$9-���o�%+!H�<[5�Z���Ml���ya���+g��'��|�O�ً�E��T��p�J(��Q�)�n쑲��/p�M�A�ge�Z�� (V���Ԯ���v�����k�Џ(�B谫sp�ʷ=��/�0_��n1vۏLy؇Y;㌡넋���J�Y��}_�g�j/�+�O�?�W�QĪ��䱔#e��/���_��<Q��1��D"&T]S$���g+y� ;:N�OL��f6	� z³_9:^��o�$�:��������Y�X�a�L@�}Rβ���Ю�����d!?o�S�0�}�s0�� +�^֜w1�~kf�����!f���GBQ�P�Y�rVB�Շڑ��r]�7l[�c��^�ov#�*�]�7�9�~(atl<� O���4͹by��D����wN����;`&���b��R%����]��V6��_s���/��L�����s$U$�I���(�}�Ź�Vn�^�(N�<F��+R�ɚKr�>#H��Q�����\]�׭ �O}�#�)|�����lU�i����~=9��G�sG�;��-h�������)�/���A�Yjf����M�4��6]����a������o""ڑ�g@ޚ�7׀�פ^�����(!g#���5������R�D�)��%%�) ���TY6�(���I",��`���Lh%�Rfݩ���\/<HO���b�_S+�h��6|�O�?L&"��ƨl<&�L�W� �4�O�j$����׫��>��U��O��M�|,k�g6�_q0�{%'�!)ȿ�TЌ
�w�X�+�Fb�*G�$�f�U[;S�}�� ��:�i��� �c:�,�OLe[�9�T�j��8�#�I ���[�E`EF�	�K2��c�G�EŒSgzX%@r7k�
��;�Q��@uj �%�eZ:b|k���#����t�kڔ�F<��F^�",�f$; ��g��~8�-��l�̾{i�L龺�^�oy�>	����	�-�9���_iU�(�S,)V]��?9&u�~���|���^��&ѝa����ڞ����u��ٺ(�o��e3��+������>z3��-h�l��O���C��!>qݢHy���Vѷ��4$��x�:%��ʁe���rG�(��A��=�AF���@1�����J��������PXH�B��D$G�.l*�_�mN���%�+]�8M�/t����U��2)q�Y�_�l�$&#�L8��`s�1c���L��O����w:pwq,��T�x��A�X����h�7�S�N�O�8
'��s\[��0������I����?'���01^���:h$.5�K(�`v���&OT�(��8{��V����+����$�3IL�Ј�j����S��:���X�d�=O��LĲ�f�3+F�U�H��Q���X4 �+��CҨP�v�T�vd�܊�H�2���u�c��t���PX��(}�&��EO�^�_��^rd;��H���C��욮��f���xޛ�)�@�[�ٻ�E^� QY�Ŀ��h�����cI�e^�}g]�E�ȇ��X�#4859{������Q�s���	ׂh���ᜍ�?/��)'|���vx{ұ��l���gu��W��u`=w�S��\$�G�	#�6�~w��?�RdҸ�Cɑ8�&jo�@dNW�A28 ��9ݯ�)lR��Vq湒��C񏻘�J
���\\1 ���AE�?���J�䭐8`Fa)�驀��Oo������4t�^b�:�*�6�:���+��MZ��IN�
�*�]��<���2�s_�}��1��t�������i�
ǔ�⍧�#����(1�����E�
��E�����c�4�rj�l��̳�g �$�92�EϜ~M����q3�o�ȕ�N��M�� Gɪ+1�,��O�ݙ�֗����x5�ձ�������+hO_O=(�h��A�L����Nv�4��k4����spCO�7N�����HŽ��ŧ0<�?_�����8��gB�h(����C-�& R�ʛ��;!)f"<�$֥���T�%j��׉��ܻU�ߺ����K�B�	Z:����o���kg6�B�9n��?f;'om�]����F� w�r�.���땨��9"�Q\o�t��Lھ�>��ņ�Ptq7S��zhs�Fޮ�ar�	���X��<�/��_ �W'����S:�o�lXH�ח,�G�r"�I-�A�mo�Ā4s �7W�åt�����B��J��<#�E;*\5��ΨLӬT�$��;��ƺ��h%������G٣����{i��� �6ވ�����d2��.+H�#5��V�3�hն)n!(�b�yyW$,v���Ǻqp� �@L�բ1/��9��M�¿}�~ݳ���G����{z���o�+\�?Z���ev˧��@�3gS�K���\�]U��*�g��5ף5�����3�O���@�n�D�LB�� �냖�(?B,I�Nw��tgѲٳ��Sڡ/63��Z JP�1}pPϛ<�>�b�?~��D:r�7���s����Q /&�<�v��)��QZ��ͪڍ�1�^���e�k��]P����� ���
:un�D{�=Y}�4�n�-X�ぼ�?b��}"�r!���j�ayH�"^��y���M���b��"��z����F��m�:���*)�<����B���ᤦ�}�����m?RrF}�Xw��������2�S�z�b��'w-�s�/iQX`�Oq��7&%�z�`�o�f~��ikM���Z����r�o�0���l?���e�v]S���\<ˊ=�Z��qw�SsO,�̩��1�QE ��a}q����.�^ ��ً'n��+��u��\z�=���LZ\b���^��ecDf %���� �c-.�6��H�� � 7X�8�RDfA#y��zy�n�Wf~5,R��4��Ѫr,�lo�Q�/��Ъ���ՂS�^��&_��"h�� ޟ�A�d\������+��l�4�!��$6Wk.#Yl�s߾D�|0�����O�����Λ��9�F�[/��<(y"�̩�x�/�6N�Q�X�|�-�{�c��������^���bg*�+�a���'͟T9�^3Uג*�}� �I����́>�_ׅ5��\�j,�¼�.#]��-ISn��T)X�Y0S6ľ��j��8�R��\��$]$��apKos�,z�!i�o�I���"���f�x�����NE�_�>�ݗy�
�����l �C�o�T0ҽ1�)�[q��0�䅘���ϑ6�.�ЭE��Ϋ��ܺx#����+��oT��J�^�V�b5+qV�ur@9�9����u� '��_����<�i	��~�H������3!��_<^o�'�p��W�e[����k�H������Ee��tY����~u��Z9����I�m���u�'r|���a�y�X�wH>���M�J���-Q��hqYQ;Gw�q�#d���u�hG�W�Q�I*y�%n��������9����������Ȇt��i�8�{���
EΫ��,]���Y�?t+�e�]�՚z�"־���NI���{���$�!a�9�܇��`�Lo��h;&)��1O�4�D��g2�=_hũ{��yR�V_���<����k/e��ÿ�U��9l��Vn����@��8�&:�l8���.O:b����J,c)f��+'J���'�]R��:��-��C�t�x�\��F���zd�m�p�s|ހ�����N��ޜ.��h-�PJ
��Y�'ϴR�4?��(�[E�ff�6%��'�$�؂���L츥}W�����􊯟��8�p����dg�3}���#���B.��R2k�AX��"�A�|�}���O�9D�V����
��CBC�K�g�x<�B�T���5(rQ4G����Λ�܁��6=���ު�2�o:E�ؘGj1�E٢k<}ĳ�S'�m{�#W����"��
]�ƣs�)F!.;-������6� Y�]���IU��c�ZWZ��"5�ed�|~VD�OuPP0��� 9�f5i'�i�G~�R�/,���M�4_�j�P�Ъb'8Y8��T�Gu�L�YQG�YBT�!G���t���G�O`\���� Uˑ��(��I�]\gq�('�5�_#�yq9磖%��)5�����G{�� ၯd������f0R�N��X���6��t� 8aj9��h302�D�ː�oW�t��%y�8�oE��y�v� >�4�	]�	12?,��9���I�(�%NMYЊ e+E���e�x�Qy�{pb*�����UQ��d�;�PCv��R�%0ѵ������ܒ	�6���YM$;XV"�K�����2&�6�]�;�m����^�X�R�!��2[@�ޠ��J2ب��|܀�^���߃��>
�k�`]�Wi^d�`��?/�BN��y `G���	���`lg���^����mWM��\�l.�C�Ə�j��tw!���/$+u�a}3h1.���垆�h��Cd��4��@��7�X<�z���z�a���s���Me�il���PT�e?� %�!��lf�R!�Rk� ����e�er�a*�7�={&�L����L��ұ�^��r���C̎��Â;֋��
���T�qߒ��ג'8.��'��������Y����2Vk1���ل7�B�� �d,����Oߘzi`?Z�I��lp^���xUl�Ӟ��?n�i}~{�k���,T�1�[l���fRq<	���J���������?�F\�e��g�A��������5_�����T�FA`��cğ�}��kq] ��q�]�o��
�\oLU5�y�� �rD{}�߉�y?:��3o���-��p@�|�z+(d�S����F��V�vU)�	hl�}�(-Bw`��W��<�M�m+�4܌X���ɿ��C=��𬭳�Y܂�9B.Mi"@��n魉W��r�H���t���+(�[���-�K�גa�Z���M]p#.�:�Nٖb���H��c��M� I\�#M�%�~�Lo�/�q5�/��w��`��9���>_�YG+ΓHٺf�f���t<�Z�7~��hr��n�,<?$԰sS�}�y8�>�C�+��9��z�������p�ݸM��X��qL&#nB����=�5�:ϱ�g���O��'B�COe�=9�Fg��С���O��%p���3�U��X�b:�4Ck6yV1���ʙUb~�Ka�;��F�wjh�?u��B�����tIu��F���(1mCܧ^�QV ������=��̽'&����U,��'��#,�h=�?Lo��D���F�{��E�I,ZИ%K����ES/n�`qm���-�Fx��O=
޹>�}t���M8u���B9��C?L�Nߵ�/@I�T����Jc�ی@e�AP��8�W7�j���%D��7�ݦ�1��^����\��=�J(*2]r���@��� }���e!�M�E�>W2c:���(∹&�ͦ>��{44��6������Ģq���U��Lͳ옴a¡T�ji�� �q�6G��M�Y��(����q%�K�І"�D'����.p2P��W�60h�S�,���Н#�l؞}���*����;+r�M�k���&���}�h��,?^*8p�����H� ��F_�4J��h�g�M\o��Y^�1�b,�b �jڎd�O�	mᮂ�@��T�G,t��fB%@`�fGx�|����Р%l)K��-���6'\?J�g�°O�SIgY���F��I��wFF�S���0=���tCG-��S[+^���b���Ҕ��	d�o��-磐�@lV$��)��;A�{$�E)c"#(��k1�Ma`�VD�aO��GS��CW����䏩�j���!H�(��b� ��l�Ҋ@�3���D����F���
���B������(�5ii�w-Z呱[d�w��L��M�B���Fϸ�v̄M�7���Qs[A��D����1'wx���|J�����e6�0`���x���$?�L��[��{�z�-�>��z^� �6�,��"�[L�'�f�L�����.�w@�~��D�9��(�Ku�M+��򸣯<� ��[��b�h~A��޷���^s���S�{�RJ��wX�.
�x�l$�!�8��e	&	9)d;[�]A�����7Z��Q�w��P��'���v-�������t@��{�OZ/p3��e\gD�6my�5�<!�;��]���j$���t4❮
� a��#�RM,�ae
���0H�	j<�����#�fA�o�5Bf2>M�on��Z��)O�'⫵%�8��QgH �Ȕ�m���\��mN��ʗ≈��Y����Vx���_�:�g�M1<<G�f/� ��0U�8��5�8Ɋ�J"9�,v-ڼe�f�����{ȥ��Mݻp3��ዛ ������2���u�A:~�+��f k�]x����:����{�+0������a%!��$3�7qDc�s?�8~����z���ܲe�hÔ.Y�sG�1(��.-A8g�����xG�>�+D�G�����1"��^q�ֹh��#�qy�j���wo�Q+4:��)O�+�>G����|U܏yD�0�i��Ƥ^B������;�%�b�T��$�^n�� m
hƤf��i?}��U��č�$���� �vWMycʘ�A
�i�TT\�J�����y�w
[fPn�.6�I8���W�գ�E��xNn^Wo���1��C�pF#|\ '����y��ӡ����v��'���e�OY�Մ�'q��y0������{�(�<$�T7bv�-�[�����e;9�ñEw_��G�6�����7�N�$��MHD��,���&��b#�e���~�!�n�.P0J0`�4��hͼ'M"F��c(EH>�E)3-h
5u@�,(qć<�S�U;J��,Id"�y�f�����!]���\��A��a����X��Ʃ��{���R=�b7��&IyroJV"�)[,���e�HɟhG��,�����`�Iɗ<W<S���=����Aozp�H��BT�^Ôú��S �Eo�H�v�q�4��ۇ�Ӷ�'}@n���Zj��
����Eݟb����P*��lW�=���/p�j��@r�_hEcfE��v��3��5x�E�B����]_5$��x%1p,ոs=U��"��T�.a���A���D<�F�>%�����9�Eӊ�`�)��45�g�o�<q�\��@���N�~#D\*f��q<i�C�E2�8~�	�~�q��F=�3�"#�b�A�Rvُ ��p33+�&���w@�F��L�4�ùE	�e�I�� Z�_���`����+�4����d�Kxmk�3sf����coj�3��eT��&˒9��݊F��`]u�.��1�EֻN�`]�׿��o:h��]8���� �P��x�����G��S��<4Y��?g�����j���	�>4�;�+4A�-�_�ΰ�H��/�Q��u��M����D�]R��e�W����>I��c"���7����+�a�v|� x�A�a�ѩ%
I)���y���R���5~ծ�4�9c��Mȥ��r�vH�a�c�0�:�m&��%�z/`� ��:.4�v�H�EQ��5P�.�|R��Z�U�<>����8�WM<3e'D�/׫��ۺ���ƣ��8��$�z�"��5Wp�?�H��������Q�l�y�Ij>�l��F�ǻz[l�L��߳[��'j�Я���鱹�J�r���X-S���l����?�|��Y?�*��Qa��<7�$y�d��i�Y�Ki\g���-���� ��ʖ"K�@�aQ��w'&������A~�|8�aɷ��g�u.�r��zf�l���?O��ll?dQs`�����É,����~V�i~a1��͔�h[_���S�;�H�B�kX�s���C(.薪g���ȵ�=�Q��|��jz�1��ڡ��i�ac0Q��(V�r��I/C��^���#<��5�>ѸB���ᰌ�JV��8>-�8���5jI�m�Y��I�UWDB�xlV����`�HVX��y�<��������!�.����*��V[�y{�H�{f�l�<%�D?���{��ܓx/}�.Nq+��!7��H�LI���u��.iѸ������U�
�H%���XqO��|!B����&ly�Prg;XDM.5��J����آ1��Ԧ�d�i�.n����o7ߟ��ʎ����$���c;OP ^Fl�.t�ߨ�툣�9൪P�xN�u���̹�.d"�a<�h �Ow�UŒ���/���Dw��.I�Z,2��P#9�x���������C�glaŒ�F[eׁJ���I^�u@H����LW�9��������W�x�W)��*A��Ws�`h�ϼ�� ��`lꮰ���&��X*�xd'f!���q��7��Kj�~�(5�0�E��K~���4Y���MF��O���������e���#��~�+�T���@':��������g�i�{�j�&Z����wV�� )�)���:>��1���;v_Č��z���P��3�U�`�	eb=�H.�S��w�'/�Y�`��;L6�%Y�?�����U�e�iɺc\|w�J�1�j��,4&�Q����Y�aQ\�k�%�>б�w�L���'�`?"(��r�I���t��Pg~��?�	³t���ߘu�p�l-.�s�nj*c�r���ooС?pY�>&��_Zoe�M�m���f�,��
�ƭ%T�xq)+X�$��6M����t/�� J�N:/2V"�|�7��]����1Ok[��Q5��Ҽ4�]�f�JPs��s�dz�h�T��V�*J��Q��y�S�0aT0�S��M�:|E�t�ǈ�ѧqº1�3@0�n�E`(~��b�P"ᩙMy�{n�!3%%���\�}x�b�WL�/�N��1W����Q/lE����ozV��V:.)�Ϧ*���xG�n����EdN�3`�ʓ����� V��蚭�T��R�_�,��U}���|���9�C�ȘhVś��+i���-ys	�\����O��XX��v��%CX�����c�õ�v4E�}�R�3(֢�4z�]ȅu\_>q�`�qӂ*����V��X�$� ^8'��.�2�.Rw�1�P��27?�G*�$��4\��M�A�Ғ���ԩa��~%QlI%��TO=��D�[�����ҔˊG׻��?hC�����*�x���oB`ћ`��_D�O-2=�.�_�x�3���	���[�؎S�AЮh��=�����$��m筩��[�����P01Te�6����Vi+�E�W��,=�3��zO��!P�tt�#��'�ݖJ�'B]����V��4"!��$G'�q��\
	Iz�o��0ڪ���a$F�B�O����].�G��tS{�Y���I����guf�j�Q��?��A��� ��t��xߒ�CP�$I���PoRw�ˡn�qdfou���c։�	�E�n2н��j<�g���ו}�'*cU���p���x�6����g"$�HWՊ27���B��]q��4V;�5gJ����	+��9�W)��RR}�Y�n��P��{5۹/�sI�$�ˋ����9}}񣧍L�2�`���#P0E�N�7%#<���tL1CV����ZE|�&.���lH"x�Dw! �WD�m�Z5;~qCoB�v��K47�5{�ڼ�4HG�;G�	�&�y�$�[���Rof���EǠ���Z��J�%VH��>��0.ֻ�`�)��}Z��:��1#d�t��V��"O��&�j��/�Rt|�3/��:28&@<iqs�WL��|�ILط��G�<�8W�@�õB8�k��hb����!5*����%��A���d�څ�Ų����ge�N��*����~+����.�g�u��p=w9���X�xxR"�hӐ��#�8��Ϲȉ�&�* ��̉�\���h��`Z�A�
��)8D�m��#�;2pZ�0Ժ_�9t_
�^�3Ѩ�i�S�y��OyA��~մ����Z~��kR���I��(9�F~��oH�jj�eӓ��V�Y�Aʔ�n�h���ڔ,fW�mtt���/�8��x�7�GQ��2Z�3>��d.{�ަr�	h���`K������s�L����m���߷=��2:,�1����� e@�	-��H���\�h?՝X+�ָ��@�Ƭ�����1����F:��<�В�'�]osl�$��� *��:&S�ҍx%��;8Q.�
(��I����_��Z=��'�q��)����?��+��	�ρ�*+�Xo��m�q]8��n�������T�(��M�U�EJ)�Wfg��i����P����5��ϱ��E6�Wt6��6ұ8��~��\��E���Qs�~(@�]|o��sp.�������T����E!kj]4�Ϝ�Ք�4�����aUIV��Ov����l�˟C����:����>�j��`���%�NV�N�G!�`�A:�����q�&�XJ���X��j�2�F^���זle�~��(��%�ȷ,���4ػ����R�C��gҢ
`���d=���L�5�@r/sHx�g*�1��6����:��x;9�c�Z��H�4��;UaO�^ѓeG���RA�Z��F��e;��d����Ӵx���h_�f.��$�Wm��2uG���`4;����uF�<s�>��ȟ���1�M^`�=,�x
QP���9s�j�讌΢����xHh���HØ��0���!<�χ{��ऊ��V�Mj��MR�w��곿����Y�s�{�d���ޛ�؂��sğ\���?�\��w��_�ef��/&O�N4�q�Đ�/��-�X���J�K�����$���@����(]M����v���7wo	 ��	�|��d�'r�ѣ�B��Xh��ņ
c�a�v��>i�D|���ďq߉j��2	�R�-��%�:��8�B���W5�6��B�1�|�rKH�G{�:o�5�4��W��G�׉(�
SH9%���%��5�Y��e%���cXu���zl�to�!�-n@2�׊�+�.�'��B��]5�	��F�ze� 4�l��׍�v����ed�)��Ӱ���Kۦ퉿v���.]�� ��-r��Ou.���/h�����0�v����k��І*
���[~��|�t�A���&�z½G\����8�Y�L����	����U�7�|S������=1 Q' y9f�h�*��k-Ρ�t����W��^�S諾hK��.��PGp��2�J;yI\{_������K �#�}>��B������$�e ̮��^̐��+�}C��o�y���B��1L�h(�i�v�aA�� �f_����Eg�*�A�h[ɶ����#-�1�X�~�A5cx����{��:��Fx�Qw��_�
�Den��v:����ğϔ*�~(FD�U�,�g$����a��!H��~-L�3� Y�p�4��Ub���{(���o@ʔB�f]ǿ��I�h�u����|P�`-I����У�I���s:�Z�l����eW�0<����� Ō�L�̾j��y@��������ðŰ�G�T8K�
~�x�9�fQ��x�x�{د�^��9��E��+�;6=9PS���W��қl��ߨ�=�ن��.�M������?䳯8J(��m.��).��BF��}FA��}��}.0ލLl>cҼ��00V:ڬo!<�s�����������������ҧTl�z,І�V�&�ǎ>��V0V��^�4nU�8'���ƻ�+�5�H���J����a�9���f������ME׻��r�da��ap�N:Q,՚��dVD�&q~�"��g(�! �ӭ�L7���u��J/���`�����4kW���)��l4��
~-��+�_q+&q���O0XH��bJ-���v�!~��+�y�p�!n��WT��u�=�^K��wx0�e�@h;��b��~q-=> ���R��<ل7���A���Bj���5\�sN<y�h��
�nURR��x!�!(Zh}�\&���"@x9�A���`�B�ތ����N�g���J??���ym�: x��+���(l�#�>^�"͡�ϤM$�q��%�4-ܢ�%���1��8zC������ғ{�%���j�����f�4�����z�F_��~�� 
H����y��7��I�
a��8p!CV�c6�]�=�eF�u���s�N���ū�5�g��rZo{�9Y���@�-2-W���ӧ�a �M�����]-���+8�)�Xw��^��d�k��'`�������,AYՒG�g؉�#�(uA�ܬ��9{V=(Ɠ�>�=�ȭ��������4Ij3�g|Ah957�ez�Z����v*�p.Ɔ5]SJQ����H�x�9�w�n������8�C	"�xYk"j�^=�RG��ׇ\�R�߲��Z��۠)|*�c�"5.s�Q�Q�
���*���:�-g�/�+�4��}�<�y�-�b~,$E�n�L7z�p��^F&�$>��"��+�uu��$��������NC��P�4�A�Eg�w3��P"D0�������h9k���=k����8;+ű2�n;��Dq)RR�˔a�)(��x}͂���+���6�S���W�_?p�@��׈|�C\�ʸ�%�+�	fY=��d;�s���"��'��0��J���L�)gQ�?�8m�s'���{�<�Zd��4�~YH�9�S=��%�%T�{��zk����/��:���i_IrR���h�A����Wc��-�	��U`�$��z4�Q��G=�͹�׸4���p��zN �����џ`�F�W��^�����W�(�MW�I�la%1���h��E9��1�G�o��OYx0k/�ejmP	J^E�n�U6n^�8��OW¹�wڌ�7km>����*�/S]�p8�#�їy��B��Az�$��Wx��~*�MҲ��;1�[	O�j�Q��f����	*�F^��l����t��M�^����7�)q(��B�Շ:Ug��He[�ݹz���:;�S��w|DБ�K<X9����&8��4��8~�������A�H��(z�~{��Y�SU�`�ե\���5��e�l���r�?Z������=��I��2�|5�
"�rs�׳+R{*̺: ��B797N~��`%@$x��<�c��YA�KX�Г�k��|܏��F���Р�WMǲFM�o
�BU�Y��"t�]j�V�#o�����c�.mڎ�i!�rx�Z	e���e�2�'z�h^AK�����ٿ���ǂj=~9׈�(wB`9n��Z��3�.=*�M&���H��}�]v�K���� �F2&^�d}q��8+��`^2p���4���.�\��:h#����g2B�ɤ_/������^,�/eFυg5L�|M���}�w�X�D�ό�Coy��ϣ�mg:wr�0A|f�M#3�_B�z&2��,F�4�m���Z�Gk�����ʐH�ދӝ���*�2A=W�0m�6i�B��ꞥ���6)��H��0,D��Ds�X�o����v�g>0Ր	��qp?7Gu����~'F�����a?�sx�2��� �u8W+Ē��3��#0�Æ)6Iw?�����
�9�l�l�B�ē�k�guX�_ph���Y�&�DY=/YԄ_k���{�*����e���łO�,����sw6�[44��կ�59ʉ��㾚�s(�0��nGd�$Ħ�⅒Mrg��9BN0�)��<��=�d�#��YtOCKvbO����6a���Oܘ�0�#TRD3���~e��:xl���j��\��TR��)c|_l�`{޸P�ӂ��.�L�.�0P�6�9Lk!#Ba~��1��}�@�G}��"�J��2����"��¯z��,��b����RIOb�]�C{�Ҁ��=q7��6h���*hC?�7K��;{����8���RAk�� ���D��#E�� �^���[�6��_0Pt&Ȓ������p���q�����{������:�k��[���(4�lˢ#?�/�o������kXK��ި��y�T��݊��|i�p��LJ��;�EX�;�֥g�+h/�&@PEQ5�Vx2ą�c�N�1��q��uSJ�D�R37����\�����Ŧ��Kʣ��fV��<��j0W��x��($�D�g@��'��`�'���t<��{A�+��|p�S���qk-��Y7���XVb* �i��U�'�W$�/�q��v�f��VE�+��@���p���M�-��y�m��h1�˃�ڢS�e�=w�d��W���"F�g.a���pj�h�+��(���t�K*F�zo��ό���}Y��%�Á��_u����|�x����Zy*��R�6�[��0��ry�[�v�K$�Y�A��h�	5�qa��` ��	��)�O�5e0�U������gV�,�b��5s<]SP� �F�B(�a���_��7�a�"�l��}w��2	���m/�C=wv���C4���-�RE�5\�N�Sr�j���zG�	�91�^�F]rΤ�����tai��k��}"H�	�G�F��X:��:̏j<����Rjb�K<w��C��"�B6���JBQ���G��G)��>�#M� ��Ó�9.O���g��7V�<jms�!�?�;�����ߟ�檂x�E�5�;���D<5�ky�5��˒���s����ط�%AϡU�cNI���?�����b�e�t���g��u�^�Rk��jp�bg��%�إ�ĵ>�S`�~T��f1d�����шٸ1��07�Ҁ1�^'O/($��cM��i���@�5�űۀ���k����ͳ)�y+�E�S1�Y���ҟ���Q��ܱ�{ %�J���Y�||O�����c������<�|�	��Ѵ-��F0��2�J#���Q��\lhYJ,oľ^@�P�d�/���-� ����yz�������נ<*#��U\�#��D>{/q䇹�Ǉ�0��Ȕ����� �O%eM���;�U������N{
^*�u滇�Ua{duv���v���M���\.�>@H�^..���0V�!����/��O������� m�۳�eI����V0v:P@^x����x��iRl0�ّwN�A���~c�g�qo>��h�&?��=#�҈��/̌\���1�8�6�m@\*sI%�B��0�,���C�TjAf�(��&��R��r����ᒐy�;�%��!�I�+v��4�.l��a�;��?�� l}o�߈,�>��!�b���A���sV���q9�~Uk~�i!�Y;4��z��=%y�/� �bJN)��؟�c�6�)�Q Q�H����BI��f*�ǚ!K W���x_h���$!�C�E�ͪD��L��E/���r�>O�à)>�z��ԋcOPn���G��T�-~]�r�o�#����00������v�|�L�Xc�����V���Β�&'EUֱ�P��4n� �mQ�|��� �{����+4�蘷�b��֗�k�%I����V�ؕ��'��Z�ʣ��]HLX��
��z2̻�~I+
+��~2�ֻR�i�2�[Z�"�FU��ŉm�y��� IْBe�T;YBD����-���faR�ʶ�=%�zޮ�+%��^<��N�����7Պ�vf��ay]*���_�1� OMi��%��ڦ4X�eʢ�:���ۥx��jO&S�����SB:C>j�c��W��]i��Ȃ��-�a�*R�|����ZZ�|�a�9�"��<m��&���tzv:~�#,�9&�{��CE|��K�O����T�������.���ۥ�f�tEў����lyC{��N��O͆݉���ӲI��X��и��7�"����é�o�e3�5M��8&nA�W'5�рu��d�΄�3��� @·%��:NZ`��W"���Ӗs�ר�k�U.�y�+�B-\��*��s��|x�j����(p�=K'�l;UԎ���07>=ʧ�]0/7���*I�u�ר�!�E���m60�z��q����|j֊�2��[��
�_ժZ�ƥ}v��/���FG$��BJ�8?�b�Ro�23�����D`~����4�#�����!G�r��_�ʦ�[�(�M���x�6�	]��5@�b��(- E*�,r�1���E���n���ק�CV����K�O��k��M`w& ��5{.�^�!1�,��כ+�ɮ�OI��X��5@�ϡ��&�?�PN��Y�UaMr�x�3!�r����� �eIt�D���,	5N���.Z�ѯ���$�&��k������ �O��1q��֫�JV��N\�0�ܱ�-�-�^���1��o�Q7:j}�|��&���<e�Q?{��l���[z�`��'�{���K��s��!����5�E�V�BW�w������P���"�Z�Nw���)>���>f0�w�Z�a`��[^�D�P����5�_P���3
��L�I�b�D7'�y�S=��Y�-�.6\�Ȉ$�Q�u����xg�z����Ss�4�g3-����	�,{r�MSKc����Kuk��~D���|����i�'�~DBV/\ �Q�z%�!���/^E�Nyl@1'Y�� hn3�V���P6����,�z�Atq0o9���ˉ�S�H#ӽ$�������*� 5��O(r�=�;DV�y(	����9qkSK��;ں�+�g�"h�(��ו�U�.JA�
R��y5��qh��W�47+� ���YA<M���}����aA��A��5�F��>�W�ˈ�DUR0���g'�%H�$���#�|F���]Q��?
MH!����o`�+�v� W$!�����	jel���
F��+^t�Z�L6(�_�T�n&<se�Y���H������pA}8�SR�G)0xk4�X����Y���3��z���]w����̧B������bS����BroAۣ`��+��,����}��C
�u��8o�9�އ�1����Tn>���-�f?�b�5��\٤�d��	h>Y�dwb�C�J���	�M�J��n�#��7��3��k�}�H�D6֎�s�����/��@�N*p
��'(p�D���P^<�n/��b�`~LC��e���6Q@�� i�(]m]���ʺjy�Tc����k��:gTR��=M��U��u(��:U�Z- �O�{�2f	3�'��-|:Yқ��UyK���E_��WJ4X���d��(�"SAxڙm}"xO;��z�����c��ۢ �nT�_���V���sfs������v�KGBQ��S���d���t��kA�?Sǥ�U�k?,��9���S�����kj��Zw��]���^[������"�����������!�&#��ञ�kEݺg�;.�E�m���m_zt6t��:r�NO����f�ka�Әh�g�в ��z��n��6E{��D�� 	���������Ӕ�SPj����Y�:V��(Ig �]�ma;.H���Ǘ�<C�Y���(R�#�Y�Qf
+�� ��>|�hP�1Ʃn]���ўbEӎ�0¡����`F��)��ڕmA�a���_.�� 2���Թ�Р�`!Յ;�?�п�^����C;��~�4a�pԀ
	��aޒ%~�K��	���m:�'n�I_���/�~���Qs|�:fNRtyP���b�$Za����܁i�u��f��ؓ�'v�����#�~)�/���l������ӟ��$rZ��2fEz}��+9�^�'T�H��}'�y�is�7��s����{`8̟ۇq��y3�{P�B��)�S�䌀�M�UZ\�o��
r��R�LK+k8�6���N"\<������ؖ�XaU�_��P��Ky�oT�]H]�)o$]��<܀��Ny�Ϣ���
ձ�2���D�a��v���j�(�;�-C��'A�軧��������o���kʞo��`a�ǒ(���'5�p"ۅ1JO��F:Q�ֺ��i4��p�ឹd.
��t��)�Yl_�S��@쥥��x����`��!ꊊ�Ұv�h��kiK�U�.S!�*q ����
y���0��|�A�$��ǁ��\�Q�}%_}���\?�����q��Mw1�v�I�}�	�È�Xs�.,>hi���IV5���Iiz'}���aҜ�'㮑>��K�`R!u}�G�{�-;�c�8�b�]צf�q��jTG?^��t
�ș�� =qב���Z4���,7u�}͵��g���[{��#��A���ޗ�6L�Ű�"���.O���D�"����Pt��(]g�S�rG|T&j6۫�� �q���vQ�h�W�����F�֛���K[lC���<�� v�4�?d?=!gQ3�4L��^��ʓ�Cm+��Χ���~5"Js������P�׆A
P��#g�CUn�f�@z&��A�wK%��I
.�8��Si�筟��us��	,�D�7��e�N̞��}8xJ��s�N��6q�/�R�r��)=d:�g�<��X�#�r�"�;š ���s�g�7˰v!�Gt��qƼ� �p�a 'm]
��r k�8�f�t���0����C�$H��\^�\�b�b��l8ƣ~^��_��Sɝȶ���LtK�6	�mG�܀�(�*�s�>������1�8�&Ys�@����W�m��}�r�k멑eǏ�_�j�����P������<`��%M� ε5̲߫���N�b�c����#$_���L���s��5j��<��8�hTH?�J�7����X�΃�ߴ:�gy����|���K�8�ʥ���D��&ٟR�dw$��ޫ���+BI�.E/����D�W�v	���ݗ���$|��=�
�FɕnNw���k�Sۊ��N\�L���x3�W��v=q��˄{L����6���_/ު��8��Q�ɓ�D�KVc|��2f��֞�`>�FcmQ�/�������[��R�)aD���4)t��5�釂��G�����{�Ȉp�(D���v�(Gu/Y@&��+X{��j��aI��z�M�0.f>���'E]u�(NQ�<|L���I�i��D{�H��j����S�8��P��#b8��_�7���$
�1+�(�-7�h����1���m_��y�ޚ���^K ���1�8�Τ8m��'5��a<>�nbD\�t1�DQB����Y�d�\UP�~w��`Ԩ�Td,TMld"
S�/T�vۉ�3��;�a���r].N����!b$^�3WFt��C否CFzX�c{º����R�O��ӕ�^v	�hH�Ѐ�!�G]N[�q���D�[5�K	`����W��E��hA�h} �������=ʟ�{1�R�ܽ9ެ�8�t�Z��s2&������
�	.�6���,I�����9Tt9����%({�j2P��Hl���OmT� ��?\�S�63�㿛'�'2X6R��і���$�=F����u��`[(s�ׁ+J���v��-��OOS`<U���]W9ӤApTFDw&�/��T�j�p6�v��'WT��ڣꙛ�.Н�i^�C��&Ź�+\X��tF���[<t�MZ��A��I=���O���|�m��ؼ�w<R�d�|b�?�A�Ь�6 rWjB���Z+�֑S}ԣ¬�q`�~����4�1�8���w#VH�R���|f��m+	��ǳFHߌ?�u§����L���A�Ags"�%���n0簩�/C��&J�[_���X|4��å�c���?	��g�����+	�Yq��`b���V	��h�o�����Tb#�D��b,i���&�=���ǊqQ�ܻY��E�hm�]e��>��K3JMmL��5D��r�X�p�U2�Q;^	�djN֘�G���Ӣ��P�e�����?���E�!�S�t>�0�����7�}�l�_"(���P�r�\��\�B��%�	:!1�e����G�N3�n���g��6f��ƲK�$-��%�]��H p~�xL_�B�^n�m���V($L~�y;���͠{���؂
�Y�x��_�~�%��)qҵ�L���c���c��X|�0� ��'�]�q3��ƾ7"z�0� �݈{\F�H�2ė�����j�$�w/�iʜ3������ߑ�a�} i-�āfIcu��9�6�8$��aZ���3�V0X/� _�yD��� o���~O�kQ�!�(ߐ�ڶ�-_=���fku)�*����Ő(ceE撶g�����PWY�D�)"����oЍ(t���iI��_i����Za�^�e��T3	D�S��O%v~�Q���t"i�r�S��݉��r�Ő�3�:��a?Y:8y7�D~�l�[�ɽ��g������������ߗ:ܵ/�2��m���"t�V�9X�_��S �� �*��0�R�7��H��w��Wׄ؊IQ�+ ��$d�ӒKm�e\\Z��3���ߥ|�x�̺�u.<<}O�T�qK�)u���Z�H
M��mP��vw�A�����o�\�*�۳_��ss0�|c�^t!���U���b�%#Q;#�C�=V��y�r��^Q�n����ڮWw��󨤅���]v�<�z��x��sҖ�1�tX�)Yg1gN`?`�'[���@�s?�S�JhN/pd��<���	RE�d�C�2z1�x��Yq����0H�@����-4M[d�8s���|2p��t���P���a�,P�"�E��VAgO"���I��-��&��c���I�IZBz�YW�6񯻝�j��i�dRipw�O�� ���$��L�f|F����j�I�x�ǳ�C���(&�ś��I�'�X�&�)��,���u�Qa��U�+�^�1h�JڴI��W4�HH�$J�2AX���bA�~�5����M�VcsU;�δ�_ID�S���i�k���$���sG���6g}�Q �!d���|��_����tSl}��>��G���$P��Ъ�2�)<@3V,��;�ւ����c�BX��K���D� �����%Tm�D��ń^i��b}��>�Z	��πR�Ӫ�SV��<�A!���l�=Z�s������:�T��	�2�T J���\��Dbe�}�2
O ���y��
A�*��g/����/�m1��3�-�u���ߩHG��j�{F^nĴA�°Y��?�(Ղ�*���4��,��~�Z`Q<��n|�l"S�,E�/d����ߤ��3���K����1"�H�qG^��l��D�
��ޓXڂ��/�/�Wg�%��~��-l��ˮ��7���G�9�-j�r戃��L��gꜪ|(�0V�w��M,q���J�63R[}�23����x������q6�x��p0��+G;�"���mg� ��AC��������Q�EZku�fm;^f��0z�Ds�V��F
�n���1�V-׶�_1f�+�6�.=	��gBO�{�`�{��݆��j*�T<q�E�9d.���P��MC ���;���|��A���#�=��U��Z>Y��$��\��}����C��ۄєb�Q"�3`�I��L-�l��
�(��3�\�i m5QG�:���������9��i42���E�6R����x5O�7���W~������?H'.R���ѝc�K�� �����U4!����Of��q��w#��}s,bW#)���w��R���Q�D�HxC%�պЄ���~�Ҽ��֤��^�,L�[��B�oA���Ci�w�#t>�`��S�9^C�h�Z<�������)G��؄J����p֞s�iSN ���uZ0���+U�vR� �4G4�W*�=w4����3I���r�c�>;��\�9ѡ�7��)}iUji�Ou�����
�������!��v���@�_+��l1���y��mgW��9��	�\��Z{|�O��t��ǀX�'}����B�Q��0@�#MN�Tv䙠�����n�f72�X��y�!��% ����k�,���
��ש��M��j�� k� w��2�	&���Ҫ�q���/�3�ӕ�����S���Ʈ�K�~ꕊ��8�)�����y"�HgN,���R=��Z0���$ݛ$�5:'zv���.iW�ۜ��e�ߩ(
�h)1��]���^WQ�c�`ۡ�e�C�v51�nF��p��\iάmk��-�ð+;��H�N�0���zlO��]C�����V��+��/���e8����.��O����X^ʒg�����Ѽ�����1�#�}s�ۢB���R��x��W�a���-N�[���S�];6����'�"O�\�:��Ii�ɞ�9�	5Lf5�3�Mq�)�Yݛ��!q0��?��`N6?�ṍCV�n�ӃkE1'�������aط���S3�.Y*K�X}�I��Q��Ӈ���?�j�O�7�偅�Â꼫��9RrFV;�|����z��\239 ��Sj�o\b��4�_P�V��g-��������ռ�f�{�]���T���eQr�8	i���ݘ��GGZ�@x���,=��`:��YS��>�{��R�J,�<��I����Y�����>?"9i�.�,fA�3IT1������4�am�}��%b��t�.�h��7!Q_�,��߿�J�E/3���rG舨0zr���K��&���q�*ZkS����Y2�%��0��r@���O�,�螢
gji���r�1��S��⯅��r�V���n{q=k�7c�B�\R�!���ZM���'GV��)Q�,&�i)�cǸ�s鳽�禂�f,�C�$�v/�G�8���	��̓���3l�R1��"�+��rC��4��]r��۞�i����b����L�k�Y����J�_a��F��'��K)��.��'���t4!.�
_����ϩ��\�z0�lJ��#�]P���5rC�'����=��u#��l�&:2�0����qx�'lC��2�H�6,h�)�˥��Gdт�3��*���q������:���w�ij?g��z��%��ub����lmo�B�F~��.�a�1��l��h�sn�݄���n����m�"��������!�T�.�_>Y��o�>�
}l���D���l��~9-"����A����XYʙi����P��+�O�@|:������l=����:8T�*o7�z^��a�L�����f���|�ۧqM������ĉ0sa�M
���\�"en�*]4-ٕL��~��!���P�J��ч���Ӵ��T�'�cl~�_j(�dG�;��P�3������e�a|֕�y�P����7Mⰼaӆ ��pG�+L��=ˤ��#����W��=ץ���ٱE:�,�U0y"�P���'����F��S�7 �~S|��2����wvi�l���L'��Ȥ�'B��.�Y��@2F�`2x�6�r�:��Oh���]����[5��+��B&��WQh��Hz�$��X�Ѻ+���\�����$P7����_�w��J��q��.?�����Z%��&����2��̑^�/�$E��R��^��G�Ԣ|U"	�[�*W�q:��Oy�f�ڐ�t�;r_`x�x0\��i���B���]����<`9'�0�ȹJL��s�����K������[�v~��2F�}&$��y���oj_�����h��� ��M �3�2o�7
P�:5���m[�lr/�mϖ~o�p��8���4a��c	iZG��R��V�1�6�'�aḹ���Ȫq�M73�$	U�j���LN[�W&�碳gс��m���a>5sI�Ta� �Xdx��1L����� ��O��te�ԙ_(B>��
A�q,������#�3�Ȧ��.r�b����=���bM.���d*<�=��R2Pe������N���x:�R\?޹���r�ܤC��OF����0k�Bi�sP�{�-�� �g�`���o���%,��O�`�|���.��hF�~*kVt/PV��P1����z7��W�T3lL��{�Қ��b{�g�W9n�0wg6	�&���)u|u�	�A�],��iP#Ǽ��\�!=G=7$�!蠰s���?u�d��a���3RMr)�?�t��t�4��(c�܀/:J�����KS�b���J�FC�!�p��"P�2����e�`r��o��:Y�t��[���T���5�{���rS0E����n�e��-���
Μ�en0�l�O�b �P�>ܖl��p���$�:�zyл�ء���q����ױ����]���z�/z��ק2�"����ZP�ÍlWW�t��3�f?��-ò��Ͱfآ�,�E�F)_V���>u.�~�q�i�� ]�s�Bʀj֕t*������7$�_�Bd@XU�u_�^��d��b@
;w�R~R�W?u�r=��	��n���5��}'rǖ9����Hb��GC]A��V�Ա�A҅Q�Y�[w��OE��8�DJ�Ogq+]4VP�����x�o�:�o��#�OU���\��
A(�d6�ݦ�BҤ\���f�z��#x)�� �Ra@H�R��b��x��ӭێ<u�geˀ6�Bʊyp@�(����h�p����ыzg[Z�-�dg(��q���Ϧ��@T�~rx��qc{:!��K�h�o�!͛���k�iR�2Y�ָ��;[�!vz4�\>"�������])�J�R�y�# ����f¬y���IUv�UY�D�5b��Sit�S4����`
��0[��-ų,N�^�;渳y��PW��H�A��3B���^����v�Y�w�]��?��g�&�2��f��:~ !��y,����Ό���G��`	�"��ݾ���f�V|"�I�����/�H^s;���v�vt�3x��}���ƎH5|BoV����	o��B Qw����?u��r��~�bC:����C=X�ڻ�=��Z�$I�H�w�>����9T�5���S����f�ѓ%����M����c^���6o�������P�է���5�L��2�Ʌ!j4c�5k�cW�d��8�m1�L���V��s��%W���
L�U7�A�i��Q<��6�R`�aʆ�-:��ױ��9��(�Q���[����vtpk�B$Qq�2���*�\�p5Q���#2{de)wG#5
���]1��wL� �
�,"b��,
|����
3 rA��`���H��%K� �+���\�`�����#�p�����M�sa�A�F����z�2���`����S�ynT�L�������l���W�,�ʝ��P��%/I�)/��ï)1L��Z7��(,�Qq��ǰ�y�Zڥҩ{��πpY`���Q��������@��-���gU�l$)&����h�x��!>�V��T�[�Fhs�&��덝<��:�{.�,��n�jk�O�{����o��8�	�Y�k~�e#[���ԉs�Io������%ֺ��K?�dԯGж�z��p�����I�����w��b��%Z�y���j`�6+U��^�r������#�� ?��=(L�����U!�]���!��6W�*&,g"g��zv)�\�b,���'j�d�m;ܛ���f�a� �Y(�	mLd�i�tT�䧯�g���|AV-��Zs3�xF!'�Y"?V/-wM@�jd�Ur2�|�ǟ'��G��;ul�g~��߱K�n N�g4�g'��k��F�?Nt��騼`�o����>�y��d��ģ-'�i��-_%���I���N�q'�b5N��(�ݹ�]@Z�wB��\��jbe�n��d�0(go�j����7}�~���6Qg�6"t'�'�p�r��K���v�70�\�Bo��������w~+QL5��w�B,	4~ ���O`�^i�M��$���AXd0�r�WγДY=����-�����?j���.����Z��H#�E8t,$�R��@u[��_����++#�7$1jpJ��s���F����ڟ�![���P�U��	#�~q��m�Ѥb�F�r9�;;����Վ�R#9�Ϝ�mt$YQj�SK۶B/����069�@7V�q�ڎ���>f�;��@{��f-��bS�2�l@�䚣����K4�Ex����0�p��2�l.����$X���I�o�E��0ƴ��P/Q��7����(Q��(j�}�M<����].6�@UÌ	:F�Gf�;H:'Y��Y���
LgpnͿ5$�/�w/$�
fR+l��lGX������E'x��7�k���ң52�N&!v�>��g2+^�X��ﱢO|
>Y��Y��H���V3��a��_�5iy��� ��>Z�W,�!�+O�� ���J�cU�ai�{�K��;2����1p^�7Ku�H��E;2ke�ԩ����u!��E6��m �0�1��=ZeN]Oka�=s��!F!c�b4y�u�8��u�շ��-X�|i��w���-���9� el�	F�6�bA �.7XtG�BL�]:|r���9����S\���O�JHUcM�x�33xI��c��p��kkb�a��� ��:8�-Ҡ-s�	N�cRv�~Tfu�WN�<�=�J4��~���a#d�9�� h�~B���U�����Ӛ>�W��S>�.߉R7rV����vm�S���NҀsݥ-����HW��NS���޼	��k۹��L�Ju�ZM`<F�^�+@w�>�!��'�E�xkA��t���Fͭ�����;�U�yK
� �_=�'DS�v��~I�g��
U;%}GK�dǅZ�Qq�Ƈo0�ö��Ab�w�� �@��b���$Z`0�8�U�=%�Y��P��� (���||���GN{��)p	1%����`�������4� 5�.j �
u�J�E?�#N����\t]E�����F㸘�ߎ�B��/�hB��x��#	ïEyS��yh>�������$A��Y��Ve#%���U᫫V_�-���S�s�ѣ�.櫀������c�	~����l�J�U��ƳO�X&Hw$��;^�@ނ����Q�/Oj��,GG��?�%S�f��o\J)��ub�!(��B)�r�����~]8F�ߓW�vR\���q\S{agu^�h�`�b�Jy���Td��!�Tҧ-��l9.uv@�<���s�"`��$�:s/�H�0�}
�������L����;�S� ��a��C�N�􏙥�u�S��5�������i����e���c����u�҇�.6`����#����5fL1*���z}�hܺA6�(�B {�%���VbIyȤ��Md��4�
��&{J��b�����R`�'�OG�SUV֛6���e"�N��g}�tY��Ey�]blF+QKt���(���cp������P�ƥ�fz@���%�R��Un���]`+�[:� �z3QU������s�j���OC���
v[\0Y$¹e+�w<���Ð��`]�t.���0��"���8F�H2�9�I?�؟2��g�M���tRk���W��tЖu��}�YZ� ��W~�f�.���A��
��A���ԕ�����Jo�Qh�RKd����!m�B��<l�OR�;(0��E��@*��@���`AV����.)m�A�a�M?!d���/��f/� g��pYr�q|8m�j���d���sk��rJ�P%�兆u����}lW�Jt|>t��A#!h�xD(��U�ed!?�pkF|�&d^��p��0��k��v�q�<v�i��2&�#�F�.���w��ev��ՙZ��[�&vжd�ʍ���$��~�p.罡�Qнl���B�N��y�N{Ջ�V�<{'�>�`���f`�М(�>̲얓��s�H�tV���Dw]%�J��U�f��O�D�:��/hK�ɐCp�;l>��p���� �b��#�ZR=��r�;xs��3c�1�eB��Z��gZP�F��n.d�m�B�Z���i*�'�>A����,��*��I���Y���yt��j!�W�q�[u}n��P���b1�^J�5-���p.\�myP���&�^
�"�7I&Nt���t� �}�G�'t����ےq�R��x�T�m){O��DǙ���ZM��5/���!i��:ǵJG�:	U'��Q����po.5�`kM$�pRX�qqڙH��w��eH^��.b���D>��s�oF/@�)��Q23RLE���V�3�HΗt�������\o�p�Z��#Ш�P�5�7��ޣ�����ҧ�>�  �(��{�P�0��(�D�pg�)L]�< WA�{�R�3���:��S�υ�[����w�f86��G5XYq����K80cgU@Z�{��VD0��i8������i�]}�p�I�����Xj�c��p��N{�F�z�d���ǋ���_U�+���ZU{�b���|~Ɨ�#a��1�������~�/���\��O���j�S8�t`w��C2^{f�A6�ճK�ˣ,�?3c[�]�d��Ъ�}��t��S^
K�Q��|�C��>������-���YT����>L��U�b�X6sy��E!���v�E���7�m�rhx��~:/��c� ���p�u3�n�y�^����o6�v�F�m>A3�ŀ�K��r���ߖ
�zཊ�|>�b���q0E�ռ�/lvo>gR:N>VS���U��e��U֢�P&�Ɋ���_�`�:��\zsk���37"o�bQUu+��� �2�&��B����s4�A(�M�0/|��^�}�k+?7Gۚ�ڃ���H�PY;y-G�S&��2��?�y>�/��*�7��P]!VI��S��U
d��|����OGs�eД�!���.CAF�Ga�F�l������L�a���J�3}���>%��O�s/ܜ�N]D�I�%��x������$�2�Х8lY�$0Z�������M�[: n�[�N��[�k�Nu���������Br�ޣ怨)���i���[�����/��(�����"9�8U�ⶁ�p��ك��� 8�7*p�I��x<��o�gtL�[��̚�Rc��䂙�?}ѫ�ż>�Q�ʊ��!�] ~�wK��2��Ux��|�%QA)G�L*��q��
{R��� �{�Q�5^��]6;G���AZ5��2� �s����'X�6Q��O]�~�h�#n��)�}(�\K7R�;�!:	hyL�	��[$hO�x��^,���E��"��YO���\*���p�`m�S8�VNR�D�gO�D"��_$�.���	�bܙ#(h�)36̱���J5Q�:&��?vQ��I�6
4����5V5���!t.�{e&9˞�Yŷ�*�m��RK�]J��,�������
.|&d_Ƕ�z�*�h�����t����\���+`�6�w)Pa���rE��q��U�D�y�m>|�>�[�Bj����c�h�0M/�Ɂ'�}���\�&�e�yȖ�c�Ӯc"�>(����W�Wj��K�g6v�R��σ��_@�I�N��ؑ�-����(���A69]$966x�v�4�?��複��J�7�gyd��L�F�ĩ!��3���^}̹δ�I���4����'�e(:��� )s'<�YLh^V휾a#��H��y�j�"�v��3ISND� �zIq���v�-��|R��F�C�PN8~���~�|28H�;eB/#s�j�r;���-�:5�#LW�v�H�C�@(�����4,���Et��>o���_nz6m����-�\�Bm&��T�������s������Z,Y�(]�w��P���Z��*�w�L�����%sz�d��,���)�2{C�/�q�]��A���#�_�	E��ur��y�?7�r���o�t����X-c������l+(�(7!~��'���0�5�X�ל0_�V���f16Zlz�Ǜ���;⪈�P
�'%H*���z�۾���eJ}@�� �TM��d�v�x�¯e�vp��!���	]�8��H��̈��m��ؤ�i�m4����x~���q��Ɛ�U�칙��NC�&��ڔ�idAG�9�R�Sɝ���!A����i���"4�I�)�o�oD`�x��t�%��}Q7�V�}��,�Z)]�h��q�c��pZ\�L�u'��z[�A�7���w=v*��m��%b�\�J�^�\�!�kZd���]��!�>z�.������TlH�^�Rc���,�]�j����|����ƣAώ`²'lv�� �08h��
SE�U��*2qV?���Oe4!?�[fj�c�]�7�^�@�-]�I#}m�	�&x�(e��F"p[#鈀�|�w�u��Xb�Q��o:4�U� m��r*�Ҝ�)�U}kGo�&3��9�����-���Z؇t+߯�r�]��sٲ[� �b��tK�-�9H/_��a��7 ��<���'t�f���[I��%nE����䪄ήS��kF���
�[8]�eX�d���kw��1��HDh3�J�^׈����nX��`�<�x��T�Ʈ�����a�ȝ���:ݕ��̿,�!��)��\YiecȜ�>͈�,�M�h��8��6X�'G2��t�^���fs�u��,6���J?<��y��)��&�GJ�G�*nBD�k��Vk���L&xU�1�[T��I�ꮤd+��/��\(�k�E%ڜ�u��K��a��7�x!�� �yj�8���f�a�'�*�\k�ڧ������d�Sǭ�%��l���G�q��e+�
�\��ucWa�=� � �tO��pi��jY��e��Jq�y��,�(/��i�t� �ס! ϵS<��}B��4�g�Y@�z���|;���q�&We/89��}c!��g9{�PF�$zNFT	PwԄ��go`�5��-�jZ/�!��!m^$�!���	fX�SPlx]Ԑɺ��-�3��4�-6�����+�8��Ɂ��N�̐'W�x���	`U��H�D���Q:�*�~_;�C��JK��m�|v5u�F�Z�C���E��t(S����4�>�UZ�u6����2{����ڒ�����n��"6D�R����,f�cA�"a"Y~� V�	S��63��o�8�*��-z3-�7z"1�� .��+*����V���s�4���1?sƎ�;N�02jF���I���ܭ��ѱ�"u��p��(G�``�p�uN:�jU���^yXX��5(贎a���(֎��U���S�[��;.����*-ZНV���/����g)yi����H�M$���x���".b"B����t��[϶&���NrL\�};6��7�N2�n��.��K��.�"��qv J�����^˘�&��зMR���(�GqY%��I	1��>��ǧ�+�sX8�]_��� �+Itajg+dFv�SH�͏z�g��"��>��@ȃ����b�b�����tA�If�d ���<��F���h��]P�yi0�g�u���\QV
����̘%$�����8	��:c����=��,}�j��F<�B���	�y��u����|J)<���"��s���LUb�i��Yj�(��*�8J�z�	�l+ �w����ePk$���(��`�E37�G�|�~��D(��X�`VxUG��W۹Z�������N:�&��ֳ�&������³����I������.��,5�i�DS1����̌7z�۬�@�~�se�p�T�DRr�1^��"S68+�lyڲlĔ֚YQ �R3�e@P�,+��H��W����}�S��X�@�L���\�����9���G�HT%���֍���:r�YiG�7����ca!y�=G�^��Z�_c�C�����95�������Tuj���ԗ8��!��`��uDx�b��4�O���CNJM��L�/� ��l��Iø�������zj�߁�e����>��{�4L��eѣ���"+�H�������I�)��̏�VI3���q����3���bm�H�W�Օ��\=0�*ˊ�YG �0�i��P�b��?�#$��K�ѽY�.�c`na�/2a�y�[<��
�B-�F��0|��������ĩ�
sj:/Bc����h�I�9!V��B��ke�P�A��{�Y��;{rj�RN���Ay�qOu_�ӹs�������O��]ل�ħb�0��s�H�r�c)j�'��C�R�]�Lv�-t�4C\���F��ipQ ZG�	_������4Ca Yb��h���-a>9���bJдpH�7�c���$B�]v <��E<u^Q�����j�ah���B=�-M�3��\�r�Dw)��'�ډn�.�8�����b�D����e��D�'P�@��0�[ߖ͒}dc�b��	Fz}L�}f���.�]��0�RV$�mاԡi�)1�+vg����ޡM�ܺa� A*e�Yp�^�
W�-Jg�^0׉��)l�=jZ��̰�f�'�h?��.�*�'�����j8�z*��W"f6���GLh����ۨ��$���n��,`r����$�$a��d"�~ͼ9;�����>8�n��߀����(փoE]LsJB5��)�"�TF�;{
@�t�+��3�r�ܘ��.Ȝ�/	UH��|��d�eb��-RX#��e�Ecz�WSɣx��)�J��x���#B]p��"H��t��]a����X�]��t�ۼ���-�o���}+�@�2\��R�?*hd�D��L��7����$��ݨ��a�Tw�DR,�>D$����;<���;5��B0����YMm�y,!�q�w�No�wc�����i�l��[�'l	r.�G�N���Hut�<1�ຬ�4�|�#�TvEɰ7n�E�H�?�n�������@&�B��؉3:����&:�1E�π���b h�/��'k~�|� �(C���O7{߉���B(hU�{Z ��m/�`ΠtZ�=�� U==c��1t��ɼ�J�֦)	uF��f�߹�����!�+�#%�L}�;a�<h�7q��:�r�b�N��д�j�C�:�\)w֍1M6���i��|��=o�O��xx�E� 9�T��fu��R9���<\�����ߘ��&��\�zo;Z��6;�����l0�4qjI��e�]v�f>An@�'
��W��*��U��OL�} l�-uFV:��̑7���T�7�"nn;K�y���T�k��)άb7�N7�l���ň?ۣ��%b�"�R���DQ��kBk
5q5)���]�y�ݖz��0�j��b���9�q��R��w�v(�@��qP�V���Ȫ��Ge~dr}�ʮ����ImI>��N��/�BQg�s�6�\N��`�_q�"d�8x���*�f���{�q�:MEےՇ���32R��9�L�²�Y ��=��j��×����P���(�����=�lpթ�\_����+�rGV����{w�fUY��]2��_�����p��6�Ҧ�V��*3�m���R�J���KR N��Zx7p0Ηna�i�����!B�\��te }��߆7����̢����Bf.�J��S���39%g�E�T�T� ���opJ�Y+y�:_d��>)�n�b��@�����\|����|��'^-������~�D�?�h�h��MMOo7,��$�m����Jo��o�,2� ����ZE���=�7��ۋ$TO��Z����ij����_)��.
.�0�IhH�b���zü������h���8��7=�{W�Fi�c�*�Y���؇�����V�gX!�Pe{OE���`��0�Ӏ# L�yy�VDќ�	�lO/}2�̫�ֵ4q���9�����oZ����2�h�	É�ߗN6v����P��X�b,w���<~n���X��C^���XE�K���\��x����\Ũis�)|P>�{�a�wCo~��'(��+����H���O�tbˮ"�����w�Υ����ɀ���w���PC.ٶ��IԊ��w���h�_����܍f��<�n�.���c�}�(m}���v�k������"k��1I3����₊8��C&���[�W��O@�@hJ��k�.v��,�Hm��3��l�yS���'3l@-ɯX�����4�uN��6ò;�� ���;{*�`)�X��*=s��&3���ǘ�ޓ�*y�l	�-��t�<yu��š���o�W�(-�QC��?�;0�Od5� �zC1n�U��kǰ��|��U67�a*��������T)���n5�������E��b:'hn��A_%�N�Ԛ�.�w���y���%�[YxAk�nzjźy��4D����(̀�W4��M��C��}�OL�z|�9D�q��&H��DE���?,1➰�s&]���w�z�+!s���*�� vx�q�($��hK8�~A���ע����2���]] E-�ͪb�nY�8�,����,�,Bλv�O����c��\����7���Y�n�Z9��:�(t����a-$�	�zO�B���G���(�ѡ���$(4��y�}=ț!v�����p�N���1���RN��?F�W�w�k�&�3���]�4V����((��o���2��[���y��_5 �Rp�<��6�a��NҞ��}V�(��h�,�#$]��A���
���G����j}2��Du�f�������P��e6Xϴ��s�;��:��n\+�UO�QU�)�#��8�u7�� do9Z�`��(Ⱦ�iYPP�9m xC�	��s�  ��d+��by�G��-92-mYIE;Z`�A�߆�G��G\�)%Zg��#C?HA����:��e���	I^{����%�l�m��c���C�b7�n�Q9jK��h�Mt�������G��qI���K�qw�E�0���;p_�ӧ�;8ͥD��.c��t�A�S�����ᙑO�g��y�Ք'a$d��-�s��wm�����^�C�$�ڕK��p��V����_]\���"D�m%$o}��)��9��[�/X��N����#��˓I��r�
�&ׇY��N�� qRڔ,�:��;�" ��J��W�W�i����iA�3��.�I�7�N�/��=?2k�"\���7⼞ �߳�6����bSO�����;�t��U�|J;Y�����o��P��T8^���&���9�"���������G�̞m��n����2��G&B�h��R
�#������tp��
w4T�H����fմ�+H�1=?0V9*wF޿�=��1���ڴk�a�s��e(V/��h�?@}�R���� ��Hi�ẙ�=����_��;�ڞ<��Wr�lA���Ok �Ö�K���sj-�+��l�X��`/��{`��%g3kU���#�T�������?i}����doMJ\�*G��Fb3�]�̢/i��&�f�<x3�����F��%v�9���5�<�](z��_�����D2X����ķ��u#9Sls���H���_�ppJvS�q0�\o�S�?��.�7�LXe�A�N)�c��Ҏ{H��0ɚ�VQԞi�-׻�&�I"�r5��ٍ�kr;7p�QM$��<�yϤ�	h�v-�m3�YL��>p��҃��a���4��73���'W���O�$���x�7-Hl�4��"�v5[n���d�!TZ��{1f}��a�
.p��y�T12hݛ�dq��&�����]�_���Q4�j)/�ڱ�F��{�1��1�V+����_�]��7�4y��glh��d6i"J�a�"����.S�������8?�m�������ɝ�0Ǵ���K�X�!T6zMs	�����b�K��.|B߷���"Z���ؒ��� +��Nz����F�5��b\dVu>���%�$���s@v)L�ʺEC�Af�1�"R|gɸD`C�� {��Q����i�T6�<6�1K�̇����C�l�3�#6��
E5:�Ȇ�p�#�7�"��xT* l5B���͆��O-:Z���ujSN�d�<xl������^Vf���<ҍ���(�5Ю��^^���
����5g��&Ig�/uU���������|�����=2 3δ���pX�R~G�9��Ǒ�r��|��v����i��H� ��ߗ����������U�3{5�L���uH���R,]ɋ�ظ�ͤ.�������p�9Ε��
��x���rZ�A�a�;mmun��<%^a�S젗��B����k乐��P[۝Y��!�������*�T^=�'�4	��Y�g<j�����t�~k��~[FR�M���|�R�e�H������y�Ũ*�
�(�8EV�	P����:^Ia+u2kF���_,i^��2;�j��w`�s��'D��K]���{O�5JCf�~����$��+����,�K�~V�a�&tz�&b~��JŀwR���>iP���`�K��MF���k����&	0�=�*U'��M�Ϻw9���hP@�.�����"_Rl�E�-#�>�Y���P�}Y��?i��9=�U��RP<��no�J�A"�����;�BبGL����Y�ED����+mjP�O�������Z�L��}��M�n���,WD;S��ۮ��8j�d�,V����A��BJ�]sђ`�?Ba�ժ2�pN�꾻_���7K$�_T��R��3e:e��K>Z���vS�ú\�H@k>0�w���Bqsl�]��ol���UEΜ�w]x�x���	����T��#WE�n)ų*��G�� G���ph�!c���T���J��I��\���.s���Y�.�$��F�D�֐P����J��#��VE$��I�o�k�i��ZD�s������`����״�WJ�3����N�|>�;��11��_�G����:��,d+�4�	<���k�B��D/���)��k���'DU�&�E|xyn�2�=��x\}����-)+�uGu���Du�� {Aҍx.��m=�"�T�N�+p�gԃa�߶z�m�cfQ�ݳ�}�nD���j2a=5m~ ��_���n`�=��bp{�n���!�������� �@��P7���;����DG���0ظ��2�'��-�f-�o�T�Z�9�++�x�I�/�����5s��\&0�/z
S{G�q�,���v�es�l���^:ڔ@p;c@2.��"�g�v7��h+~o���'K/d%-�����C��~��V�K�z|�&�ϸ/�M��F�䡝�.+���;Ma��v}�#�
��V���(P����bd//+�6��=����e��D]=�$����?�l�-S�(��f�I�n���nC���t&�]�E]���)�G�>�+*��ui+م��)�?b��$3d�����%�����k���e��R�2c^��2��Z�1��v�OzV�E�4n4��Y%9j��]�UݞG~<;�y^�D,�#+�S4�/�Ӕ"���E;�$����aK�CQ%�P�����9�b���d��zr)�y)x�Ъ&fN�W�T�	��lN�}��=R ��`俘�\�!�aKm����u3O���Ό�Ӕ����1��A�|o��t����4�Y��1�ʾs��k�n*.	f�lKe�[��*T>����<B�&Ya@\�fAL���F�m����P%6
�DH�R�E��Tӵ�3*u�z]�̂zv^�uD��r~�q$����I�4�y��N�Y���Vdf� �l����P��,�'��-ex�Cf���K��Y�������w�~Bz�9o�vm2����0/b�?�n�%nĠ��c��1�FĮ,�]�U�N�P6�z|܁˹���h�zs��S�(����h>�dxkpΪ���<�4{D����I�ÑͮC�R��̮���,��������r�D�w�����@ ���v�l�c�#.1�S����ߵ�0��e����O��h������W��A���N����O��BzZW���؍�=jPf �xcdf�^�qw|��=�r��7!X������߁T��� ������& 8H��!]����>�n��ekx�'�t���U�i���_<&�<Ͽ?Z�;�����L+��_�(�Ō��>����$�i1~���~���' 0<ۋ1��6M�V�/�L�"���zP��Y�b�����(�X�����'�z����%�Ѭ��Dy��oX��|m�ԇU�ߠ ܬ =k�Ud	\��� *�奌*(4�7o��:�s?����Z����o�Z���h������>c?'q7���%��;҅�N�R���>�&���*���'�s���K���.#0�;Ј$���[T8�����;��B�7�����:aPZexe%�L��P���?�o�M{���6���d��e�.VV�va�����F�V�/4`��/'����K��~@��
�=aɀ'�"�E��m����()�B%$0E�~��^|D ���_�����z�!��2l���J��s����O��`���h���Z��IORN��DdҞg�BU� p�iT!l[hՑV���sɪ�����+���ｫ��4]_&l�>XpRx��m��.RL�/Eo�_�<wƙ]p��M�,|��w�0�4 b8�-@�(yq+�ӥ�RF6�O�=0#�1�~��i]�߯�%�pæp��t���Do�7��g
="e�,.�`����idco6
-*�Ze� ��C��HV��VB�*j����)�X!9��CU}��Y���kZ|f&�r_ټ4�;�$#�H�	�t�u���f����X,��J%j/Jq}u�V�/��N���h��v����t�}�{I`��K��.Q͓T�J����c<��k��T��^e����������)E�Mj{.�S��|�(��h���i�o}�}.���m2
	UjfBZf�`��c�5�_؝��^��'{Sc������w24�O�s�V'6$YW�D�$V�E���w�� ����(�j�	��^�(
UU�>�xa��NC����p=Y#�ފ��Ju�j�(�cx9� fս�,y?L�r��8�u���S�yN���5dU.V`E��RX�xu�_c�|�B	ϳ���j����'�4 �R�W�ٯ�\�d�n�3�K�w�bS��S�/X�Ek˦T��)*A�[�,��ty�R���S���0UNv��i�U ��ocV�'�G-��}�R��]�k�F(QuH�Cx�滿,ch~Bv���#�L�V��^�czɬ����=C(�jg-�����$3��3�	����lL����H�:�r���u-Hn�S��MMK�*��~���v�G�G���n�p��q��޼����y�_�I��#���rX���f81ן=�/�[�Te��)[��)��{'�P����J��q�1�
l.��%�覂;Q�z�O�O���W���q��Tm�`�.����
�a��շ�|���n�0�2�#���^-uI�Q�����Ā�Mz9���[\�}o^ݨ	�c��ϖ���
1�hl�� �����;v��w#��It�3I��Xb��E�� fn=
��D
�H+�B��O)�K�"r�)���NV7+,;~�G�n_�G��Ӌv�"K�9��r,]�xĒޚ��Al�02�OJ���Vd`����7��=�EfI��6Uw,F�.�x��T�����G��=|�Q�����L�����8� �RL�:�{�C���3�@^�=������ ���[��0�(9���8Q9Z��s�]R���N�C֓;{+2l����_�ܤ|�F����)��b(�D�n4}��/X�w�.k����ɩ.�*���	�EX��o���O��"�w�>���:�E�O�@��M���F a������@�Y���N��	*�j���_z�إm咇n�ݺQ�:�G����.l��T�7۷#�g�9)�[�a�A���&��̷D. >�YM����'�ܼ��w1Yb����8S�.~m���v:���K��Z�f�
;���F\eE�|������ �(���������w&�u 6�_V+_���2�YB��y��[�Wt���d�ɬ]$�K�4�D��/�R�� d��B��fN����q��0��#�6~��3{U"����%�y̷DO�JR�9���#7�e�d
��7!V�!�<~+���/�Ѓ�k6�X&Ky�n �k��RB��0�!�;6k�~Yx[�~�P�T����`Ym[��0z%"y�����*��D瘙QN0�u�E�֍��U�+4��;���n����Z�p>z��PL�ئ�^����U�l"���?���iSO|�5��\�m�P����Ng��M4�A�
b�-�V��2�=�����@��l,�[�K���#�����<`�8_(F�_$nW,J�ء�H��ay��`rC-�I��6�#�SN�@W�0,�����d��V����\�愾�9�k���d©ֻ�C��m!ؠ}���ɘ��S�:�8h7͊����9��{0�.�6�ˈ��1l�|�����ΐ�j����������H&�dN�e� {��	:�7�E,����M	ީg��D�W� ����!�h��>'�3}� �s�̍�'�1�͔V�^�
N3��Id���nٟ]�fD� :�9҈�C��r.J�����_A�1�����'��M}����8�]����q������l]�/�!��$!aN�n��2��׸/$�l�͍+����j �2�+���Ld����_v+R�����4�&�Y��]\��9��7b�Q���jI�l��͟{ ����8�⩈o��Ln�¡$tS�G�Cik~��"D�r� l��A��'U����4�?|�p~M��f|���/)����E`r$�\�|�ݑ�Ʃ"_MII�WzJo�KZ�?���l�z��[���+����h5�X$�dOy�W/B!'��Iڷ��D�Jtte���|�z��HS+(��]�w+�9���=�8/����^��$�r����t$,���(G�v"�?|{2�=F>�џ�8��#tˑ\t�m�j@T���Y��V�;2���Ui��Ct��!���N��bt)�В*MX[д�HR���������C�:��jV�彛n�4�NO=ę�ĿG��r�+
i����˄1��~a~���}}^������{�5�H�ثXh�O��
��̴̩{i���'��:���9���[�>�=�0
����Z��OR�mj���!𲃒]�&�
� �W�*��ϼ���Ʀ�؀!r:�Vq��R����5���0.��ɤ��Xg)V3%�"N5�����'U�d��� Q�Tb�]T���C�?u���%3�י��*o��L����ڗڏ�=r�$��;Pd�B1��
���,���~�k�u�Ӝ?.�b5pVK�R ��`��}��<�ބ`�[�j�=CW�W�ǂǷ��������6��{G��nd�=��`U��0� �j��˕F�%}��7�V�S�x$�JY��񅆣lW���c���`�.�k��'�%��PF���������x�a��>���ڳ�@h[�&�T����]h4]���:��M2�NT Aw�~��� x��0[ݛI�j#�N@^#o��/�e��yv)�z�&eGR���2茲zq����=l�b^oV�#�t�y;��h�JzH�xء0���\f�f�TNge�2ъ��D`޷�N-���'�/r��n�}�pِ��Q��{� %9��`������Pq�|�N5нq7�)ټH�)�
����D����nF�p��'+��汨Ĵ]�i���ХHKwu,��z�!gC|��������U1� V�u��fk��QX��8�~����W���E�ف7�̊S�g,�$�*R�S��7& x�@�c�>��~��r=�	qF����}��Z4q�-U�Jꃻ%NC��#}�f�D�G�DMc�%�=���Zd�߮��}�?A�E���Xx:��}�f��5p�m�N����\O|�4��2M�d��+(&���R�@б}c�)i�P*C,�8J�ndt\	Xǻ���c k����Yģ�u�^ѫ� �Nm0�U!�*�${�D����I���snXh���&�Q&A}�� ����6M�'gR�s�߳�y�]��kʎ5s!�q[��"a�x�XF�$�y�r����5B.t��������L���2�%�k���V���`A��cAP�>q�.Cw��ϛq�hN�
 �؜������^A�Ƙu�:�Ey�!q3;���A����2=^X��[�s_������[YTD�4�Q;�+4�\��˒���ش��g��ӽ2��v�	��k-\�	r]YKt�.�wx?��>l�����֘dqch�"�^���%"EBo�lsf�*�Tgr�񕝱g]Ö*��6�u�X�Uo��~ #�O�����KY-�z	�?S�ϊԗ{&.}���iK�t�	irO+��e���Yf2�[���.R��U���R��0�_�R��S�������{'-�Q�{�ƤD�fx& ���pf)r����60�[}��B0u� V����/�d��s������Dh��o�e8�0�T*J�#�b���r>:�o6�i��]?E�4��?rP�`/,ߥ����\zLU��p��~�Ƨʄ��u���|�	z�Nb��h#�Lt��}
i��5�6A��c�\���p�t��HW�ӕX�R)��#��8�0�P�Ҭ�(8���GC�38�m����k��{���R�pA\�Wa�Xg��}�bW�W+g��S[W0��	�3�k�u;�f��h�%#�פ�r��P�tE���܉k��T�e��%'-���N�]Ǔ9ü<:ac�/���~�����y�~}~�F���C�
��d�G7��y��p��js��&K�zV�[�ͻ�!\�U�ťe"_��̄�lb��{ ��h��9���t���$��`�^�eե{ڞ\?��yTG�'�~�>Ē�X �����W!�8"��ߧ�q��с�;���=+����Q4>��dՋ�G�����޳J^%R�4���+��r�q�}B��oN  ���ք++��
�/���n~F������3��/H^���{��'�B�=	+�׾7"T�<qwڀ��4�T&p<y9��ٍ��
� d�b ��J�d*Tﹱ{+�ś/~���_
�)���`m!I<��m	���M)p��G�a�y��aE$��"��"U:���@����Z�=4���&�i�'q�\����E��*7�m1l|�V����^��]����o�§`.�:�<�BE�������3/_����mq�i��iӘLU
����\�LB�;p��Հ.B`�y�U��%W^���;��fA-:J��R�Z���w<L0��"lN���@c���*ia�=�6p47R2(���q㋏����I$�,�t��B�p�wd%�v��cO?�u,k�O��A��Q��&ko��˿�.d���]d#�Z��c	&L{�}����rˎ��ݭ�6�?ᾩ6C����Hg"�b
'|Ab�v�nLIy����ף.?��z5�l�M(b��=�R��o�rȸs�~x��Ly�ޗ���	���*����l��$�&��W��G9�<��,$����6���\2��S�{Iò���]�f�U��$�r�:>�.��IJ ������׳�����5�Fs�8Y8|I>{P�jǯ����5�9�Ss�J�e2jE\�k���w�G���]�J ��t}�T��y�z�?�l�	�	� I�y�=��E嗯X�]bm}�'���i}��,�$���h�\�&{ ��S�=��~�i���+�߯^�t�1��T��k�ě��W��'��]Q{��d藙aз,��0Z�(2���=P���T�I�B� �Fb�NW�^�/�<j��M�W��3��NSj_�)	�E�vUV�Y����t��+�#�uD�N��;��{��yH,2$s=�`c)���R�s���p/>/�}6�bnq��2���̯#c����}/ץz���Ԥ��#�RSċj�jU$�3v���9���C��9m$�l��0��F&���8���0�ț>�;���朳_���φ��gfƋ.�Я�cn�W
��-��^7��� �=�C������7-)<���m|E�DaX�P�Q�Tb ��N��ϳCm{���ꂲy�7��HQaIMD>l�e.�G��,��w�u��y����0��]�
�Y=ngo+E��xԍ%X\��}5�4X��*��C������u�m��y�Fn�-��=X�����BD��9�n����tڳ~�Z�nFJ�r#�s�����-;����`�v���<��n�/�(�����"A���3�:߮-li�ق�������n�;
�g��E*0�/�ps��R9�%�DfuyI��F�ǩ[���K�_��)��R�)��q��U�)k�тHE`<�[D�	���'Z�b����46J���c�C�}?X ��G���G����	ɍ��|�trp�Ê��Ζ�ῑ�{� �e�$����V7�?[�8� R��On�T���0�T�(����#a{�L�����Ot�Xx��8�zH{��b�=��c�w�d�9��]�ׁj�������-�.���~�i�� ����QO�'gsV":��Se��F�~����#���!Oq���I�v�q�zO�^D�8�臘�la�o�]J|����������R�[�P_u-�\��q��?�k�8�r#�(Dc�l׺�k�I�/��h����x&���s[>q��Eb�w$]X�\��ރ@�1��xϪ��R��ƀ�3��h.Du�g�����ܙp�,���s+�N�mPW}a�����J��<
O %�i���kw� �*�¾���a��6�A3���w�冣YT|��W����r9�� �����r�0#�sC4r>�&5�F��m���gtQ��c�	�.��l�0�c8N��g�2�yi�w�
mt%ځ�K|�qy-0�e!^(Ij�\KGX��O�*�y���u�����7x`C~�S���#sa��\G���%)��C�6�F�.�VeZX�Wh�:P&��E��׳�1GAd5�T���z3N(��D��,!�C۳b��E�KrW��TI�{z����^���� ʎ��d���w���$W�B�1H�O�M!�<'ö���丹�Η��ytaQ"�d���Z�y]�yG�$x����x6�r�#e;S8t��3�L��sE�!o�m]񢝅�16XD ����V4z9(�T`zI����0�$�jS�q�Sp�S���9�/�@���D���_�h���4``Z�l�1���ǟ˩��E�yD����o���A�g��l��Q^��?�FbF)<���p@3N���dY5k�����M����B�o)0X"Z������mi��*&�zFD����/���z�I��7�X��6�h.��=Ո6c���q��G�E1�RƢ�-��O����l���|�jJ��t��~ᡈ��wɡR��Gx!�3캪x�яlh��
vLf�7(K�)�~����g��"h�9)Mټ�*�/�,B�aA��pM*M|	�C�i��z���z{�'W5�z���}@�z5�:�p:�f�\�[������$sHvg��Ul��v����%~\3E�'n��a�C��1�L�U���t�d��T�����M�\��wt�:{��`ѯի('\�dX��W���40�r���j�����#�q�����1#:`��m:����\��}�Ւ�̤l;��y�Ik����rM��#��yS�d�)���i�#\2�;�a�h�-H�(�̞Q�@pQ�͔��Ѿ@Mh4���k�p����O���ǩ�T׎�,�����ο�yf�5�<!��J��-]�VzW�M������\��{K�%g�$+Zv�U���oa�A$�2g����J��3�|9'!�%�|t>��]A!)�Tt��D��w��d��m�(���S���KK2�)M�\5³��|8P>k�:ꡡT2,͗Z����8&U
��gGO����d/30����cQ�n{�q���um�H�
=۬����T���ov�	%�ǔ��:��Io�|���#�3�kG�Z2���K�{>~��nO��]�'z���m.�d_%���F�Ej+����a�Y[�\�$@	���y��Ak�s�.�ZЯu��;����x�OK$�o��z���9����x��I������ �� 9q��D#�p���]�!ojtl֤��v"g��M|i���X�ﵚ����{Ieg�Vz�p�.��t���l2�&ȕ�q؁ɲ�D	KN��O�n�(�a��%��Y�����
�KlB?���{�Ln7�d����=�%���Ȼ��l�p����`:��rEl���F:�
Om�T.�#k +#|gט([$�̞`��]#�(�O%�A9`7����N'|�rp����(%@��/Hl�{��Z�
�p�4��,g`��������T�J�o]L��p;��;�s,fҿ�*���З!k�,cI;�5
78��;U����x��5�Q?Q��QM��s	^^�h��b��s:#���Лt���n�g��Uk�����V�N_�WČw�[v��ZB]D��d��X����$�-���|��>���9ȍ�Y��ҽ���m����X�y��һ�Ft��)���&h����#N�2;���E$i��$ ,%dA>�)A��; ���=:C��`��W��eZq�咃Q\�L� yy@�� \L�F[��(N6�PF�(S�*��s}��_d���P�e��oR�b�}:��K,��G'�|�!Ԣ���g�������G��a*w��%�R��~�� N���:FJ���0���,�v��$�2��b�d��տ����M�07td�	44��U*rL<P��O��c��5��F���G�7&�Ҡjk*������衡��[�V76y��'4��Lr>��4�#���E>��2�H��>�3o�P��&�)H�!������{���F�J��d��4�a�Ď!\H8`�aGn
�
��V���h<�8���m�UE��n�ro���f��^�B��Hs��n�m򆑽H�;A�Ts���Nm�R�Sb"i�#�h�R2��L��x�=<9�_A�cB9�x��`��_7>_�\�J��2a�[�25�w����9�o�㢨�(�_�a3|Wh���VN������
��  �Π:�g0���0����V��fK�b�W��W�9(Ugk�
c�S賜,H�{@̽����9~�@z^���e^]!�luu�#��I�x����-Et(��:��%e���YҔ��a�lJ��������h��`����5�4o����S��������=��F�dV܊4���{�<�|�z\B���#�W�jWD].��}&��,�0-�;�)�%m2l�t^�}��4b�٨C�V@���YtۏE'�X�(Kg�hHS���L����?�;R麤*x���~��o��}��2a<�W 2'�)�4��{�O�+OJ"���NI-�TTG� �>��z��J[�`����[Ye8E�P�3#YV�RX���"l�56&�d��U/�)EXy���� ����R\��$E��}"6>�X�Py�Iy ��췞U�L*49ˏXQ�اzv��[��4	�no2�C;��]/�X1E+��S�s���ŽM/v�ۄ%8��+-�p��D�o���k��3���ڡb�M	��Ņ���'b#��8�n7�5]	�3�U� ui6[nf&;(�;h"&��H��M#��A�����p�d����~!7�9��*�=rlc��݂�G��WmO8���.6��s�*
�*�ѩ�,Z�3`We�Җ2>��F��<�H�Z�>JL�k��mk��/��C6��X�j�K�S��ѧ��|.(gPj��.]�[s-�.�g����b�B�kV�jp�O����4>CB�f�g�[�N�Ri���R�߇ڻ���O�B�~Ƶ��O�C�ՁфI>���a�E�i����V�*�ķ6��Ż�3�n���˲mKpW����Y�9�))xj�2@�	 ڼ�a�rS���Z)�������{�i�fA��'G,w:Uޗ� �������3,#�L1�	��o8�1�W��w(���ѫj���13�4��,�鮗.��L4y�;$�JOԃ?Lߵ���=��o>�M9�^��.>�<3����|Z����Ƽ~�N�"���,��(b��8�'ɔ ].��P�o�i廤���J4:`�q~����7�|2���::��Q�*��\�1\Q��Y�uOH q���r�>���M�/Z��ٗ��).�����,>~s�a!m��N�-��`�n]x#�"[]��_�g�ԵR<x�ӏ/k�J�:EΒ-u�iol>�	���1J��?�83$�^!׷�h�F��b鉔��؛���S��12���]y{���#u��N��큮RL�,?oZ�?vg��^�\y�| 
]�=:�:_���{���4K����e\.>#il�^�>;$�Z��܌�6�@�
C�n�!�.~Ew=���^Z_�9�F�p(���-�{_���\��%�cW�n��=$�8%@V���F^���_$|m��1��g�ٓr�\�[5�LpF���
���h��{+��'�xk�#q���s��Y׉�-/��k�
;4D���M�jB`y�F�/^߄]1GMN�I_�Q�Z��+��?>]ϨA\���[].��y:瘜�� ֯/c2��)	*���K����0J%(�6R��&�" �w�V^�Ub1Cf��=9�M��9��A����m�J��Y
@/��ҝ����g���zm�[6Ɠ$��}D;ܯ�~Nl���&� �38�x��r�e�qf��A-}bĨ�P���'	�J���ۂ��8Aa�#| �,�:ϳ=�����j�Y����3��@Rv���RbRk��#��!HB&�A޺�A���Ԋ��%!�r����3���Ʊ"."���Pj����?�'U���4ܻ�㋪u�-~���[������R,-��X�U@U��4��5_�dv�0~��!��ǒ�%rOD����Q��I���|���)��4fxF��w�s��]�/���D�2���[9��ciA��#���C�N�+��e/z�^���� ����~��f敕�c�Yp+�,ʐ��@81��w�h?
iBIޯa�Q��;Tk�Yt2*�Q3�B�&zJ��m$
?�j��iX�.F�a^�e���Üƀ�~�$.l����;'Ѥ��_�7��ŷh-�^��[��oZH��k����heb�)Ta�V��c�(Ǥm���w��5�[a���N�.T+v�x�;6}n8���^�h��s4�FP;� �E��W=�8���
9yYT,��@L��?�ু�Psr�4��$Yk`��ԟz�&�P��UJ}�;pӸ�����,&�9 ��p���Mt�g�6jG�w��x�E� OX�H ֔Mmc7�W5�*��-4� ��Q� �\c�h®����_��	�am~c��n1RD�P�����bJ�E��(0�,�аy)b�`� '%_��2��yD�(9�������0��]j���ltp���z�5+�{�\\\-@��~�Q�{8�j�_��7���d���l�د�0� �L>I%��b,r�su�@����zy���J�,e	=,��t�0��jY���N?ѳ�X�f�9S#1Xk��$u�f���ڧu��7��_��B���Hg-`i��s��9�M15m�"��{,�a���$	�|W�Nn7���.f^�tt7ɕ9�o�c��%K�拈v?"kA�v�)em�bQdy#I�o����s��>��p�%�XJ������F���ӾT��ANǛ)�$��l&*{�Ҝ��U�3Ӈ�خXi�>���B��&�Zp]�e���T����z��5���!>VIȵ�K q͂��B�v�2Sy%iL�!��+��Z�����������+"����O�mȝ��J��br~g���ۊ��ٙ3�:���ؓ���9�q0�_q�b�K�P�ɘPE�A�ڗ�g�~e�sA�_^+ s��C�l:l���TD{�`�VO3�"��sy���`��Q�v#�Y8�rye!�-��Q�;�ޟS�O�5�`ڬH�;�^���^�]�g�]�b�9�]y�D���"}�Yͯ���˔�.EPOt�$��H�H��:��Ǵ��@�[I ;�;�D�6����{D�������@����Si+�_D���"�z���6̦+y�x�s ��7|��@�!LPE�0?;mN]SW����6\)�xd���um�N�v4cw�O�Z���nc���m���$*�]ux�!L�0�[A�/��o�-e�yy��yq�z����[@���"O|&�_8T�-M&k��C@{�������y�m��� l�pZ5��B�D
a*0��H�Q�ާ�2���}B�A������t6r��~�3|����g����c�x��S�I~�=j�J�G���t�-o]�Y?'.
؋����i�kj�	���h�3U:IBɼz�n�6W��3�c+��e��~⁝�{�l�h���)�dvoڒ�Gѭ��	w��q(~���(�g�5�R�H���;�����y��F	P��i��q���\^o A�s�Th=��R�}�á:�� ���uƾE�ʖVS}:��ۻ̓A���VX����%r���S ��;H(s��O�_��Uǌ��7>o�X�mZy��`��
C�ۣ��GS����#��B� 6��H�[�[ss�����.�D#��<�NI��'b��aa�g ��5�S��lX�8	��yx$f^^�4������!bC�Q�];g9�e����5�X������O��}��žW�6�����~��kJ�\KH��Cx-����'���G�A���.��}�e1+wg�w��������uW�:u&�;hY2�E�FڤG��
�ss�'B!G4;�.j�䓫�(����@���qO�D�|�8��^5�y6J�c$�qH�M5Fv(	Ⱳ��67B�jŅ*��Җ]�D'�i�a�,EN��}��]��!U��w���B�"�X7dW�Ќ���J�-@oO(�j�x���$-.��9g��@���%Gb}�3J����;|=粊��Q�;�����r�/K���m�����XQ����~���Pv�U\�Y)&��6��Js롿�|��~a��Ww��<��y܄M�')%&M�D�M.W�^�2�� ��������F��v{G9�s���/��)��{c�M�w@�I>F��������[���>����\�C��$&�h����H�-�:!ǣ��_,z�X#�n�
PH9�jrC��B\� _�L��a1��h!?�� �>n[�H� 	�z��/C�$�����P�nF����c��Ddg��9٬c���(	���ł���c#s8>�ء�h�`�f L�f���oy�P�o"���F�����@!u�K>Ya#MO�'�W;`�=�;y�di� �l�&O��z�^��6�iN��2��>�w�~��<<bw6����&!��^Yj�MV;�:<?	^ν� ��'h��sI���8q�F��;J����.����G���`Wb<O��J���o��CVy��O2Q4-�v�)%<�*���~� (G��cuJ��p�?�ҁ껰ܛՂ�v�A(-�|��+��$L�'���a8~�3Md�|}�;砗�൭u����F�O�n��ʂ�:����U�R{�Ba����L�V�巕:����đt?���.��U����3PR�T4����&EB~�Yb�?��'�����9� �a��n`QA��qrG�t�jOW�h/�n�6sɵ@a"lx���H���dEg������U|���?׋����.7㹚�?�m{��3}O�t4P_3О��'�/�x�b��e�9��G�9�(Bk���%��
0@���@�%��/B�)9�I���
@O�h�5�p�+b�x��څׅ��Q�R:P�&�`�����:s��rY��?z��i�Q��?T�q��K��Y� V�1m��r�_.��0� ������P:�ᰉ#d�bh����oY�H�V��9A(��iUΰ�0}HTO�v5�F�9 )�^2-�O�z��F�b��:�4X�Oj7i6p��%`��R#+�ݏ�W�/�)M!�;DK�C:鸣PM��S���DbaHS3"�Ú����|�Gk�����+��u_Z؋ǂ7�/�E�7�x���V�<���%����3*��kV�܆�O� �n۠|-ϧOj<K၌ ZI��i�<b:�J�8a;��&�����p#�����2����3cFڐ��L��6��}M�v5��<AF.��Ƅx���/���uG�ʛ�>#X��_����k��h�����Y��1�뵑��;�31|}��Y�Pz?��VngG����|?���0�_��� ���4�~�Z��Ah��sK*G�v&\ۃ��"�����Z�����O�CZ�7��΄~&�d8���d=����K�-V���a�9:�Z���M9�z�nH,Nw�t嚷l�-Euش|��@�u{��:��=���K�xը��hH��>��$��Ȧ.��9���a�|��~r)�����B|Y�n?a�o��S��V^Hfت�K@F�9&�U�F��3�5����G(��@���PD[ �c�ǌ
6W�߽q�x���+�$�4+���oi;�i�mq%ef3F�T�:���Dr>�`/�q=���������=�E����i;���]��L�*�~���&�p�2}�ɶ���wgҷ ���'p��l@�z�f����ER�C�r�}��'�	Ȏ�W|YA���q�bM�M��8<���I$�5O���V�?@�NR�h�����r��S)�dg�G���ڒqКꁚ��E��-��uK���`�z��@R�=�h!��=�Oa�E%��y-��h MW��P���f�	e��۷���J
Ƌ�m!�j8H�0+M��I��|Ѡ�����*���ȫ�-(#�=b����K�����8j�i�Q���IԿK��]p0�����L��{䚭��K�l	��g/ibU*��M��O�\3��;�Fv�"	�����	��J���-y�3��F���FG�%��{�bp�Y R4��<���7�ӂi�s6��5�C�B�o��T��_��/Bz�[���a�#����Uj-ٌx8��&��-<<
���{�^'�n �Iܦ�9'Ni�>��b�'�{�HA�Kp1|��
\W�<w���s��������!��⣇��}�����>;��MA�Wv���T����� ڢ;�7��T8�42"����s����p���c��(��=�[ͱ��G�0Z��0%!����7�z�ۻܖ)�v���-ӧ�Oh貍g;�8=[�~tA:����d��'W�:IH�6E��0���떍h��Xo�U�V��g�_A�b����>"�.�\V����0E°� ��T��B6�zr��_>Q�����;'��6 �?5�{o��73��K��E(� �H?!#�Kn���v̓$!�eg�����1�h����)�ܕ%3�<ET�>Փbf����B��-��vl跹��A��:��}f'E^�	���[w�v���С�;$tV��|A���m�������ʯ�y����)P	�v�ˤ���SJ"��*���4\5O/��4�>�������3��B�(e-j����AEb�q�fh�0�m�b�G�"9<G^P�c���y�Q����"�O��'��!�r�Z���&�����t�ou��u������	�ĩ��z4u�_�.��
<뉑�g����1c�pIѐ�jp��T;�n~U<՘*�T_C�m��Ʀ�d�G`-��Cy����6@sӎv�i�l��+.Xg;;�pV��f-YFU"�Ƚ
ɢ/*>fl�鴭w���� �z���f� [>%4o��s���ŪK���.u|ˑ�3�ᒈ�bp<z��5�+/G��XMf�������X����fy��N�����SJZ�CvP��{��z���[H�^�M�((��<����}�{W��K�YK��	��ٗ��`^�ɷF�1J�v�s^��2nG2�����%M�p*3ftZ�|ԽT�����_�P����o_�l}�����n�]�F�Of�
Cٔ_�U�{���k#(gv��B7���
@������y�O�C�<Ѭ����(����f��)���bY��u$�1���H�c����\��٦M�}/,�cʿy���S5�&86��:+{3�Y ���d'��4�ђ�H�������W�|J�GH�f}��㫶a�k:�1S2e�@Q�̭��6
a���e�X�+@��C{�)Lu4+C�n:�u��ށ��|��hq7>qD@�4������&]�����.��aQժ�p�y#�O_�ʫ�m��Y�-m|�p����P��m�wEO��4 b
�;��t�r*l�R����e�?�A �Ά����e3�O���`�9�'i�)$�\�Y�x��n
�P|�:�6x";�����>���H�~�k����6�g���Z���tg�4&�Q���s��X=-%��ɑG���a{���h��s�7�<U��	q�IY��13�m9��8�F-�f^P�uGmO����:�-D�YG;�����uz����w��� ?�@m��3�Qﱕ�a��b��Q(IE4L�k� �-�	��Gٔ������f{�q���W���������d9֠�&R���"c�&��Ǿi�I��~t�K$<��>,��>Z7@��È#}I"
��`S��m�y�(�ۣ�~�����������(Y��u�Yu���|"�=�H5b��m�����=D]p�ϳ}�p���ĿS`٠����9>d��h4��}�#េPu�>��W�1��� L�ۨ����>.L�b���X�M�њq���J�T�4_K.���u�G�y��2�Gc�p������PO+]���ڄ/-]xw�}�GiZ�'�T���-��ʇ��Ce��P@����P��8�'�"�q�3��"���f9a���0� -U�Y����l�*&��]�f�{S�<^�j�ч)Z�:+b�8_O��:�H�f�7ʟF�����tw��1�@��X�
BM���U�0��I>!l7E}g>�$[<�F��R���guu�F�}�B5�؜@���{����}f_�VkO1��S��:�k.�S�+�HZ�atJ����n ������Fխऔ9C�͖�נ�;}͍�잌;R ȵ�H*�N6��
|h�]�@J�g��.�-w�`���p�F����pw�Fj�U{���M�B�)x���'h�^��3,�=�l˝�_�م�>�h���gQ����Ѝ���V��6h�eo�/{���^g�~��bd��C�\�q�Q�$&�(�����m�:�"�ZcI�RӒ/Z-�-gm����m��3e��`��Z&���/vWA��dG����]K����W�/_f} b�;���ǒ^a��w��?>�Ɉb.e�����(}.��:�EYbW��zS�y/aQnD����	����N�5	�m�ڠ�&N̾$�vP̉��˝"��Z�XI๭�®U�}�S��ƶ���t*<'�:=���o6�-��3HsڂjS�����b����'��R��%Ԕ�K(�A �}�Cu�
�����РE=u[t�e�o�^A|�ZmE������6z*�H�S�x� 슡.��<߈]r���'SP�1Z��ZQ:�|�Ⱦ0��)3�W �V�$ImU�_ �CG<�Ob2���&[@��_����h��hY_u��z=MJ$�Q@2��i�gyu�#ޠW	d��2�fɕ n.��Ze%]�z�h��w�Dk��58bi.þ���8���B�VBM����j���I���p�u�b,� �(��
�Ո����[�<�� X�@�G����S���f�ީF3�TQ���a�����TwhXo���V�ݧ}��n��m��1��jX	�?E��.�q<v�έ#�Fb��C�q�y���䍄H?�{&��i�n���f���p�D�zC����#�Z��}�v5��/\�� &MR���
e��P�uf^����|^���6J�Z�o�K��j�C�FD0��A�C!#��V�������S���4���� ����7�`�d�
j8Ю<	_������\>�=n�p�R<��;�����7!%�Le�<�����.}��O#z��Y�ױ���I�]���Eف�1����@�R�DH�����\Ļk��@X
Ȩ�.��d��s��D�µ�j\�Y~�����﫴�Vud0�>QlJnP�O������n�AA��΁�"�����!(?��`����v���(�������e��(�i�?@�_���d�Z�t�{`:^!O]#r�]![�r����=��w��Am!�A{�=�	�HPJJ���O5�lˍ�K6��/|��\�')�g��r�9��/A0�f�����2{�L�	0�GW^e�v�1�]z��W�A���Q�:��s�aO�G���g�`	Zc��Ї��b�c��@i�:���Si�_ѼW��Խ��t�2�)a�Oy���=M�ED���[��g%đ�5�Ύ���XW]n�9Q�L��3���kj� n,[��@h:N�$	s��X��o��;���(�G.
�	G�hF����@[�4���ɑ҂���S�zC2�lZ�~��'��+��v�o�b�W��I���gE��MfE"�	�8��4x&�|��m�DNA��̒�K&z)��'�X��ɰ�����y��dn�0�������7vh͂@b,��T�!���O���5����s{���	�J9՞2ň�ۖ$-!m|�d�7�d��ء�~z���x�E[P���a�D�T~
��8�qQ0JQ|v �òX�5ގ��YD-��w�����p�ma�DϞ�t�ִ�Ѕ�o����v��
�l�͟��č��5�0���̰MDM�Xp�.���9m��J��^���(:ܺ�h��Rx��p����
�����*��<�&�19h{�lZ�e64G��H�߀�*�4��?�����S*=i�����s����wȇG~-�!�)�u���L��T��2z�k��f���8�ϙ#Z��6x��F�=C3L����1[���3Y�8�Lv�
|
�H����51��n,����Q�+M�Q&'���*��p���ԁ��}ȎO\(q�4��?9����V�G���!`�|�[ߺN��j�,I4\]�%Bي˝� K�Z(8�l�
�6�/3����T�,]��?6�"��4����+��5N�c,���S�uzX����l�U�\
l��k�[�kim�F�Wa}Ӟ!���*Y;0�*u~��/��?6��wz�f�z]@I�D�
�X}��&u���ZI�5�L��V�p&�\`����Ъ �y�LR�$�f&�m<�	��M�K�pJf�G� s��<_$5��-��o ���Q�p��u�,+n)W֞��3��~��a�@e�{X�	��9�����X�v�`�s1�����h3�`W�D��cx �K��b��m���-��!��"aN���d�r��Fڡ�n�%�v���P��.��a��>��Ґ�s�,,�K�&�m��
n�=�L��;�\�R�o��V%fR��P�.Xi�(����2���p�R2��l��$�>���?�&�1k�L��,пs�jl��i\�yc*��EH?�5�Lk]A��B���B���,J��6O���L�M}��\A�E}i��f�^ER9��aة�~y��K\�P������o���#0L\�"�8�-���Շ�D���!,����vߢ�պX�q{�s���{KJ�T���os�[�?֚g|p>�b��������Ԏ@\�(��
M�-�E�ؖ�՚v�(�����}�r��a�J�'oe�[��ӷ���)��rm�:8χfy�^!����"}�,��E�%�\U�������Cp�'���6ۀ���G��(�Ѹ#���@����}j��x�P�Ѥ�F���3��<�n�Ld��́����\&���0�wpC�R@�e�����Y%""�7��ļ��'����M�C�@X]����C���N�Fl����e�T 2��t#ʕĤ��)G�>��L��oջ�Qo����sE�����'�a��cQm�F}e���'� �yE����"���\}��S͖���.t�����F1���{zT�Ƅ>�/m�n��Y�I���mN�=�^2.�U*�z�āQU�xec�u�`�=&����Ϟ�
 ��P+�e'��o�ߔ�3i
����	���ѡ�`~\jju @�y>��B��W*R�׹k�D\����p�)�u��ܱ���>����g���������Ϋ����Pf���b���]�28bF|�(��3���e���4$�񛆙bT] ~�R|Kh�.��j��������5�j�Vk����E�Ɂ����9���� ��*����ƶ���h(2.���kT���Nƚ�GKn��z�{�i�b���4]u_�N�� d1�NW/)��F�i���:�����i����Ǟ�G�v��g�
�����}�G�D
�:W���Že��Gz�3�(��b(���Եن��9XJ��b�����M�I3�=ǩ���y|��&�85u�Ń�����n�*�{�T��hO�ų���m5��k�ڻL�Z���io9cyo�-��/V����P;4�i�S��T�!�Q����8tj5"�\R`V�[��oɑ��vh�Q;!�}QpO*&=,M<�����-�'�~k���x�hz8��э���1ba�??q|�<6o��iA��w������������/J�GZ��m�j�f/�Ϲޞ�e�z�pJ~�Ǥr@J��bd#���n��t[�m���<{�M�D`�.cly��?
E��d�ה�Q�^5�,��֝0ߟ�m��)p[_<�����-UD'�fL�R���B���3��N����i�� �X�#���]�̣Cd�>���p�nl��U�9�X��!LY΂��`R	�@��5��@:��]�4��K�
����7�t�'��[$Ғ�#��P���"�=S��,ݜ�F�o2��ǟ^2���L$r�\*��ǐE� $��5���&�]2`�w֍����e#����awyz���bZ�t4b2}n���i�j��攏.�D��R�t]+����h��h��&�&�}t�O�D�gy�{��Q����m�ˇĤ ��)��g��jAx�1VA��<�7��~[ ��|MYq���(ك(tEPe_����lE�O@��h����|{ 2�l���!4�ް}X���������u�6�pbKpC�`J�AV,�N�	�$#y@�F��hG�����!�/<=��S�0P���ɀý�h��&c�泔����ЌmF=��ϯ<_�#��<f����0�:Qve��NV� Gk4*[ǀ: �Ӫ�9t ������$�4��R�3p�,00G���82:������F�g��Aa�=:$>��y\D�2�E���Ů'�6C$�tC�Z��֕������pd��p��Q<NU#��H$��+ڒi1�����|��ֶ�-��%����PJs�Ds��+N�n��}7zN�����2��}դ� ˧D�`�3ʬ,-��}p�A^�6�P���8��i`��ȸ]�6���$60������?~b�c���7�	�rK�[A�y%و�Z�1�9a���TN�ߝ`���:;*9����O�9GDw��qV/�ܜ� D:��Q$ЛQ�wƻ�o�i�[�K�lU�����(4�A����3��|����c�Ow�zC����M�@ߝ�G$�x\��*%Xx�)rA,4u�<5�����g��"V��^�z>��}ԏ+4$A��U&��G��j@��eDNu����fU?���޽"au��撒�m�=��lSY��3�C�v?B<L1���Tti"o=Ί7���F�2�ED}�:�Q������^�����
�2�� ��7��.����jT�����
,@��x-�Z�����2�#w�R��q��[��y'�gx�FG�V��b`_�S�y�D!���ɿX�&�?�� ����,o�z<15�իƬt9��x
���Q��:�L��H��As��DïJ�@�D"Q�I.�� x*�r�wg�8)@g{��$��ϖl|	��ޅ��i��Ko�������-����,��.�i�PV/�7Wn;Mի��M�OV�_.�k���q4��WT+ƪ^�Zt@3�� 觚X�*�3	� {:g��>�R�������=�� �Fa�>N�ʏ^[�G�_~E6CM"l�9�.K#�Us��g)�����P0�=������0���w�Dv�@��}�
g+���ֺs���ʀZ{�����2���}�9qY�	���[_�>�U`�=�byD�+�c��U�o�*W��ZB��TC? �T1Oo�ev�a�C%���Q��:)۰[̢�^�����Bt�(��[7x3٬�'�<Em��O�
��HB1<�]�*׵�'ƭ�"*����|����hs�����<�ʘ"^I���$;jE�,� O�*�������a�ven[��N]T��o�B\zʗ���h{M����5����d�������6Uv[�%�7"���c[���eڄ>����>�s%��YZ����ME����)
��*�S��9"��˫�mC�jCjp��
�&)3K����P��@���˻�jq��kY]��b�N旻p~��+�E�H��=�lϓ}=�1����E��c��E�E&�����is�MW�N�@�N~�$ͪ�A�QlN��?���6"��Ҕ)G�''�����(N���!�[�����D���BS���b��)=�(:�M\a�Z�ܫ�F������v�l��؛l=�f�'��6
:��K�g͐�p(v����W�7)~�}.3�{���{ğZ, 0���"n��آ(�"�Yc;
�c�Vֿ���$�V�	�����5]�py������~��D�oΈ���Y_���[h�yr��oo
��S���1�YZ�yW_�:�L�LCYN��{�n
�ڍZ����s��F�c7�f���ȑ�^Q-D�"q��JOu6�-L���u�:K���&���Վ>�q?o�Ė:��vD�,[���U�=��$��#;�%�Pt�vw��b�Ы�9!������My�C��1Y����b ���x�H��q�4D�R�9��;P�����c�2�a\���_�7+ٶ�7�Y�j�5�nsa�u���Б�.wq�Ս�5{"��뙟� [��}��;���$�<ma��y>=��[���QI&j<늶��T�o���x�p焎�n=�&G�Ym ��8���X�Ma�L�e���ծ%�z%!	Ou�N�P�ݱ��J��y������ۿ�;��^f�=g��L'�{���P�����4z���jMc<����[ܨ$��~�M݆�b5�a��P3|��ָ2��:��������Eԟ�U6;%;W1��A�|/��w��c��y��M3�S9���~��<n���ӊ�k}��Ν��-��{������V�m�'wb���EUN���?���	"u��qXj���i��M�)��#����������q؞F��T�f��-ʊo~ *�@�PcN7ǘmueM�G_d>R�����Z�v�����7p����RA����-s�L���Y��'s#5\k�j� !�]�q�!fud��{��g��NV�^]aV��J\�O$4��U����)�zN���b5"'�ֵ���`׃���\�1*�{���z׸Pœ$+om;�3�?&�?���"�3���:)�y�H�wTU�R���?�A5K��iZ��0X����Ŏ���*���í$}���=L�:����F�C�n���4���B��B^PPvL���7�$�lQ��P*��]H?�:�$7�؍_Ų�,���sFm��R�H=Jt�ܭ={��.y��{u(�(��ГbPy x&ȼq����.[�:<��c�x�ʙ�x$�Y��U@�Q�(Si�$6q�T�DZ���\h;@�ӏh�@˃�#��6��Q&% @ԏ���Y]�j�ʊ�q�R:ݮ�-eI�Q�|Q�7�*����|j�1�~cW	�R�%Mh�o�HƂi��]���nI�D"��r��a:�Cq�g��0�����v�돣/�G�Ī��`�x$(7����-������I�7���94���:�㺁�#���qq9���@*�)�}��]$���j2rN��.F_�j/Ӟr|+�r'?u RB��vM�e��&]��I���<���"���~GnW�ۯA�W&;���(�)���
r�Y��#���P?��Sjp��������#n^,xrN�,����T�*�<�t<�m���a*ֿ��r����e  >��:f��ˡ\6�����;���_K��pTV�u\o�Щ$f䋋�=�vP��Ώ)O�*[ս2_��xX4Wb��نtK5J�:��!�&����=A3�2����*�`RD�J�c�ҩ�b9�����^LDC��R�j�4b%���	���9���?8�F���H���/��l���3��2T���O�9��c��舼Pv���T)�1O{dQ-�@�(��X���&ַ.�u9�%�)Ƚn�����ɲ��χ_N�3���?Q.�#c��1_	� �ַ1��F��ۧK�J����,�.WM�4��Y���o�� �B�Ī	rN&��y&Äl)aE����梳d��� �ᗚt���uog�nV�<�P�`�U=S��7;~S��sv3���pw����J�WW�n!�2K�+�T�˾�Ra���W�U���߼�Z�e������iσw8�B��p�i�ݚKw��}x�@iC����@�O�Z�՜��oj0��j��*-.o���W<M%od�4����,V��y�W��"O� &��Ww/ul/z���a��l��n���e�guG0��c��MqA�U�pP��ut,Q��������)ӵ���|����/����ؚ]�$��b�v�N�Ysl�����(י���X�p��x��YO��k����}���o=A�I|2�n��˷�<Ps����8����4���+t ����O����[E����Ҹ~A��[��}V�P�(w�J`�5[˟���!s)U^�ԟ �
��<�i��$S�$��EqA ��Ԥ��ʑ��B�
��̄cV�M&�xPi�]\�]���"䞊0�=�,e�'y���l�!*.sip�z�����N����s��$�+���1Z��?���|c8�ν�W�6M#U�[VS��;Y��3��.>P9�4X�Ou��6ۮ����蓆��%<P�y�<O��f�0j(X�肯OE�Usw��g-��&��Z�*F�C��ڱ�V�bR�BJ�s�G�a8B�4��2F#���'��ί�����; ���lf��Ǻ?(�!%ނ�K��6��lbj'h�^��F῞愗(k(H��2@��E����1�a�dyA��(""4��%���z�/T��P�L<[�
l��rTE`��U�ۋ(u�x�kH�7'C�`2��%M��'��b�D+9N���g����B�V���lฦ�RQ��D]����8p�ԧp���R�T�,4\��·�5�G��j}��d�V������3a���<��-J6���C�� R�
�l�"?
���座����Z ��g��	���\6��f��{�/aKft�ӬN@�P#Ŕ����D��G�������o��6����/3.�P�r�+�_`H�ը��Z�xy���:<@g�Z�0����x�ɨ��[�Yć&�G����^���������	޷�V��t����a�d�Q�
U�ӂC*�=e����fy����+#��jn��(����D���nF�H�^�c��p��<�tn{[pr�=�$^y����B>w%�!7�"n��$\�1AL3-p!�vH$� �w�l,u�I��inç�qc���]l�!���CF̧l��Z�fUTi0�-\�q;A��t���'� �Y׫7�������2۔��db�-�?��l�o�$v�#��׫ɗcz�@�����rjd������B�!.V�@ד
j���Ģ�jL:&Ź��Nb6�)���:;�|P!�� �68�y��i����>��o�0}��;�O ����ڝd
2dp<χ��65�4�<23���gċ�7�2��pI��A;�A�E���9qƿ8���r��_Ǔ�?�;Ө&m;��ԁfw�'�����!����K4��)��ԌM?���)�̦��t�'��2%�gv4:Ě�(<E�m&%v�n�xj��^�K���Z磸E�3��Г���EC>;�/�r)�ѭ.h`�񃬃_]��[y��G�F�B��
��.��^�"_-yx��{�H��ݝ�n�U���`��d�?�(��CGx�[����0�!�Q.��sA�l	���Ǟ���K�'ѕv�@�eH鱊Bz�'wm'W����F��㺝�]Q��	� Ԍ�Q�:�&
��R��_AP�����TC\��R$�������ϸDf����Lh��T�{CH�s�+�����C��3N���ݳD)o��%���[+M��f�֍{�
��A�I�V�'�6����2����J`��KX��V����S�����M�nQ����E���x���[�RL^��F�u)�����R�T,���ȱG���(���X��Z�ɩ��HM����!|M�%��R��!���Q��ͷ�p!.�1��[o�xj(sϡ����������t�����'̮O�ֆ�ZAب�j m�7�d��^���F���l+9�PY��t+��4�s&�L�Ϻ�'� ?жgVþd���֦pqJ42�0����N8ew��SO�s�;�K�ii_ՍXl�t3���E�S7z���;6S������E�����_F����^_������{��'�ޞH� ��vVp=��~�����>����Xڸ�4�>(���22�tX	�M<aU��cl�:�7�_HD��6�V�_vh�Dv�̭wHBbdG܅��*���"��m��l�v߸�M6�g|��MB� ʵ��&���|�X�Qj�6��� v�sZ%IB���zT�R|�ҳ��#��B���H�-�{Z�t��f��EM�a������q��� ms�?>�e��y_Y��tq�fˈ��!����ß!�
�`��������.C�^���g�%��A��	��`UnPB�O�\��g�#���.a<���t�9o���pjx�b_�y+�������d�6PE�����r⋜��lxx]Sq���qU@���/���L>�EuӾ{%����ܡ:�����q���<��S�2�H�O�w%>#�P�:�L8f$}B��Wh����O��}�LV,>� ,����^,2eEy��w4U��റlڄ Fa@[�X�_�Rض�N|3���$������m"+¦~���"D��g� ��1o�Z2օ3Þ��/*<9�$
.�tCͿ�a�����ٿ5l����ˀx>�;��nߖ-�)��՘`ǁ�Ji&�1C$��L��j�Q�W��AH�N;��C;Ĳ�������M�H�M���m}�s������&��X��w�f���5�����{u�:w��G~~�PU�*,mT�� (<ғϝ\�[?�����Ҏ�0���BN���n��|!f�v0��r�BŅb����4�
nI��Ak����V�4`C�4�xJ��%��m?9�ߍ�t;\t� �'�Yk3���>���()� ���zƋ�=!]��W�O<�I�Uyz;,0��u������O>��M��Ufu��\��ke##}�K��,����fJ�"D�^QgcҜ��q��y��� ��U(E��dP����^�	-��a:��9��(� @&>e/;�h��Qm�|�g��X ���$-�� *�z�s�w�~��4vp�ڋZi䁆�:E�T�=��Vʪ�N��nf3ZMm�������?�H1^��UNb��1�߂����6,	~�3-v	�M(z靦?OKG�D�&v�| p��ބ�n"�F�e��FJȘ�N�&f֝Jԥ,�+�i�� ?;3����&" ���r�OHr�@b������3��Q�A1�*�U� ������Q�q`��|p�}u&�эb�=�[�����K�;���6=��w���|�R�����8�Pv�����j�|u�p��>��`˭��.���m��	���J�v)R� oB�?�����Y׫�֞�H}}�坬�XX;�� �/|���N��X���z=-b�9��CPM�5�D���pp,��-�W%�������h��F��9>�r�q��|{��wE������H~�x#�W�yd"����t�3�Gx|�^�;D!��C��J����9f�9f&�AP���D%�5D"��t�����R�2����:j���c>h�^fǥ��;Bd��۹�	�B��0�0e(�.�
�5����F'����4Q)g�gx�=l�l���ˇ}��:���GK�5���$e��q�cz�k�~���n�"����;�d6�L��KF��"�L�;��8��.* ���q�!�Y��e7�8,!�w���"���Z��(�\���X,�z��;�*�����e���t�������+9�=�V��+�n����4�>킷V�~1���"4�z�)Z<?��r�(�����,:��o"��~UmynP>�,�/l���,���檥����*��(���:���������>(��Q<E,��C/�&��V���Y'�|j��`]�G���4:$��$�Z@3�j�n�\)ꗭ�О$R�A��`i+�h�PV)����oG���s�Q�Ǿ�m	-�ky�1 �u!	E�e]�6_]�_���y:�8���o�y|(B�5y���|v���$r�4���bÄ+/�Z�Afؽe@ ��$1��{�8I7>����]�F���ݮfB�s���Mq���k�u���C?�Z5%�3f< �Y�)O�����0+PPF�����H�������U3��g�����'<?��/G�'�Ԛi���uҍ[y\fCo%O��9U|����]T�V*E�.1���'��8���d�M�+䎼�Tܿ�^ �}���-N�
������6K�����.�j�ɾuz�C�;{̀f[)� ���x���N;�J� ����3� ��ѭ:L~J�
W�=��1"D��-a�ǵ�B�*�R��Y�FX��@<m�ٝ��#��Ms�o�ٯ;�s��\ ��.�0����b�f��R��C`��������sBK��P�;+P��p/M�����xֽ��g�[u-���G�,��%��w�1�;]����;��֌����ڸ����i {�rVg޶]�Y���k.a�Lα^�)͠Mp�2qU$��S����oK���Y�����ܣ%�F2�ߦ��5�C�(�ztH��@�����=�YD3�����ۗLc*^�����>�/�	��#.RȚ�������4nEz���;YW+u����\+�+?�~�$�n�2�T�i��f�����6W{Cpg����G���d��f1Hz �ʩ;Rc8(�b��;�x���h��=ę8I\�F��Zy.��uɷk[��ث��o��M�Fd�U-w8�M~w�����E��ٱ	Y߭�匑1���־�:s/��]�٢�dq0�=��k@��9j�8J�u��=�Y1��C���#8��%-���2�Z��?�'Ї��Y�p�O��Ɇ	���+�=��[	���".NC����@5�:U���˧G���U��4%=�a��ω��9t��}H�}J2굱�9�|N�nDG�n�$�p��};��š8΅
� ���3�eEl(�w�ER��ڂ��B���EE������ɖ�c{�M��ݰ��,�L��L^D���a3��O�.N��̂Q~D�~��֣������_�z��y�c̸yR���T�/#����4�8��	@��_�/����q4F�߶=gp�g��p�EH$��}[�G�Ǝʱ�b.��Z;�Ң�o���Y=.���v*B <�v�j5��N�l���r����|9�.���5��V]�T I��i���f����~Go#��I?�����nҸ�=�6?C�7�H����#B�K��a�K�hY��G�Oϱ$���q;vޤ½�G�&�mgDz!�1%�Ra�����cj=���9��ʮBuԘ���a<$��Qa!/Q���7����G���yn�i���)\����Y��A?�%:a�q�BZl3�\���vq�Q���ٓ���'�=Ϝ-4�7�wEq�KA����A}��>t��Ԟ�y�{���r���*�X���x�jˢ7>C��;����IF��a�D�lǛڝej�x�8R��&����*o�(T\��_s�4���uX���N>2$�u���I=�/�,yo�s*��N��tw�u��)�]O�S&0���W�w���Y���k]��	�0dL&��:�L���4�G��.q1��?i
-���Pt<��ϙ�ܣ��Ϊ���T�I.�1c���Jկpe~�#�w��%$%�f���O+z�e��D��b���>jxckX:q�X���x�y��n�j7)���փ�?+���E7�b���3����~з�+v�FMf��E�(��l�W7w�"�}}Ns�)k��/Z��^��;��st[� ���������1{�e�ΧJ����R���N�0�Y_D䋼!���T�pQ�&�X�k*�/ÌkO�vap���Ƶ�\�2���0�mg�TQb��DZN[ޯ�6�G�
�s:m3B�u�u���W�,�D!|H��~9�͏<H�mE�(8=g�`ଶ�[�'�R����ǭ����i�M���-O����ȥ�c���oNnc5���ǯȿz����J���&���P%�l���P�ۢ��w���=e�b���hH��Zt\J�� J@A\���U���P�J�R�a��Y.f�>l̶���-��G��X{2?�c��zǭ��4$�"��M�2&���;ڜQ�޻DĹ5��`D㲎gX�YJ�&�oZ��Մ6d��L������o�=�ę[U��`�� �8�E�w��>��kO(��k��U;8R\����Nܥ0��"���q��]�Ι��UK	�d�/��̠h����Wls�7��=��i�j��S7:]�wҍ��M�@d�l�8M鱝�_��H,K�OG�PE;ez�kT�[�r1xD�ߝ��J5.,�|&5��x,zIz��.J��g������P��z\���`���'d�|���[~ov�|c2�1N�7���&�Qq���*�"w��r.$�E_�����1��m��jU���!���at�'8r�U��i�����"m�n�21�0���8���˹��c"��Z�s��[9$��n�5�b>�ʫ9��$-�#�ҹ�F(G��`lz1X�*�+]���:�5��X�^���ai�`S����X0���q���[�-M૦�U����H�� l��!~^v�RD�Կ���0�59k�БZ����㬻�� �ܟ���X,�=�Ջ�`{��q�Nc���9���b|m�_�gNX��C
�˧�,6;|�]�0�*�&���G��aw��|����Π�6�z�ҫ&�M��*X�~y<��:�vF�$�Q�f��+���ƨ�T�='s,�
=�Lw�J~�NW��� 'p>Q����RE�����@,�l}�SY��͈x�і��O�H�^�օ��֣ݞ5��=
5*f�$hr��q1��WeT~��]������j��0�^�D<��s%�(�`)�K�<��7R��^N(�QQ���������(����:�`4ǙfnW���"���k,u���|O��5������"MQ�
�칇��B����H[,ln�C�z��9 
�Ic��@ESx�����h0��^��{C"�T�� Vu5��~Q-$`�.�Z�X�@���ncF���4~,���J�^ �'�e����αN��!�`K~���%_�CMY���-L�e��+ٳ�WЃ`1��Mk��^VVg>�޷,0�Vi��"���;w��*U^h�&�
�%�c���9Ń��o*��=��� 2�JR1���vE����~X4nL��a�=F-;3����D�4���Y<NX�S��L0��R�zp��O!��X�,b=�sv���/�MN�$%��_:q� Kp����B��ʻ��^���r�|�_�R�H�y�K%��8ֻ������;K������ٯ�a���rY���8쥑]��hn���A��- ����_/�Ș��s���!����X�Ъ�T�9�K������KI�̅���ɳ�tM�`L_�1���2�q�~H��~���n繱i�|$鷺X���VL�L�M���<��6ڐv��F͌�� �;Z�!q�v�,�BlR�����EG,�"ً�Z�]�L�k}0pA<�tt9Ҷ6�),��x-<����g��k���|�i���!���k��E�4��\e�?�Pn�Ȏ&��E�Z�Y:������Q����!'H��4�2 �+�ʹO��C��L�A�*�lF��l��D��HŅ���;ґd�q.j��*;0Q��F��@JI��
G�(�&��6�p���R�T��-�Ō���U�JNN��ܸ�_zV���@<И0x��_C �	r�b��������P�����R�BS�"tZ�����E�׎	�B{�C�y���?Z�-MQ��r���&FƟ>���%�.��5��܍������%ѣZ0HS�Ol�㷒�,�
��~��W֑����ԙ���@�S1j@�]kXP00�?cO��cI�iyZty��*,�I�h��������f�N�Y?AhtL^B�ףP*����Nޟ�>�Hda�ä�Ix���3O�.3~(����������JN�����6���nI�/����F�MxE&3���
�Ȳ�'d�i�j�d���Z��E����&��R��s4�4Չ��0�ء��Ρ�n��я5�J%�Ļ�$u��o��zvR��<,��#;���F+A�ԝ}�~�ݜ�}!D��)��֮����}1ݳh�o���O[�>��I*Z=��8/��!��2��
*�����xO�醻2�ʟ�fV�u��ӧ� ���mF�Mt�j[p���Cka�&�vq	��y!:qP���5��:��H�?/O��������b�r>�t"���z�e��^1��6w��u�vk(���c��34�c���Q����>W�o#�_���L��=���Y%ܪ
�[$��9i�� ��%�,Nֻ��,J��A���^鐲EK �%�6�^���G{ۣ׫~I��8�H�6���B��d^p����SO#A�֎��%���R����C�s4���{(�(�WɃ�����"�_��쵸�oNﳣ�܄"핱��Pj�l>���0˻vgCO�7@Q�	�	r]0ɜf�a����/ n0�i{ �'�cIv�Z$�d��xu�a{xf�[����2�DF�E������t�̽�|�Òq���=�]B�8�Yଐ���{pܘ�uה��KR�7���s��24{�Bs:��?������*�8�oi��ބ5+��L�;b.W�aD��G(,�H<�c��_{(X4a�����r�f|�^J
J_P�6.��;�=0�",D�5=5�mU�!b��M��x½�u"(���Di�~u���'���8�{^)q(���Y�Wu��zka&�7��J�����ä�y]�\�=l��~�ex��2����K��=!��
�rY�]ew���z7��9��E�� �D頤O������*p�����h�V�e<.�A/��bz��w	��)���Wq�����ۦ�X`޽�{��p2KG@�Xt2�n9ud��ϻ���egy��4i�,��1�_$?fB�rL��,�%v٥�����m�"��{Q��	lU�/P�\_CǺ�@�H�a';S����7�8��M#R[`���J��-96^��i0��G|:��B�@�:P-dX���m���
C"�id��G��ͣ�d{���9jW$0>s(���hyn�f��S�*	>�[Y-�~�р�m�C�����p���ȳL����2��tB*��3) f�����8/E'���2��p,�ڳ�ڼ���#�T�d���b��y������	��T�n�6nZ'n��m5B����2l��
���0 ��k.��ǁ�c�~�n6q#��2 ���pp�F���5+�?���m�k�>w�)�S���6���0�#+/m�P��]3w�B�cîqsx�yn��f���-�.n^�S����]�-�@���j��49m�{�qWuP�u�*��}G�@9n�oJҰhD��̇{�œ{t��<���S�nÛ��,���d2��C���]eז� ]ӝ94S˅�E����d�)&+��($��S�����:8c%8*p�Meby<u��Ou}~��6�����&��[*�E$)OS�����$�S���GxEV[r�yȺ��~Sb���	���[f��ۀ��\ӄ�!h$�D$�_��PR�3(�9� L�n�|l�Oܖ�P2� �h���Ԟh �T)G�����Kk���{�2d���]��D�U1�$~o�A����b|Cq�A�pˊ�h!y�$4��ñy�75ڕ�>�����i:�S�T�,?�aW��ʗ,P����"I<Z/ͩ=���`��H�|���2�i_��'�J�ا��(
��ľ)"��tř���Q)�4f �ٽw��cJԬ�*3�MWJṉvk¥��a�q�AnXe�x���X����b� yBc��C���ҭ��`5N>�Y3\�
F9��@��L%=��]7Bm�
n��w�i)O����K���N�|�:�A�3b��M��1���m-K�$�²����̏���ӑ���uoyH#ꘄ
YSe"������k�F�w�p�[瞈W^o=־E�{�r軴V�d+y�um�YvY�pA�ك�9��-=��JU�1��1E���<�����
D$pg\É>R�&26nӨ�kex��3.�-WOMpP�󵯤�<��˰��Y��-W��Mk?x����+���ayKك��K���	��Rd�!F�9�n���]�q��c�8ߨ�M����6l��#~D��@=C!�����V,NX�9�Zw̱�l����:5�<���k���k�7�I\�+5��]��v��5]E�����
w�X�~<������C�y��r��o�A-P"�$3q<�{9L� A�Z��}��S��p�~Bd�U-�	���
����׹a�����MH�*�$kD�p���r������[h.�#B��Mu�"~�tK1�I%��o\�r�m�֘+`y�)ĒK[?[]���+��� Y��j��E��?��Z�	���m�TZ�}�L}��Ӄ�c�$~�@ԕ�*��ʻD&��Bf���#�G[a_A�B{k�H7��ﶄC(�q�X"ǵ������@��K�<s�<<��۔Y|4bj��J1�4�J�<�J��׷ʼ`[R+�kUo��9���Bb)lI�M��2����Z�u��R�g��hC�c|��ό���ݢ?�XH5�����C"c#���%eI�����蠌"��Ay����:	�ow��S�˳MՒ�h���IG2\�q.r�3ί�E�0�Qp��
�,��$zǎ��_��@ ~�;��d�!���>��v����Yh�]ѵ ���G��k���䲪����XcE��Zj� �&���n��XO�,��˘�233t�x@�BA��*�hoO�W��w������h7˝���w�-�Nj�Evp�gkP�m��!����ꊌM�6;��_%jq��ՈOn�����iWA��v1�F��"�����;��n�����<���/���w��«�i�o3wz��3���Lk�lb��S\�s�G9�<=�@}�Q51Y�K���OG7����������5#n�/4
�M6��6iG���?e!��@d���[\��x�'NY1s ��/�1�,aL"���� �Vt��~1���R���F�0T�ɓ��r�d����6I�d��9�UW�X��c?�2��B��/���l[�U����b�Z�I�J�%�rQ�^z�91{�6�&{o��������J�_�|F �n��(���X�Ӻ���Ò?������"��%���!��b���O��#M��/�""��:���Uq��[���4�=O[���Ԝ���	~�N�����]�� �-��>9�%,p�rs�ʏ��<����t�+��_DA��#�2��S9W�d?�ǽ�L!���ms0��\����ӓ�a��2������Ƹ��J�����L��­����H䘞�4�E�$Fg�s{����Lg���u�i+z���F@����G9��֕�!6���<'L��3��D-�Ғ���~�t��dN�ج�[����V��!�-��.!�8=K�u�|���z}�c��x����r�C����4��kٮ�j���C=�m;z�dv�6Mx$�l~y��*Wds 4(�Xǃ�nn[��,�2V�y�[	�~0�*aٵ���hP�:�/4����]�):X��1�nI�ߨ�aQv��R}�y�2���].\�O�WC�g|�֫�B����o�J��¥U����bF=��6�J��B*O���|3�m�����n�D��>#hY�Q�tX[�S ��Tʬ�p5���f����Gy����g��k�1��P�����*̾�oR
��w�	��:��I�ss�z@�f��N
��EA����8���"�N$�2q�Qb+�U���(ol:�Y��\����qʠm��L��]<�rtGp�}oBJI{���&�x�ػ`�S��̛I�j�H�
���D`�JQ�S�p����B���*����;T#uAx�����s�b*R|�����d�08���1ru��P@��+	���(eT!R��8TI���t�� �����}Y*��ҽ��N_��ꢸ�b��L���rԦ�7�؟����o1!2�gx�k�U&*����O�,I�<��#j�2�H�$� t�+X��F��]�P�wx��}�_�e���d&�$��V�d|�8}���R� �OED�HG�����[��k��F�f&%��j$�F>��:Ol�\c����������og��@�E�),�)#$h���xm�U��c[�����:������T��Wg[�uz���_�* �����0aS��5���m��H�N����j�p@��d���hY�n���☁�FM_�@��rz�����Y1�'�hyPN03�B�h3R�z2��D��W`7��ԋ6���v�Y�사��RI��: b�����̼��s.�Ѱ��Q�g"�i@�>[��E�t�ӹ_�a-������1���ȔNn�ʱ��X���=��nE��+�Xjн��C������Ox�ߐ�CSDM���z�O�D��s�K��T�*�fJ����,�ώ%xJo|g��D����Fq���ڴ���8�" ���/g����C��+��r5��� O�#G�~?�D���Je��c��PC,d�ځЪ��)�n��� �CZ`ģ��H����O�|m7�jfP�3�.E����}�jB��w�L��h;�";I��x=�U���p � :�M	������M�q��G2=��4>�W��}�L ���+{h�7/�Y�@D˴�c��i���f]�v�J
�}�?���c�侰a�׽��`'��� &���m�[�
�cvɍ��}�bE��O0y8en?j�-����s�"�G�h���q'??�֚9Wŀ��n�����k�Y��{k���N�Kv���6Z���kaS(�Ӊn�PU��b���l{���̈=��' Ɇu�e�:�R�u�;�%P��3:{��<�߹��,���>�I9��O+팮�̼����3Q�2}#��<B��W�����Z�1 �=��@Rf`�{�G�G��7$�<����v���ڥ���(���U���?� �>�YG#0����W�<�2 ���)gl /����ǀY���ɋ��i���ޘ�E���cK�foɈ)& ldb�KA_����ݡ3Ϳf=B?$k��ܑ(�����9@7��0R�1���h�q����6P�LQ�<nm�촙�5� �������C����}�b��p�	�Ar�W�-��"����p��WjF��<G�Wo��1ٺ�V���&�*GDoCRd8�Vڞ�1�=��7��+<�	�60G:�
s���?�Q���,k�*Y[˦������X*EhZ�TMݾ�YVaQ/�3(aj�O$>}�S ����x��AZ��L�R|������
��v7���0�Q�U0�����»�N�r�]��E
�qV�*x�Z^"�������QJ��������Dg �b̙fA�t�L�|X��B�v.��)/�2�Y�h�dRsy?e��H���q���3�v���Y?+�}��j�1q�@ҝ�b���內�(V~��M��m��)��V��G:���%�|�ܾ������ZUQp�֭��v2������ю8��
�G���Ey�s����77���K��R���¼�,a��nN<^u+%�Ȉ��v�G�),����A�!y�����t%�i���%&c'>q&+k��d����WL�6V,#�j�^�O��H����+M»�6F��ޥ����X�'^�{8������0=�9Պ�q��V�T����N<��)�p��=��%�F9?*M7U��Z���CY�N��9k��@oyu%K)��3�4䛰A���m���&N1t��"���z�T㈕:h7��j38��ȴfEd'?���h��}���H��+@��41���m�.��4���J}Mi�TG���i�YX�%�QU�&�
�B#b���Y�VA�;�(@���K	}��m��t��~�}���u�&�˺�T�#Jْ�Ș�#�ň`��1ĭ"i���58��{V��G���~��n�JX���1K~�ԧ�	ؐ��	8]Ç�� ���a�娊�I�W���I1-��͊�ڕ�~���K��wM��\Gm�m<���O�|󦕊B/v,��\Xb���뫵�q�,j1È�u�^:����Ӿ����$�G��g'E%r�P�AӲ�ٕ��!�(��J��F~�	�x$��xa7�Vѣ۸�%"�1@�/�&�m�������_DH���/��:>�"R��+ݠ��S���������jን��S���$��>h��%�q��O���$��{�ޗ�V��)���#;׈K#��eh��ր����ӨͿ
�|K��^2� �}7��w���j����r#US�&� 3��7��ܲھ�/(�i��d[I*=��T��-�~�k�K8l��2\`��bV�>�4�"T޺�:�����"�J4�3�[��l�N �!�vm��3�D8�B��L��=� �9��1�}R{�,���I>z�U_3��	�G��Ҍ*[Ye�̝��c�� �]�o$�ɮ�=eX��/BQ-3b'�g(�ʱ���ɴ٣��W�5�ʹI������.��E߯�S������y�Wݜ����mI��p�$�^���z��P�(������@���t~�0HV25���O�m�%��Q�,��+
�ٹ+x��&M8V�_�X�nX���&�����4G[/��e��s�Ja����6}�Xs;B~ƕާޚ�`eN	��#��s �b�,�5R\2���.\�	��S�K�����(�����؝���aPѕ5͉d�3m���\ހ�/���L����g�+��՜���(��hW]7�mΏ��s<bPO��@*kФֳU�3�mm��<qԿ*�^ԇXV���~w�W�G�Fe����u�=�$�S�.�<a��?���9�<ݭ���A
Fmʑ}�vh|5���8ƹb�����b�����R&ig��2���+�W���\7E`��SS�X�){X��N�㙤q7.0�~��l��M�dxط䙌c=�
�P�(���=;���z��嘠����[�6��������j��NA+��k�xo����cᶜ�N�]|�m5t~+��V��7��%�9wg!�9|��勒/`r�nVH0m[Wa��Y�e"܏���!�L�1����.MC\��>a��5�@�g�ħR�w�;oݑ���	#Cy-��ӫ���~��|{Q������nB��ؕo�R�+����rϭ�|`�8��0/%>u��A��[mCP���������(LS��c��%���xZ��!E�I�jB�U�m����Z�Ǉ)����E�kz_��7\!�>e>-W�����v�:N(>���)�ιU����4��v�p�3�Hd�.=��bB2'MP� .ώ�g��˥����eG��B?�#�����Z��k8�+ ?���
ƌb��Ƒs��p�(ȡ��:�L'x$1�8���Mtqf_����{嗓X.�:��n��y�E죰��S���o��>TM��t���։���ܷP'�N�8��F���h�5RVF��Z֡.���ϢPO���r���x�S`n�Q���/{��(��_����Jxi�H�g��̈��<u'�iV<?�v����1ADqm7~#�o����9T=VU�MrجԬ�� ����S��(^�<򃽢�<��D?���{V�
t�oIZyb�$���]#��<̙)=��Y��x���I��g�RxV�E��y>�>?̀U�|��@�����6K{s��7�\4l�r��8� \��7���_�B�t�;ߠ�1���z��������5���Fq�C���(�����'�Qh��M�I*�	��t��s��K*j8}+�o36|��a��`!�������
7��<�[��8��K�
�=�(a�Iģ�:_���h�E� N��FK����q�����,�,9��z ���~��L��x�-�<�!��9G��r2��m��I��t���D�^'�+��Ldbq/<љ���N�u�g
��p����!�h�d��n��u�m�~C��gLrdE��qR.;�s���L��iQ;4��)O}�JuWY'�!5�)��N�5�'��w72 �*�0g�fبg�n����S���^a�k�ڶ��kR���W)��xg�G�G��9[���I�͌�۵'bcT���ȥ�/ {�o?ɞ�],��U�6O�j�g/�V[�����9n1�D)g������U|�:����s�3?���mW��sX䐘��G	�!��F��1��n��M�a���d$ҶBAB!&���!�Ls���^�����Z�aݟ�s'@���w�Gl����m ,%�g)�{����	1�!u6������B03��W��j����9$���E	9�����A�f��i���������}J��k����1��� �ReyFu��o�+>���f����0$���?�3aGo	���%��d��ua���?�@[��E5r�6Ѵ���a�s�?�����4M�:�������s+x� P���e��a�{��*��e���{� �'������[~h�s�s�cð����ǟ�'�g�s�X6�V�1�� h��ėg-6���ja�����60+�bEF��������!u���Ú�2�"�����,Lx�t��	�
DS#�ǲ���ˏ
Q%'��͊[r]<�KA�b�}i�ơ��j�r+�׸ڌwrKS^���$3ݎR	��0�Τ�����<*n�<S)9z�5�ȉ
��a�vD���#Zw1tK���&��;��̈́�}:�b�q^q�6ԍQI�'A[�bFl|*��݊Q�\���_���n*X-(�J~U��7=eg��ʦY����P.|�:���.�>�'<�S���b8���G�eoA���߿+�,1�+��GL�R�� dx���n�If�m�d�g�ʳ;ž�X/A|���=�s ?>o��Z�����:��u(��v�䳳d�ӂ�ӎ��8%7�o}�C���M��^�����g�M�J�3�6e}Kl�C�*����ſ��4��+m�8?Y]%��'t�"���j���X7)ګ݇�Y���ʺ��7ِ��sczڥ%?�%��2������+!�����I��]զ�S��^�BF��."{�9X�� ���iG��})O��%Z�G=oR�ߑb�J��M|6��K2Kc���2���5Y�������Iޝ��e!�V�-���a��l�Ł��;<}Ck�k�%�Y���h�mjjʵ��ܦ��ďu�Q�Kqg�[%+��7�K���n��g��Bӑ)��j&�|ʷ�m�$��'yp#�
�q��;���nx�Tk�uӸ��L3��HL-�f,]0���B�O*)u�1��j�o�	w�3ʨ�.�紓q�E<5��������q�y�F�{�fy��9����gp��#37�+�E�k��;d�б����j`��ߏ��<K�s(4�[t����{�1�R='������l����9=`��R��S��o�]T{Nd��P
�9�C�g/j�?���"��A�,�n�W�����a\_��򭉕���R
��k���1�F^P{���A肭�� /L�d���j�:[[Gc��%��#�M�ƶ���fco���G�j��Gf����i��
��O����]��J�XJZ�Z�_D8ؗ�������Iy�