��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g﷬#����O����v
p���D�eq��萱5��-1�5;�޿�^��)�!B�̪�#��].� 4�� ON��ZU��+��9v��d.��kjDL���
̚ӑRQo���2���dU���$�R,�Y���"�Ḥ�T�<���:C�/(b5��N�����Oڸߔƃ�1|��e�!o���9Qz�¡	�* ��1_e��H:bx�>����s� �@��q�Q���(�3�3�t��[nwH�t?ev7��T��Rm��X���	%��D&�Y�)o����eV�Ԕ9?Y%R��4��I�
�yNTI��W�Rv�6^�]s���L����	��ѳ�Ar���}b��q]����b��L��Mʏbc��Nh�fS�Q9)���rH�}t��s����U�$��ͳ��8{S�7~@�C�
&%8Z�e2x��"�J���:���vc�,aD�ǂ��� ��R�)�6�nƧ��EV��������g�x�v�ڹ�p�w���u0���ҟ{��V��v״���>x��>y�m�;f�TӯF[hK�)��'��겏�1$,j� ��"R����j�S=�l.CM;w�S,qO��¤{E/Q�����i9�/Z+H�44�	<%�x=أچ2�x���UO�>�cyo_0k,/�q�ϻc��ЗMu��&�]m�S��I�ȟ�t�]$C���5���!xp��y�yer��H1�T�9W]�5Ԃ7(���) ���������Q�w[�O�c���!g4�OV��Χ�J;M.o��/y8:�,�s��-⩽���J���s͸��;�7U���B��KMn�p6�M5]u^|�XܼV4�;R�H�:��N�v�o��hXѯ�躃(/�
�e��0�I0���FL���i�W�ꔌ~}&�?�K6����h�^h�crE�*(f �Mhc�N��̱������ y%�q�d��GrYʓ_6p=L"C'G[���S� ����c��6u
)w@V� 	���$�RR���������!R�zO�����󼄖��Dɗ�j�🩾�⁴�u1݋�r�Y�>�� ���gg�t'Jw��_$@	�O�V�-4�E|�Xo���#&vc5v"Z��i��<h���L��M��6*%c���K�71_ڥ�W�(���;S<����B^C&"�V���K�$���� %ڋ�Q�ȷ9Q�\:AH_��F�J+��v�#\u���`͓�|�6��'A{F��ܺ��Jp0�sN3����:�G���z��{[���"�3)r;If/㕂��#D��ܞoD����:Y�k��B�#	CP1oT�Mhr �� �w�*e!C�9�y�1������`��2,��^�jc�Z���&C���[��w�eA�WF35�0�1C��+�|T*�r�K|m	rQ��Ţ</	P!��x���`��q�rW���-��Z;�b��w��R�����m��Dp�����#���DP��	�*�Kk��V]^}J�)^ư�C��m���������n{t����DdO��~��l1��&�7�>(&��Dia���ٗ�?�[?f����9J��G���;/�����3Z�#�D�92 �%?t�P����&��]鱼��'Z���F4����0�0�v�+
?B��_���&�d,�|�k���z�M�˗{��"?[=����~�Ȼ7^?ҙ+��'���q�3�-!FsH}���"�<F��9�g��������6�O/?�sS�=��ϴ���c�Y#�u�4ΐ�..�}^\�x��)�&�hJ<&���g��LWXV!�bL=���o��݊�=���&ϩ��z�//�U}%KKN�Wi.��v%Js�8Rv�Xժ\y %?��i�3٬e�}�463?җ��&E/B
:5ˆ߮Ԓ�+������!�C��7}�XH8ԥ������" x9���*����n�, ���Zbc�Ͳ���*a%��o���zA�7Y�۲Xրa9��Z���$/��-�h��)�t�W�R�����9|�FCe
��������U�x.���-=���8	|�D�ү�m=�>���;n�t_J�i�qg�k�$�e�B�nE�a*��{0�l|�;�$�T�k@�q�Eのo�%�����Mu�b�JW ��E�Y����?m��~����1xkxݪ^^'{�g�k�&6���U"��i��D����rp�K���	S0t�7G<��ڎ�j��L�����?��z?~`G�I����<3�ޮ�a�2�S}F���ň��4���預��3�u]�	H�7o`�T8�s�ʺ�$o��S��h� �9�7���޹kX�;�ZRU+P�JP�Z<���b!�6��K�t�6haܴA��E�������6��nh�i�gg�⮏כCu��J���e�4�7�H��U�������}F�_
���z�7n[�~b�
?�g�}��^}ȑX�V��$���iu�Ư�*�AZv?{OVHt�Ѓ#~�Wҫ<��{=�����`&�ǳ�@� �ȰY4
��_y�ԼΞR��m���g�vi-�ps��v�j/~�j�Bmmزή�1�/�B���:��+�����i��E�| ���x��	0�놗]��Ϊ�[���'��ϪMK�T*6�_�HQ�Oc�*���1�^{�
o@�?�%Ņ�ڞ�L��I&��������U��*l�5K�8'�/�S�k�*{�{����RP"�P�#���ڈn�.��,Uh������.�c����@��I5s좔����Hܤ~%�_A:��Q(o���`�j/{ձk��{nNˉ�D�>�'Fe��}3�Ƀ�~!��&�f��TJ�{`z�[K�E��Ė*����F��e���	�T�84>m?��ಜK4�uIOY�����j�ʓV��R9D[�;o�n3y�ZϷ4;q�ތ,����@G��-nE�d�~)#B!�2�L2��x�(�g�3��@G����8{��vq�6��Ȅ,��z��Py޴%L+���Ģ�`h��Dw�}�*z�ۻyiDn�:��g'���&'J��d�:�5f:��ИU�"D�WP(�
�P�ŶS:�ߦ��1R܀���*�`"���Zm�l���[[���Y��tM��й�~4��<2��\ߒ��9�I>��I�����J10(�&1�!u$�-p�2>ɝʤ��U���{W=�D����X�+�S)f��p_.��q�M��s��:S����U.a����}U�z��a�	��/m�^�3�T��P�u���թ )-a-�R.�g��vR���<�25\�LRz���7BR����^��n7s�I!��y��j�wl�����>G~ E�]�8�)�K.@���r�=��n��0^�HԢ5��Ey����3�3��͝��n�ԥe	�q#��.��4�6Ƈ�!�f�|��'
�M�m�֭�$�k��:mv=gC�#j~�	�@eM�ѐ@ȏD�m��J8fÔ�*��߮g-����#�+B��gJ�Rѳ6>O� �z��wTK��@��bʘ����H��S*���k�«G`�tN�d2-b�[�~�Ky��$1N]O�#�Y�L�$^�n1F怿p����r�~��7FL-�Q�vq��e -��X�?�/N| f�%�E<�O��� ��b�K��q2�Ĵ� ŗ �V�k���Z	��X��>ɜ�oS��s����f�-mC�[b�G����/�˅��M��:��>?5����·T�$����𓿔f��@��en��1��'m���ʻ��U�'o�б�VÅ"0M���^y�s�c�<&
�R�wדOZ��3t��z���qZ?��B,Y!k��s!ࠛB��K���gځ4�a+�r����gYt�S�t���r/�9ɦ�� #W���[.T��?���LEr�l/x��Q����x�5�F+3ke�����gތ�D�G�����1;\�)��^�hĆU�TI^�~E[�gm1lAe�x���I�\~u�M��em��H�����R��0S�Y��h��2���[�l�5$ɯ��8o'�Egc��+�|��A�ZVt���|�^�&�}�'����4���Oh`�M�P_�٣�+�5k�ō��%ⰫYrP�kP@����(ŧ�b�G(��E��ޕB�Bc-9��AU�u��`͇wY�xP�(f������:��3�~Q_�Ί���p�dR�~^�� ��8*��c�ɇ���]kG�R{�6O�jXd7��t���� ���~3Y��}�$��@���!'�n4\ge)o�!�[V�Q�-n8މ-]�gh=gQx��4�?	M��<�Y��M�I5y�*}���wv�����N�,͆�f����o�l�X(�	U�����~+O��y)��{��w V[^X����/�L�`k�ΊG8&	iuL$�W���k�x�hR��C<��RA����EY�cPA��s�U%�@_u������d�j�-�����z�������ތ��w�Z��&�bH��4�HSԭV�w~�[ s�x��`s+�n<�o�I���_$����q�P
�;�����Z�릏$��Kz� 7+a,J��Ѡ�ɸ/��8n�#?L�~�%�"�.N�9��;��c���k�9�vY�⿒"?>�����pk͘��SA�xO�G,EF����L�f޾[��s�+�@l����\^D\A�(۸�K�LP-}VntmP�j9!e��O�h%#�����?z���K3~����J�{p��ޑ-�K�=�Ԯq>�R�}qrzǱ&Ƈ�V[Y� �$-)��,���'�ΰ�Q��4� ���� ��	о��:� %s2E���mw��)V4V[� �Y�/*�y=�-�q���n�N�k�����.�q�1<�^�t$�u�T |5l�Ư1�]jxb��u���E��ϯg�*v��[R\����U��{{@"��Q�E-�%1�WD@�����8�1Y��.
",���2��N$E7N��iUhN��M=�dau�tӀ^��������ܘ��N �&���`':��;�XbX؛qѪ=�mh�g��0�y)�A��I�ֹ��$��	�!�d͑�^t�nRl���L�V���8I�5 ^����Jl*�O_`AR����9�w)�KS�>dJ=���qa۰�}:�ޘ����R�`����F�4=_r���SO'�OW��\!�'���~����bӅ^�U%{��)��[Q��ĝT=L?d+�l#Q������V�B�u�������&p$�n�6����~�[�����<�E�ل�����]n��y{�²��^bY0���JC������"��D�s����-�~�
m�*R�)o{�s���eZ�4c6�@��CߘdN@��7��_p[�m.�ɍȩ�ڧ&�#0�ϬK��ew�g���F�ve�y½B��}}_��Y�Mw��N�|j�c��$�uQ�M_ �^x�M&���D��JZ7q`�D�nb�����r�+�n��(w� H�R��>R�6 F���t����ݿ�����4��_c�}�ݯĄz��{9�W�WU�5�9���ᣝh�����h�"g�Z�\�d����ӗא�q>F}�q�������#r�D-��CQ�z	�p�}���L�Q7�bH"�dv�D�׊�JTv���Pj~4$q]4�G���$�z�Y�0x.#�L��n�Gň���5CS���XC'ˡ��"%��
y^��e.\���@�JsGQ�\�cE��侷�[�e�Z�D�Fn��hG������m��܌���F��S�ܭ)!n�ٮ�7���%�0�R�Ք&Ӎ��{A��ӳ�q|����w�HM�`L�w���As8g�](�|��ӓ�����wh���8��)�������IC���Ew�}�F�L�A̭�*���S8������+	�[� ��*�{�?Wq�=4)�5���I\](��⤣߇
��H�Û�f|��vp!Jo
�	�}�Q���nfHp�,8̦�f��ٵ�� �k��8��5���m�����A�����е`������A�o�̸E�~> �[��_�����,ǉf�=m�K	沤jf��^����3��A����c;�[�D�7�[�˴������i���ݫϒΗ�m���H���n�Z��6}�`��t�(��d�Ss���%Q�t7F��k���W�st��b_�Vg��|:�#�^�*A,A�U,�E/Zy��#�䖛Jq(9�i$��AX�n}i7��@@��.|-�����
@aN7���w�G+��Xsq��U��67'�|�����k��Sז7�E�wF��cs��^)��Uq�َZ1��x0�"7Y�h{��G[R��#r���џ���<N5���#��c#����B3�����Qzbqal�<~!�m>c,V�~B��C����y���=k�����LwΚ%��K(NU^�/�C�����r��-E�̛�{��"�b+>��>1Y"�p��=�s}Q��I/��,�/$�������|o���� ��SG��!}1���5|$��1���N&��_?�,��'����ޖ�7#��%����?ܷs:��ja��?�=�γ��Qxn5X��o�/���e�k�f�k%=��Z���;��W^oy_q;�	���S�b���m	�,��)�̠](�a�}�_N�|%=aC������y�J D�����B� �^�:�3�Ÿ;���4�0(��^ܼ�O��Y����4<����i���R��̀^ʄ����	���
%,$�	��Pm�Qv}Z��G�ç ��75�J��5K�w~8*�'W�Zkه	��
�#���Poh�k�X���,��j����á&�*|�w��*�b�PG^J��z�N9)ﲶ\�)����u��˵�0��G�c|�;O㈎ɢhuz�ϣ��,�D�S>>,L��nuę�l�L�O)��q�\��p�i@λ�:����w�$���5��f(1�`������ �F�hT��D��m�w<?�WH!e~Ᵹ��\�-��C�U�KEEj��D�4�aP��C�v���	0r���ښ��ΩԽw����������UL��\���f��1�^��*��������ڽV�E@��籦q���9�?�?�W�o��1�>5*�t����1���#<����̭C����ַ6	��$qm^�IB�Nx�̤�h�Kٵvڀ�1wm_����l��W�#�ж9�r������H����:�- շP֡�S:YCL
�Wi���E��.���x�Ҥ�H'����k��$$�B�0�[���
Ǥ�U����5�9���>2<o�C�� �	��#T�T����� ���A���N�� ]X�����%ꥨ���B��ڷm���x1Ȁ�YēYE<���P˖��IO�pQ�ȪQ�ԫ�nR���0����7����*��p 8)XRƵ�uA��C�a�c>�4�J��V�]�T��S}����Ϧ�!��%��{�0�hN��|$�ce�a&�<���qx�*5��!][�|�� �R,:Pu�T���h���l�=`��#I2Ij+�|	{a���K�j�!�1��O�	�)�~z塳.�cq�p���<DN��ց[�؅*G�'Ok��s��iԗp4�[F�╔3�����"�%�''�����'g�h�u���-p.���&:!&8{32�@C��>�)K̀1*�\DJY|"i�B ���1q1�?(��w-U�?�Ih���Pa/N�tS�	�HA�{�O��P�G�.���6�8R�B���U;3�iq�渁�e�ד$7��a���(��\;Hz��<:y%2��J��',��	����h��wF�̽`S�B���І߭�>��@ZEv:u���X��,������w�I(^h�*����)�$>	\��d�����/e B�RX�ǚE�W�MUy�L�;�S����d�6CI=�iDw{>�a���z�"�q��y�]*���(�8I��~�n2 _~�t����`,�o��_�t :JJ�^C����큆�)#�r~�-?�ߛ�����مCn=�Y�����O�^�,�x��|T�3�w�yW�4 r1�{h"��l�TA�R���&o�}//W�O5@0�ಐr�*��/��y���j%�N峼��0���ȿәX�Q�4G�k��~������O�[��ny���8b�R}���,՜�MQ��JE�Zʮ�*�'%-�p��K�n�����R�9�u:刼�L�6(Z�^ۛF����p*��%FX�~���l��of�0\�
�ֈ��N؟hȤ�*3��=o�Т|d��A�Ѕ���l1��=>�C���6�(K�.v�%���M`��z.$ ,M�u��(k���EWI-Y�n�o �����K����s&��b��������ۼ5\xgk}g�,�t�6�[�g*tZD�Y�B?��ΜO"���ڧ�l�;�B5U�Vp�T�|���x���:�aw�<O���dA��)X�+�VU��}�G�g�2p����w����$�v��f��u� E������<�[�n��J�c0f�|Ԇ4m�@Vo/�ØE�
��!{�v��K��k.12l�
��z�r�`ߵ�֭:kf|��S�E��j�w��MW���RC��$i������5
p�O0NG}�Ʋ���/4b���?�(�1��F0@�2J	���8�� A���M@��e���A��~�1`⃌j3>7A��ʹ�.5$�@*�����*�����D�3m]����Vp�}ޛ��ϰ;��[�U{7`��`\��EPPE7!?@�4�2�A�:��xo!�4Pg����d��R����o�+����|����f|�ٲ F�	N-�U^ީ�53��	Ȟ�Oq6#���V��\>|q%=$�q�j�U��{0�\��k����9bAت�Y�ȁF��b/`�m:'Zm.��m��[� ���G�4����2.���"��-�:�jr5$�x4�F?���c}#�L*;J7[K�]�uq,P��C�K��*sh�ˣ�~��Nk�7��4@�*��3�(���	q�
�� t,=��˳�䭾)��iթXib��˭J�\����|S{�|y����A��=��\��hܬL�jֶ��3����.�4֙�d�z�Yt��N��gH�mgҜ	�!�vgd�+l�g���^((�?� M�^�l3xI���k����;S��o@��"�H�@��!�]��Fi"��sN~�0a�X���`��I3"U,�H+j���:�{�*M	�x�:ܺ.� ��&�s��a^uc|����R�Φ�@{�c�if{+~�����9oh����_�L��@�Y�h�$D���F����<���
�7n��7yb
{ϙ����S0�P�/xif�a������GR�'���
�%<sM"K#��G,���݇c(������*hD�9J�, H��I���c��̂N�3�;x9J�BO�Uq%݌�jpt�PF��l�9��Cn�:��h
����Fn@G'q�7�]M����R݄9��⍡u��U�=��߻}����\�����a&�A��31=*�����g%�4;�A$��&@އ��CKC�P�f�?����aS[�	�G�[rl��[C�Ap�!�������������Uz�'*�ʽ��� {�jJ�@� ��/�>Zk5�A���`�h@�3#���gAE�?b�q縓ǈ��Cy�~X�Z�7��Ip�w!Z8�(�'�=�yx�WT������\-�Zo����t?�ڻ�K�P��Ie�~^�J��`�pSǻ�y{s�N$�ul*����e�v��V�P�F�}p��C��X�a_��,��C�$~�D��9T�ޠQ�F����p��&w���\g
q}�}��=�A�J!��W�8�k*�f2�-LazA��$f�.=�n�~ÒiYr��A���D�Z����(����NO��v���0��hr�E21�E	�in��w�h�����ng$	�C:/
ႊ�8(�]�Z���X8������Y4��c8#�a���[����Ψ �$��[���qP�d0a~�`��hՐ���Q$6É���Kt�@2��J����UL��e=]e�Q-��mF�I)�hDi�c������T�P�qKq1`�h`�s#i4=�Jlg���=E���|Ѻ��\�=ő�lv��]�f�L6����TY �t��ewU�&��%�3ozA9��.�7���tܣ+o��z1��1�fg���h�uÊ.u������DQ�u��f"Ĥff2K�D�;�>�R}��y�W���9$g�����g�Z��ݤ�D�F[���Wd��<���V�zY#�K��{Bj(��*�v0M��oU!/|�(<^ީ�O %ځ�G��Q���ߴ�(�6�R�,��J�B�Z��n�j���Q�֌�~,�w�.�!>f�^�̤���z�-����$��c.Z�R OokG�[b�$�M=7�I��$c����ZZ���`�1VQV2����N�ˌ�8 ����=un�ɳ!s�� �AEN@}�S�N7D�ѝ���m��U�63_l���{��U��b�R�6kT�����hR���0$���i��)��஡E��>�b��_5��3w�o�rǎ��|�.���?B����a� R��$���ǞR���k�zun�bCZ-7޴���2�ڜ�<���H��c�Im��e*��<�.L�2���Z������#��\,��`��%�pn�3H#�4��^���7��Ѻ�e*z�b.�R�D�~��M�T���>��5���ŝE���g�<��/M��6�հ����"	u+T�T�b���VI$��PU��/�M/��O:��д7�ݾ��������߾�zh�s-��q�̸�����E�oa����}B�	�yB�� z���~0N7_�>w���qXN��. ����}j[�?xߩ��X�D�~KHL�\AI�2�% /�?��;�t����P$]�~��6Kda!��k�M���{�=	uP�7�0b�'K� ��R��K��frR������3��i���7�Q~0�V{�ÿ�/x �t�ş����U��Rc� �+�������s�� &8�횉�F��-�M ��w���@�܍��'���9�����9,��e�$$��;4I��U@�O�9w��k�V֠��\���r"��o[&�S�����6�G�����)<e������D�A�_�p�͍�k�!��~�QFr������LW���{S�|���u�-n��s���#�sA�x��˪��0�M�fM�Yw����8��vj$1G��� `V�P�ν��&��7��KwJ�X�r;ú�xA�<��2m L���D��1Hw��MiRկ/�����<�޷_8h���I�%C�)�R������k|���:.����:e����Dͫ*
u���w�J�-�{��	��Z�F�a���e�3,�g%IԎR2w
�U�SFR����_B��B��ױ
o��|����8�k��p�&�ȝ-L�`�Ҩ�`g�[l7ۍ�T�� ��A���0��P���� ����~%�%��R��Lہ)��J�/��/�5���<H)��0>���U�#-9���[B�<��1�����|�tD��K�h����v/���:#�Z���=��+G��
)>�D�LL*[���#�!5���<'q�����w9���wwG�J���8�>��)� �ڝ���8��9�$�o������(��.�gk&�UN��=�MY�Q��˨��LӔF9�����ĥ\U��yjk�0�T̧�8W1���d����bN���?��਴o�Qv�w��ZU���\�`u"`3�9=��Mɿ�n2�@����s�8�=�Dc�6�ޟUF�eT��Pu���N�A�SA�!��Ҋ=[G��S<���]E�K��|͔��5��/�g�\9��/���(�c�ے�tmm�����R��/�5%�,$��T%JQ���ϒ$`~�~�އk��%�V�LN�ej�@�����.��܂���"�e�:s�x3��9m�^����Mo2L�~m�iF�"����v�9�o�}h�^�O�G"%��V�*��,�1_�p,l��'��
�4c�q�Bd����/|ڞ�)a�q�d-F)�oÁ���N���Oi�f�)�$5�nܣ��6�k�����/yX��RE��l�
����0v"� 8��H�e.&�[jƘ�:@�<�Q�s)�� �7A�d����LY�AS%�!P����7�.�$��;����@�� ;��4�Th�w����1�˨T�~�].�՘f��.����I���[��S�I'�Ǌ�U�D����Z�$r�ᅀ�i d�|��z|�ڰw�t�q7fxp��@�޻)�q̵kz^7#�֜��UVsd����Α��"��f	 /ſ���[O~Ņg�֥�h��_�޶��
�_ � ���b�h���r9����J:�>�/�꬐��� ���X�ȹ��a��ӝ�Ջ�8"�ll�N�����C�0`�zj7(���_ѹMP`�I�_c1���2x �qF�հӼ�r�	�����`b��g�2&3��C���!x��|�F�{��Ixx
�����o\f:���w�c�����E��*�0���0���V��fe�@���Iq8z
m�l������� �3�Q��Q�a�zЪb#O ��gbY�ՓD�~���m.�&��3���U�m(��	�Wb�,ՎYcA���X^�:�[�����0,���dt��Ȃ\�K�.�K���N􈲭�����%�w����닭R��SZ�R����'c�Z�6�wKb�X�!(\��V���k����Z4�X��m,�O���t\Nz���-0o8i8�U��C������N)#3�:E���G&��oޅ��,�W��:P�^t�_��9ơ�����F���f������q��$�q���'�O�q(X9�l��������k]��F]�M�B`	?-E��A�'&&)�
gҳ��ζv�1-:ƺ�\*�/��t�.�O�ꩌz�YX�/6c,Wح����݈��q�N����avXmZ��_���yO��I�D+�Ɨ[�����@�Q�$h<A���e0�O����l2Zom�#�'����C � H��#$�pc��wf����{�g:4C����z�K����Dce�m��-z�Gl����~��Š�Dy��{�D}��7`�x�����Rqj����t�OQ%0��l��c[��
�"��A��j!��6�,Q/��]D+K�y�t�Ծ��bP �S�un�t����|�[�B�,d�D���,�Y^ʼ��y����M��Q�l����Eb�mo.M���+Ƶ�;	�;�px.�.�R���?���
���ߞ<b��>�!�	�D�j;?���I�\��x��m�X��r�0�
�"�:�(���@��n�6p0h�𣷲�x� q� �(/��kfU>�
F��k$7�G�J��b�QLc���c.�cj[��~M̶ ��Z�[@ǁЌE�\�F������ګ�p���Mg���;���bB�b�o�%s�����3�0ѽ���H.��|6*s�=Z�l��j�#.Wlq �i����Ӎ.ǯ�,XNXp,�OѸ$-2�b�y���_�k9�5T��xs�@-�~�ݟ��9a�m�/���$Whv����P�.�W���
Ws�a.���cP����wf8䱴���W��F+�b�mz����qPQ�`��/��pbW��=8��D���(!���| 6?J3��q�$�m�ht�6V��z�}M�j��
�Xb��F��nJ#�!��ߴ����U�P�{"r+��KR��kɓ���Ū������P}%���������N�:'E���W>Wm����g.?�ȁ#�������t3�J��%�&W�������]����7A�4lM�ӑ���"y#K�צ�:���s���,�}��3a� 6��^�GR�%>����d爒E��'U2��.!]�ʏ�挕i��h����r�=��N�3���g�NC1�m���INh�]���)��V���<���P;zv�_b{����!HV�r��y=��+^��R�T��dZmp�`�7�R"��D
=y����3��O�	��������nA_�BT]x���_�+wL���8����dW؈��l��m�č�Qm�[=HBH�YF����G�e��IA��6��K�T���2�|��eRč�Ht(��]TՌ� �Qf���8[�2]p���9;��y.^Mr/�|��X�y����u7�"h|s}�	��
Hŋ�Z{�1��z�n`]���~���vrj=Ơ(�F�k��:����p�tzKP�P���#������3���X4H\��E+C�|U��>o2�����!Tn��������ըS��֗�{�A�=�� ��$�Up�?v�NC�ˤu��^����9�˱:�ԁ���$���ß�(r耕V�}��"�X��cD��I���Zf�
A9S��^�=��%l6fmH3w���(��:��d� iMSއ�]\��a͛���SL������}��|6�(X�z�e~�$��;���>~>��j�-��x`l�d��ѥ `:1q���$�G�R�SΠ�-�a�d�s��¶z4_���K1�~SD"ꢬ���M<Z����+��]��Lsy�kz�����"�ꅬ�q\���	jz �#�.��D���/:J%��f'/2 �n�SB���F�OE�u�_��Q�͗�#����=W���ǩS�i0ùWz��v��ٛ������r�T��'^mxV�&���L$���D�oYa��NX��!���R����NU�F�/��<�2�)��Hh�
��f���%�����B�=�mG��7��KnOJ��h�O�����,��"�2�As����ij�XN~�����h'H#���Z����l�>�r���*�f ﹭zuA�����Z�d�M�*g��_^����2Ou�O�{��M��ά1�vr�g���4)��<6yӵ��P�h�O�h���:�Q`?f��ą�GuuB8*`�`�r$�JP�ЩL[�Mt�����(V)���j}��Ggrf�� ]�X����#�mI��]x�9�����|cV�l�w��F�Zw6I���f�E��3bE6�I|h �g�^�l�s�ez%8��8�~U���4B��B�K��q�HB���|G$,�K%C�P�IG��+=�K�S5b���{-�5��X���~'����{��|��<�[6�W�*T�a5�-L*9��Z'W�v���`7�ٺ?f5���`r��k��t}�MT�E(� E�Y���w�=��:3��kt���(�Kd��)�>&���)������2/�ݩ�v߲�g�@��U:�� e��t�u�5׀��}�c�du,!��`w�Ҽ�����r�!�����:��lM��3Q9d��}���^޴�D}L�:�_T����Ys?������£b�z]qn$�;�xʋZ��mS��HH���Q�P���y��HɈ����uM��C�iq�o�'��^�eճ�����`X����h����\�o:�`�r�y����?�A��B��(�� �/�|�)���#f�u�����҄l�#��!kWDrh�/�K=a�lk���R�dsW>�߿پ�l�T(����u����u0��pg����W��7��ȡj?�� 쫝�*���8�RH�������W���̗A�"7�吵Xc+��YR�;_�/rIfY6��'Y�q	 '0%�R�끷H!�Bm��Oh��o	�~to�3J����{5c_���Z#CvC�\��(/֥�)m9NJ�v?�s�f���R�*A��8�a�v��/���I�Ȕ���#��C&�j��$�2���'!���Z���N�̀�>��x�	�e�!�|ȓ@/�d��N`'~��i�PQmCǇ�6�b��V��=�����(SӦ�G�U��������ߏ�_���/���8U�wg��U�PH�f�f0%k4��p��3�G���z<.!=K��WF(և(=Y���� ^�sb��΅8�W���<�c9�w�]�-M���+�V�:#�?��R΀J�}ʝ�c �=���C����k�/�A:������މ�I������7T�{����V��3u�3+�`���&����{!/�эB;xw)�O�EP8tp�R4����6]�� ?[/Zk��{���d�61�@\=�um;�X�c Ӄl����M����V�;CI|�UW�{3m�N���4W|�?��z@" �Z����i`�4i�����q�B��l��	x�9;��N(�'�4����ݐ�J$�ӁF�͞��`���Adb�g���gޗ�t|ud���h}�����-K�wWU���_'.NÊ�/ZNmE'�5���$��bX���~n!i�)�e� �8t)�|y5���D��!eu��ݩ'b����9+���Q\����n^�o ������t�f^ia�U�8�Am�j��AW��sʚ��#�q]�����m0���'��sR�蟂�� ��6�`��D>�r
��oS�n/�@c'�]��$$�b��k�$���j,J�[`3+�CR1�珶��>�ߪ�)�hn����)�I��%]�B k�L��ش��T�ǚd�5�:J���.7
�aNf�u8,�N�3a�6�|m���&��|W�={3�}�r(ĐY���Fsp-�38r��L�[/��䁢f�o	!�S�=����]��N�g��5��a��Y��ˏQk�O�4ieK9pp�l<{���H�:2�)��ǧM��7˶[-"ЎM�N���q1�0n2{2����Rb����˵��\�>���m!``��F)���B-�d,]��:K$q��[��21;��P����sN���?4(�=���H���.m�rb����W|@_�|�_|��'GE�p[��=0dL׎<VV*�\�R�77*K��݇b{il ��+M�Mc���'`�y��7jv�o��z���u���9/3@���^xkY�8�?a�~ �B�C`��2�q���` [@����Z�鶲��хD��1Mϸ�*+	v�����2����^�O&i�� ��Tq�6�(4�!�N��5?��gƅ� ���b$��v�p��aQ|2v�@�a�h�9�Y`?��M�0��`؏�z$�������c�>Ovn*�� QM�J�m�AR�Pm��5�U�l�\�k��ݹ��#�U��?�q�;�����2R.���;�B�xM�<p����
�>��ı.�l���Ȫ0+q�*]l���({�\j�d�#�������b�XfZǬbO+]3N3�T���l^4F�˳6Ų<���O丽)�/�5�^=�ab�3Z8K0K��z9�������x��Of�@�*��th��N�����!��e�R:S�$���H��JP�M�s���4��tE��׈��)�ؤ�#���+5E�iDW^;�Ѓ��ё��T���������}���g1<�zI^�o�;�V@d�����rjr��MP�`a�DN��A��	ŕ�F��.�|4Q%~���%�5,S�D5pIք�� ����*RÕ�N������-�G�|��)��&r�����ta�'�:�h��R�h�ϸ�}5��Q'X��Ķ�l|��gA�E���|�Fg�
�`^K�<��-�y8���V�tg
K��0�N��ʫi7\�"�gqxW�a�s��f�Ƿk��|�"��_��6EQC^p��_ ��E�J�
���u�Vm��E��XӲ\�h�������h#�9)��%_$���R!'�IV�e�=��ۼ����`�ɵ��ā�Hp���]�0*��X��e�����d�.��Ӕ��a�/�J�R�:R���IJ���H��FCJA'�lQb'�8����O���r}Q��x�~��)�P��p8���e�r/��-�����޴�8�kQ�5W��{� �>�,ܻ�>lw��$%�������GN�#�l{:����&;P|v��!�NΌ�w>ضb}��y?"� �E̍��Θ���t�Mhzޗ[����H�M���HW�Wn����hX(,�'���� �1t���si�%�"���)�����s�$���!�:K���eo��!��1� }2ak	�6��L�&J^	f%�
pN�&"�K�2���e����xhnod�dISx��>P�S�v�lY���k�R���F(Ј��r&z�#�5t�5k�!n�zk(�٘�T%k3�J��7u���jRU�:24 �PA���@�9�L����8�8fw��Ƀ&�ЈЪ�i�a���F��^��������)w���ȏ��%����v%U1����u\�`ꦅE��7������Q��������v�
��?�XA���p�+{�\6o��]P�
�M4�RU��]� _z"_���i���������`�e{T7�_<���P����M��v̻�łg:�ᨮ��
��v��=�����ǌ����_bL�FNT� P��[4���-��~�aP���,�z_�ä^bN\3Ы\F� ��3.�b�
�(� �Cf�==����4%�I|��K�|ڪI�^mט��V�s�&��%��C��%6�b��3@^m2��~O:VE�uе@�_�lZ`4�Ͻ�����A�a����?��΍�����V(UQW8P-���#a�<��gi4��s��r3�]$�ڇ�lo������ا�Eb�'2��!\y�m�2�|y3����b�$��3R�N�I�c�ޜ�:���C����o[�$��;`>e�نL,�9�E��pC���U��`��#K�$-˃��z�X�A�f��˾�!=����ҝ�%x��k�$�ڃy�zj��