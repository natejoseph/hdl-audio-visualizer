��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�j*Ɔ�r��ӒO��m���=�0��V(��֑^����#0@��{1��PT�A0+E����J��T����qv3/N'��
R��`�pVv��9@٣b�o7y�k��1G��"Q	q'I#u�]�H��8��2���ѵnv��#9�j?]$�(�z�O!(H ��k�a����(�V@A5<~�	������2��g�l
��2�㵝b�8����̟8������(O�bM��jܡr���i�|���(%�,W�9C���;)3_!(@�Ye1|zty����n����0�b���,T��H�CtS� ���Jt������u��P��+�&0����ԞO��C���}�G�cp���㸙[$wwr��q|�a�z�c��O�"��6�t�MQ��8��p~���Y3�s\�6��1�+P�3/�Ǘ��9f���}u®�>�YAY�-��b�l���^N}�k�j�����Gf�s(;_]�N^�<
��QO������~$�2��RYY���&5'1��!؝6�d`��@3��F�����E�u��Z����>���~$���?�2���5X%����{x �N+���<!@ݡtIς[Z<�e��,T�#7,G�Ӱ��M�"mo���,b=Q�^��2�^��&sCpLW�{
�$߹ʦs�EaOD �+�@��[ڸ`���ƞ�:EFZ�8,���}�u#��ޥ�� mg���	��&���Ut'���QF�Oc�����\W���h�(���l{t�QP̹�����PEw�[s5�#�Q,輥�k��p�����îzg�w�N��#��YD�f�a՘%3���䥔3���ֳ�מ�@�}�����W�& &]��TS-�s���0�O�Jj^��)R�X(��N��F�j�]�6�=�f8�^&4��=k8D)}f��vm鋏�D/�����R��L"�%W��m�ǩ��I7�KyJ�J�ϘC�h��	5)�X&� ���J�9�@{_�xǽ�r�R{��}��Q�M��IR-eT�����$��%��+�p��I���d�b,�?�G'/Z�ba=7��k�7}��}����*��lצJ7�WUx��xI�I�vC�z*��LZl��6tBzN�3~���U��g���52�-��������`��o��ő0ҝ_���w�]i��,�'/�+�d�xb�\ 8�h�ZZ ���a�����u�|�.{8���������"�d�5'��v7����E�`x����Ut�fɱ�mJ�)��9i:�K�"R�0���L�����"��y���:uS}�w ���m�V��c�^X�ك���6�d'd����4�l6�*�b8i�,m�%�*����Yh�ۿ	˴����fVSY85��ƭ#h̸��[����	ˡ�aj�����	U7nZ ����͘���
����딆)^���U����� ݒ��]�d"�B����,R���H�������V��},&.���ԟ+����T
T2��rg�e:�4�=�D��:�Q�0��(�����W��1�ߴX
<�� Ǫ���yyO�l+���	�o�%ڕ<��Fwyͱ/>+�6�n�=���6��q�V\D��d�>CѺ�e��~�r��&8('����RFƞ��xC�QM�Y�O�f�M��je9ؐ�������'?֛r۝A�k-J��9��rf�d����P�9�Yס� ����E��tv��g<� �
r�N�{ǒ|���.�sl���9����4�#�A�U�N�.z|�t��Sl�f���5�F���-���  ��E��t�~*� �����g"�O����6r��9�YB��`w��X�����4FtT~zժ�p_��0c���M�)>��tđ)(��*�<�\��B������UV����)mAgv��-�:����E*��0S�M��">cG$�I�n��0���wG�!Zx��}�E�㓛9F���J�+֜�ݗ��i��ߍ�����,1_�r):[([%z8�Ϻ&����|�T;d���'?1�J�S��!�^%��H,��}���q��/*��0i��.���&.!aH�!���U�qv��Q�`G�0i4�5�C��ō��x���4��L���p�$JH��]�u]�a�;0�2�.�~^q�4l��T�i�@�o���֐z@�@:�DX�����ʄu(t���7�m�'e��@�\J�e�(��y�Qb�]`=�	�r�Zh!zL�{��2�=-��=�Ƹ��5�e@gn��l����&,W�X75��k}����=Bq[Dh�M��:s�dD'Z7-�$�	Eo��py0V���+��1�I�!;�"���@�Fh���dT9�S~��D~���W��
g/����שCq����ؕP1��Ц���U^ f�&�Iq�N�+Q!Z�D�Ɯn�8��������Ӿ��g�����,0G��~�˭�ʨ�	F�B���?��Q<&��= .|Rŉ�Q�z��h��كU�f^�����7�&C)y�͜/���j`֌asI����a�ǩ�OU'���|5 Bd&gl�4�
�<a���!=N�1G|ڃh� .���h@�Ɨx�Y�7�os;s�0���]F��>��W�|�g~5`N��"��`��� F���E��E4����\�1u?��6u��'�n�5W�W
�Z:y����e��Y��6�w�s�鐂N�l�F�9!E���~h5��a�Ҭ�-|_��t�X�?�i�#���t���!�r�Z���Z����cgh����)hId��gD�h��)L� M�$a�B�x�Y�u�Z��{v�V������t��]���r{HcE�=F���Ey\�6D���ˮdr2U8Z'4�i1n�3PN���)7�ݱc]�;���uE:#�3jlZ�=�(-zפ3F��J-L��� B=�@�D��wO�~���S�������CEn�U:R�� �A�G6j������-�}Z6�G�y)��y�*Dc��w �U��AD6E�5��9�<���˃=��o{#L���)���y���Ȟ�\n#
�qk�V���G!s9r8�h�p���a$���(���DtX[3G�>(��(A�"�Da�Ҭ�t~��8���P>0�c�tBw�#����nd�����T��4�ԥ	����jM����Χp;���.���!O��W�%��fž�����Z�$[�(G�W���E	i�L�@��-D!p�	+�=u;H$�7"�<�|a��sƉ�b������U�Vc6N�D�!�[�(�k� +�{�ǋ#��m���W�5�"~˚�5��u���B���	%�^G/�<Ԍ�_�6nLަ��
�7�
��T�$�昉ВiaMW�����9x�0�f�h����.�����k�AG6���4�T@��/��Z�I�8W1������)_:�R���"���������K�s��Z2���Z�����*P�λ�w:X�T~
��ր����4�I-K�;�;t�XHZ� k�l=����y���W� S�`�Am�_�- �H���Xc�"���� 'K��t��Ov�: ��↚���ZA��Hx|O�����"BO��]x/o��/c�p�������T����v�)!!�I�C��s����:oV�d�S|��Z8�޶�N�r<�~�M���K*��.��N"�n��L/(� �����&�+1������s�<fP�4�lJ���65н��]��B�8�`�#�mN ����õ�̿��z ��a͆
�23Ͻ�:z�r�u��B
�D�'M8�R����Y�;^`h� w�s�8 ��X��O���U��/�y) u4��&�?=�X�t�B5��"�43PWK����y9�꿹�	�p�9̻��V�L
�pg_m��{:���t��`^�����ν��lt��%�]�{qr����L�t7��5_K��6���Hq��kw�1�rlH,et�ӷ��j{{��L��.���$U����<4�
��$���s^�p:�v�s���j��4�{vל�t�������K��U�r�@�$aM&t�Q��գ�����$#����?���ƺ��q�eO����i��͋���ە��1?y�|V���Y�ߕX�����Ԏ�<�D�nהN_�5dJyRGD�ɠZ�f��蓭3������6\	��9�\]�4P�94`�g]��8�<Ŋ_L���8�<FnZ;�\In�U�����3
0���l�)n����>O�Ǔ��y��w�TMk��	�aҍ���n1�.&n
î��� ���䛳6��MM��`�ߜ���Zn~ID�tV����j*�:G:��XH�t���0m)��~����jB�B�k[.�"A;�{��J��CT����!������nܟfK>C&�n�2�cX�;#�1�̖�3KW��O/��!r�i����?G�_�����h��m���qN������1��0G��0�[\b����!D��W��C͔)G)RZ��g54��RX�㪬�D!�䃛	�� ��̃���,��j��z�ż�S-�؛�s;L�]!u
0����(k
$>��\*f���G���1W��x�@~���LA�(t�?j�v�QsE���xeF.��
����H<�{YPfV�b�Z���Ɍ�����^ �q��љ� �+�H�f4��6��t��M�V��LK=��iR�<�Kӻ�U�Ts��{���S��쇈՝��Zw�(��f=�&ޭ+8�����e���k��<P\�%�����E5Ɏ��nb�qNb8��JBW��'<Al��A�q�$�*��Y�*�(F� �U�� �B�����˽��G?f�H�\��sn�#�cĝ"N87���v>98F��� P�FwQ���{�!IwI������l����i_B�N����pt�����x�_Q�3��a����ݤQ9�]�u��/��
���lŊ���L�蔲�ᤈ+��	r�>4!Y�˕Yn!Zq5`�'��3H���u��Yb���e�r�x+�o"��룢��֨8O�H��+(. ���b9p���B��iWsqߜ��Z�@��~a�9�B\?&�����ԭ�H�LR<Me�U2F�M����iwp[�-ʭ���Sǒ�*e8'���CMɏ��E���C��4��bS�U���jS�{���r9�k{����4�l�O���c(����+���_(~n{�	 ���ܝX��=��F4���x��6~�ͺ�Yw^c�h�`���^�a��/74�x]C���+��4\HN�ߋ��v�F�v�ײ�c��,�0�BUk�yM�t�C�g5p�Qt� �~h���rd3�����g�ؘ��70:54a[��E5�@��D�ƞnW�S���6��v������Ж�l��Z��oA��#`I�>z�xn��U��b�^�,��p~�}ž��da�C��Y�{�~כ$9hP����Z�K�:��Z�Sm��A����0��<E��W	�8z�_��Ph�U쭸��BsW�?��HY�(�̐�(��|���%%��M�x����Ȟ�[�덪�H���@�޻65R�x�e�Ϸ��x�Bx�� �i9�����w��k1@�x3�!���#*8����H�}>��­��f���aAx�Z51�RN2\�F�[,�9���|�VYQ� j��s@�� ����n�?hk]NM��<O}'�_�Gyg07)���rk�B%��f�[�<cC�\_8����)`W������0��"�����9�Q�6Nz�I'�F`D��ѯw�y�P�:#�E��o	�O2���*�<9<�Y&�ܸ�w�R���*ew3:��d�19��|�9���]L�p�T@�,$�P$*�zZ�1H�X��u��0�0	ٺMpCU�٧�HJ�v~��,���ZS²U|�I��u4���Z��שo�l�^�6E5_H��8ΰ��K��u:�J.�����h��?���Õ�������V~��Cq����\4��]E(�<�����qr�� P�R�?�dC_��"R�W��85�����m����@��^�Q�	���f�\e?Iw����ۣڵ�Ҁ6����1��8����V��\�\�,JZO��2:�0�Nk4r���ҿ&v�w�E�ŷ�@�Օ���j�~��O"y���Z0������\!trН�fJb�I�X��V�xYbPIm�p�V��~U0m�	t܈��M��hC]�Rԙ>��}ܪ1�I[ڟ�Bx�a]�M����8L�Gd�AT8Q����� �=rJ��NwY>̍��'!DX]����2�3���F���XQ�)�	~}wr��?j����;\�qegի��'��0?W)�����Mi.��X3L�c����{����»:���E��l�7��H=?���
4��1�:��kѠ��d��y����apV:S)��l��)9U������d-R�\I ��ak�k�)��$!�Y���L�!p/L�`�,m���E���g���;Qm/l۰���ߢ)*�wqh�2�qɩ8#�~m�n�I�}B\�{��7�#�^��fP��a�V%̦�?k�������k�v�z�����U�KL���I"i���$!]EU�!кJ��ޢ�ˁ���)/�}M�N��u��:G��ҡ����ޱ�oP�a_��*c5�}e���[�g���o�����}&�%zU��y�����"�ް�z�p�ތ���c�����N���4S�
�}�
��g��dʾc�p��w:Ǧ yG��/#�S�;ԡ�1c�Еg�C���/�B�{揺�x���.���z�#K�T���tZ�v��!�F9%�� l~�x6�����+޳��!w�M�S��~=�UMnk=w�&���s�,Â=�/���Ĥ�1�\<Dp�<|^<1�H2	˯�ԯ+��C�J־Τ]�is�_)�����y�-Ǟ_A��܄6����h*P�K�t�N�y��Si�Y�C��Z��5���9Ǖ�����4�-�� t��wGX>�����#��âo�=%0�r�.JuAտ���3�P�E8m�{!	䀀T/vXO����}���o�-��A�+WNݕ8q�nܥז}(��	�\ ���c����bߩ��#�V7���T%:I aB�b[��Y���{�	�r��i���7A]��5�v�������i�F�kڨE�����BB���>Jݳ^�%���� ��6:7�h�fNp�h� ����9Z�Q�yq���#,�
�2k��w6ԩ���:�h�B������o`�&X�
�6BB�ٳ/����y/ vp�8;��M"tՍ�2G�A�!G�S �?KCV�b���GACjAD$��/G�D�NU��G�Ǽ&9[����mה�kPƆ̟Xl�U�}���먮���=�s�@a��D��h�O�sPpm��u�3kSU�<��\��V���Cg�>�����)�z4��	@@�	&��x�E �`Q��撕!AA�W��(ZЭ*����b�vV �͹�`Q:S��8&���\�Ծ�t:�Z^�k<��\)ؒ0�� ��j��b�"���u�Δ�E�Y��;���ABD��jeݙ��c0>p��.���c�OƊ�*i�ĭ�W��/	;���\7���G/T�B�K���d��'߀���G��������!T��ǻ��j�3vɂ�N�ڀ����F��#y&^!WH5B�hB삻����/���l�'�k�jsQuǀ�{��0��IR]�����p`(�R�_u�B�We!mW-�x1������GE_/�^��Q!������������h�Kv
�� ki��Y�(�6ٰH����5^`	�/��d��x�٫�]vC�;�Nq����5����OҞ�HeVݜŞ*��ad(":�5H������D���g�'��n�Q5���r5d��Õ�����܊��)���f�ʭ滣�s��W:�3^-��#3lubb�Z� �c�g��]�dq��7�	��rV�rC����@ �^���w��<|J�����<;��~��6�E.Ri����;�=�2la��+D ���@��:FY�L92y-s��j?a�����P���XGe�J#Q9�����}N:h�����N���3������ �b�m�!����|HH�g�Q��F��7�9��/�C)��f�����L�`;��Mo|3`�Čz�wE���xγ^;i*�ʮ@9��{��Re�e�E�uٖ���)�'��8���4�>�`J}@~LAU��<�@O�����������'(�X]��>��y���R~"�K�s�+��!������J&x�K�GN�p��uj�=CXrh ��c����"�sTBu�<�
�^�E>���.�� a�ULF��"��V�a8�����kM�]�ܪ�A.��`�$�	dR�9�}z`Q�����;}��ݿle�j�2fC�(��RP�K��*z�1�
��!�����2$�m�C�-����o�Q!� �x�U�8?=�;GF|7�Xܕ9��,��)�QBQ���	��5�4�S)�LzD\��Dy�U�[���X]Ct�bX��X*������i!�?��;���-�K dޛ�&;k��SŎQ�c���@�eAC�֔�l�S�ǅ�)#�V?F�WH�,U����C%F,c�i��̆��@o6���mFǭI@k��s��v�+������_��KN��<������5�0�h�=����LuF#v��x�b'=���s2��������D6��c�d�VtU��֕fs�8B$;]c�n��%GJi�$�������]_��q*b��m�#
\"��+]ڰ�6�!Ż���?�&Ż�Fq�^�N�1��d҇Q�I3�������~^K�2b���E��`���1#�/�}E��oS�s�/�D'a/����7W�ҕ}ĸK��M�G靬_�{�r	$Ln9kc�)�靵P"yw(u�& 	�)l��Ҁd���j(�@���M����}�����~�A�_8y�o]���p�HBA��j'���G���.i�CT�R,�qj���0����DQ$�aZ@)�=�t� Kql<�[A��ɮ_^�Ug�2j4ɪ�7bQǫ"�g�W�L������w-
��w�4��b�A.�s���Z�&B��!��5c;�Z<,�3�,�፥A��X��Z9�xKd�\�4b��$�xE���o�<�[��<MA,��������j�,V�u�H�!f��C\���>��{W�t�.}�>�	x\#��F���;��d!�`}��N�:�S.VVH0� m%`����<N_��d��	*P[�A�L�e�p����kmJl�+�����#�*Cf$��N{��[hz��bD�+���<����i��_�h0�ZF��ݦv�ϻ��0$FQ2C|��K,����<D|���'����8��_����nO�ľA��#��6�C��{6�'�2,N���6;���K���61\΃uB��B�Tf�/M�����|ތ��M Me�Kv�7�J��yui��z9�h�E�OF���Y����r����ԕ��J��@��?x����\;�q�wF�ō(�<؂g�P(��((����E)Io�/���b��jr��;�1�r�|s�L_����$(��9�J˵S�g��^i��[�O0��Q#����^&���8���S�@{Y���N������G���P�D'+G�-p5ڙz�g�H���r�>yf�N��f�i���H^���tG��S�>���?r�p����$�4g���멭Z����vg�%Y"���ʡӄ�`'��Z��\�'�Z�=�1��C����:���9O~���y���6���w�[�� Pf
)u���0ޒ�#m>ą]���?�(Eh��?Pg;�����(��jnd�h�R,�z@Xq���k�7(�lD+[t(�X�aĉ7��߸۱�Z�Z���F���a�s�`�w2-����_����T&[���x���r	�~TaA���(�#�5�y�<��9Z�͆�%�_-}�=9�n�b�50���3���Ӛ��o�0ڛ0��{�(n���q,x+�6���"��{'s�7�G��?�|T�6#�a���@3���[�RyB�����2�,r'~So%��/k�h��+��/WĲ�w̷��[Vi���ah�)U`:�Ӌ�t������*�E��']����#��a�X����h��%NL!��vO'�L$Ŀ>�{X�o�~�D��s  j��xN�¯�r>v�G8?M�,�1"�o��+*�-�u�k��b�Sɱ%T*3���}�	ނb�z��'���#5n�[�ֽ�a����y(<�p7�4�b^AAU��6c�?��]%`�C������`T�L�oI������r��U{T#�cF>V� JI���#}�ho��M{�<D)����~�av�:=a��*��vA�ܗ����Uͥ�q��{^�}�p�І<��l�C�
��,���|�@�R@���Q�#��+��%��SB�[b�<�j.2�GL��m�[7Dml�Z��j���K
=�J���M��p�@���'�� ���O��e�;�c�`)6e���ˎ�2�2s��c�f|�9i�x�����#E�K�8S��K�1H�gA��>6m-56��P�);~�л����1�.��-8�Ǒ��v��	KSј'����">�6��r����"5���j�.��%Nc΄5<4�@@���;*�H�;����J�d���O��zO�2E�����Q��j�0�^j�1J��i�@�d�Yí!2����0	��O��k�ٳҌ��u��hۋ>����^���d��C��D'�J�4�r����.������Xʀ�Pq�����v����Q�9�h�=:2�\���r� =>. �2#�n�i�h��x�[��w�ߔ�=�����c��[��-��<�;Om?�gd�� ,�y����X�1�O�~�˄�I ���r�;�O�=������c�r'a�� ��1O?ـ��:jᰛ�`Q'�X�_L����(�|�+�KaД�ҡ(�gH�R���o���&��zN��ehɰ�N�K��N�Y�F�MS�ՙ��[����Gl��> �ND+�,ĭCH�La��G�v�F ƫ�E�,�����j4?k����3�
���N������S��?����'jx����*�	B�ZC�n+��"��!�@���@�>MZ�sM�{H��%�QV2j�`0���eP�I`��+*�N�vO<���ChhB���"v���K��a��b�������T�S�{�S��;�E�_��+ņ�k���DF.!�ts���������� ��w�G�2B�QL�I���=���:/�T��`Z+Ĭ��{�$�XddD�l� Q�vz�W����jT�o��%��Z/�4�*�,I�;Oˊ�q�9w#J�E�3p�ώ4 �z�2TdM�F���'���Wa�=$��%�n���C��d�JL�V�>�.vf����މNmT��~��_+9ɷ��J�"�����Џ�F���B}����v�O
�C���%��LW��%qCP���J=����cw�`<lEу����1��ȹ��0��D@;_��j��*X�\ljcD�c����2;��b~��|�fVF8�����Mp�n-�!�������m�3�F�	>�U�h��TLq�D��Hۑ��1�F�<����������7�Q�wS�y��+�66�C�a����1������QEN�O��&��-���oS&1?v�m� �f2�hXy��RUL��KN�{(5�!ܓ6�&폤��L�;Y䞎����8�B�}�<����.�7=/ԅ�Qf}�}�z9PyC<�j��$%Ӟޥ�Z,}*g�x7�7�ϵ��������y���K�]z���^y��fܠ���"F/,V��K.M�X��A��z�Wϔ���y�Ǯ���}Zk�3`�7#�I~ȥ��D�\K�Sh�A^0a�?��"-<�*��|~0H�J;�?�W��9�q�n_B�-n����ƼT�M�l2:�2PGa���(�籌��kR ��<��ɸ�k�`Y!B�dx���R]�$���=1qs/�Y��� ��/�̛]�*��P`lg�C�Ę��-����0p֚b�H�K�I �W�V������	m�� ���/3gG�+��3����'ɓl����}�.��|ss�N��+9�+�>�Ho��a���Ƣ����"&e?����~��8g�;ެ���n�[p�b�A��GĤD�pĭBD0X&�mE{�Lq� �wԸ���{�h�ݔT�G#�|���eْ�d�ITl��0���б�b���H$�Xu����S���ev1/�� T�Cj�TT��u�r�@dT�z��Jex!7bgj<�6�޿��; $S����!7��暲�x�IxX<��0�z��f�\��9_��Wg.�Gf�z!�3O��b{�������,q}\��[(���¼kT��:>7&�A����.�͐UgD����8�~z|_����;�#l(px��p-��@�o?�����-�`�_7����u]�C,>k���}�љ6k�+O�*��hl�����C�E�C�/���%������5�w�-:���Hգ_�;�8�3��^��}yt7#F�__��XZr����J�S��nb4��$��^j!c�*>����I��v,�0
�#�l:�?��i���O�[Ѹ^ Zg�Ʃ�=rXd~��FL\~?���E�u� s�^$\w�զj�ĕ%98�����S�a����M��pa�N^ߠ��D0��<�J:�β?M�L�5��,E��/V�m;W���M9��n��yk��Y�E�5�d?Qv�w�x�c��p��jb���g9��&���^\E�$]	���� qA��%y��;-���no��F򕋌�cKkU�� .�zzf�A��גf���+X?�^�V�%����_~�_���ц�,�����+n��q���oG�z����6-�j�L����15*�,�r��h�S�1E<�i��j�Z� ցT����0�R��=�өFs����j��96���@?m՛�V�����ś�޲|'ֿs�E2�QR��P1��������9��ByB*8�6�U�`(��p��j�;&���S�9m[F��`z@ˈ,�cp�Ǌ��y?�c�G]�ƚJ��Y
f�����}���=giGP���������PD9���* ��4���S��PZ�]��������r��d>k���w/��-֩Ζb��G�1qՄAU���Z!�K�Χ������[,��Pa"���/�Ǫk�����^!������0`_~8�JV�B�li����6��Pa:�scwm	�=ޅ�\����P���+���O��p?ϝv����:q��-\��HB7a���J�w�bm��E@PI�2�X�[�?�Se���X~{�_�>�(tl��
e�uv�U`�oJ��%mo��S�x�o�x6�(�m)�:V���K��P��]t� JC�`z�����ғb?&Fi<�PU[r�5��g0�����c*�;��������>|�cSWu �ͨ�tD�O^a� ��05I)�����x�aοM���x��rGZ-���������'J�w4Q����FK���Z��Y��+�A�07tR��c�t������p���m��+:jm�O��D����N�K�V��S)!�2�����d7�2�i��Vy�ɱZ�ӂ��Lə6��I�}����7�rh�:�K��T3�y6A�<Wkz�S+���͎����p�h���E� �U���� �f��[�w�8�̝̭�q�i�!�0ۮਜ�-����Q�M+f��$~T0��:�,�)�"�6���~�D%�2��4R�:xr�֥z��cƚ�w}�4�.�P��l=d��mE��T�<v'8Ap/,����9��3�y��gx،�xs	�;����~���$g��(|
��
�6.ɜ�X��n�P�GT��)/}��Gp��a�1:Ή�I������D(�e�к_������b�\���9w�Y1�L�)I�#`M��4�k�|��Xs�Q�9����s�֤��A�~����F��W �
*�`�k3]�KLyܱ�Jg��Pe�8BH��F�i���@%�����j*O(q3������^����`;�L;\FϷ������R��I�|�g4P��+����[5c�.��IY��s�O��=9<��8�7�t�n��/�d����-��ʞo*n�f�
9�l��w�({�������t��cM�
N:���z�.da��z�lQ軬����m������뮲���8�F�0Y��ۅ�I�:���Y�f�Q�#�|uε�x�MI`�uZ�X�fz*�<V'�./b�aa���Kq.��mwt9rf�hːHFo�1����a�����H"�~��f}O�׎r^'Q�*��Ϥ��
��B+i���A5X�:dq~,��g2���=t2v�t��mG�!�HU�	���p���`�d���jx����ۘF����+0�$�p��#���M>j��cTɔz;݅��U'�^��ߚQ؄v�����f-R�Usbiw<����2�GIo����݅�C��!r�,��0�`��(����D���B�tz�w+�^�;cfC��Qs��jCn}x*����B�����E��m�����#�F6�t���'ź�!�w%E�F>X��p�qC|�)x$���?�I�A�<n�4�Z�^�])�Y8���D���d>���S�zOHX�����B�Ԥ�sv);%�;��~����#��Q��acY��+���N��Sc�J��m���w��q�aF�sa���f�Q?Vӽ��~���獅��q��i^��_�Ȣ��L$B�>!���΅Lsg|ɔwwL�|���V�Lÿ:��5���	2bG��U5
d ��� ;s7�v�;���-�窜�k[/�4���l�? t����,A���d���`➴�V_��������o7�w�s��|w���[��>4���i�����Qlg�ܛ|{����O(=`�5O���V��lL��Yb�����R���1�r�Dh�~9���6�,b<�+Z�:"ƻ�ʳǊi���#��&�~3�{��6����&�l͘Dpi�F�lNԡ�)��H�4���i��#��RV܇.�������p���������uo��;��H]T�#d����_~!�#�lDB�+s>�@O�nК�{,�H~o�~[�=o�����.&V���Se��y��@�VZw0w˃���_��[1'�O�TҾ͹&��>�~ގ���Z�f���K6_i忹��ԭ����0=��}9J���K���N1�Η��X�&�߿�oe(�/��\
���Ź��-���Nc��Ş�#�����"Z����k����64g\ߖ7r�x	@
#!&�,�uW��:
�w���*������!h��o�An> �!�"'���޼o����)��I[U��&����Vs�H�Ǩ&4-�����9��i�������G��G?���� ���PM��v�;J�f��?��b�_���/i�X��p����t�ϡH�J�����~K��m��I�o�D����{�b{~@D���S/�0s��T�	0��/	I��~����Y ���CR��T$%}w���F~ǡ�et2�B`.���*{w�� ���x`� ���� k"�r3`���m�!b'#���js���g�4[�q��'��5�[�b��2��]X�D�C�K�Y�����$�y0p��Q#���AA�^Bc����C輬�H��i�*�$��;r�o�0*���M'<J�]�������@.��� 2��7��k�����SZ{_��� a0���d�J$��Clm�nʙvgE�s��?(0�-Z\�:"^�k��7n'_��!��.���p�-3(�R12
fX[H<�B��n��=�xBw�^��b	VX'��P���wn�%��)fDy D����Fn�=����w�L����ͿF^���vN���W��ʒ�q���J��-3������|��!����kN<$��dX������W@���f�f�$:��%U�lF_]����fO�� �xX�?ֿ�Bw�▘~����$���w�^�@n��Z�Bf4p����N�ϬP�{J֧�����&�]N��'�1-^��K\Y�����`��D�T���������@��5�Tw%�f�?��rh�4�Xl^P%�S�${{� ���]^����;�_��]Xx4�n`Gm����];՞��0�+6�
�7;�ym
�n#�	
c[�Y��:�R���~%fqp����a��h�[f���S�G�*!s����pD�?���������l���f�����5V�a�?C	a��♍����d*��a���v5�a�ry�j�����C|bcJ�n�^ۼ�m�c���°בI^�>|(��mDJvL����ާ����oK�3��,�����;'e��|�B*���xprszH����z��D\�(R��eL���7sh"�t|�牏�H�%�g?��S?�������?���"\�@3�rΙ�}>�0{������uH��,�lu^�e>7���*��|ń����� a��{!-�������z��\2t���6���|�k ������Ԓ
^9�X�mi�qۣ �V��9�YlHި����@���E�)�bu�c���7��=��۔�H�}r��xpJ� ��G�-�
�	�v;8�-w[2�v�C�_Kc�p��x ]�|������}��K��kI�u@�̸�a���;�0Q�c�s�?h��Rv�� e�չOp�	������4�%�[*?1j���*���M!hB��������d�^��~�K�$�e�����T!D�Ϟ�'M����6� !�u�HӡWM�=	g	�;se�SW)��~���l"�7���y����|�����(:L�:�l�]�Y��)���ڥ���
���Wr���NP��7��]���U�I_�R�ʟ	����D~b�G`�(ė��������X�v�+2gJWI_z�+l&f��0�{�.��ܸ���¹���@�h��?Ŷ1�X.�V�{�KaV��-^}������ꭈ��'�e��;���n��Bf�A�h�H�8:�Cs,	����!����������97�Z��_��m��j���uF}x����]:�X�5�B[K�\33�:x$�����!O�?���܉Mj��*1�vy���^�
L@l�+��(Y�h�3��m�v�r�=_��r�2�q.*��3���xKmz8ݏ�ϔ�.̽�f�2����l԰�u9��g��Ш��of׫�ȃ^\�j.@v�:j@��h�W����w_�1���O��Wr����uX?\W��@�v�ڟw�9"�Ȳ�S�uR{/�Ɓ�?��*��+�j����]���H��x�1I�!�{�M��^�g�x�f�&��i�	��[�:�l�6����j�nĕ}�y�j ����Oړ(�k딤4�l��R�q���?�m=E}�aoCV�z�B6!�r1K�k���-�W8yp&�/{�V�������ё�<*>x8:	|�U!4���eGx����̴�r�Q��w3�.�|��-�)D�hNO Xa=xT�5�kP��6̏�,l��u��|�F���}Z�uG`�6c^�_Zlqh�ɝ����$ٳ
;��Н�I��٫�p㍂R��<�\3���܄2��fc��mq�rZZ�y� �?�#��k*�:�,�a&��E ��9�7�o���BTJ�W��@j$�$oe�u�&�\��AlᥟN�9ڂ���C�E�b���5֚�@�M��2�a�R:��Y7O? -07"y�H��;�n�Q�^��a%���f=d���1��`Ī��^���/������~R��%��V��G��x��|z�P)�2�ϖ���H��T�����#ĆSh^�1?겁��ǩ;�ДW�lg��FIfq���H.�Mh�F�J	�W�[Hp�~�$M	 o�0�Q�ƏMo��#g;)-M���lǱ�(O�E*W��`����SP������dƳ�����0��`�鲖;�6�&ߕuگ J��Jx)e������� �k��j�Q� UAP�?��0�N��E!8��_�$d��_�E��Kef�D��^)�gDxx��=��(�Mc�Ǵ�p��Bs��y����9����&_Z�a=l�+������6-���㋈�!�H�pU�@8B��2��+�.����7(]t0��+C6�Uc�.A�+4�/������HlD��Z	��٭����="�����?y�_���0	b�R����;ܶO ]��a	�Wc}V�;ޱ68CEp����Z��RX�Z�00d�T
p6y:$J4��8v%|�f񓭂X��dlՓMC�m��5 ��w�7X�^xh���]��{�|��� �h���4<�Q��S������DOkH2�7Ic��O��	�� LE2b��U�%f'$��BZΓr��T��ǬP5�
�@յ�����kln�q����$$��"�5��e�����x��%`m�Z�<+3��(xߜTA���C.��_5#8�����W� ���ܚ���gO��Z<`h��ѺD�ӄ�Y�ΰtt*�ERf?�zKsx�C�|��Ä��Ey�;����%i龰n�Qg����4O.���fѿ1q;Qc�yd�V^��h@*m�j�Mb��Hj����UB�[@-�rX��Y�l
!n�;�Lm�ׁ����� �C��F:�?AќE��)�e�w����4"�*��v��EבpZ���}�6�O_�Ki��cE�*1[�r��Πf<˟���^�@\���V.�C�K���r�+8f����8c� ���'H���Ӏ�{90V0��a�k�GG��<"t!����n�D�%���M��a�GEk�y�^�vgSn�C��8i��8�>0��"�&�����W�?R�c�bF�m�`����Ȣ)���^n��y������-*@q�>��&�Y"�6�iO4�HNf�OoQ!$�|����@�B�2d�\ktУ�������F~Н-je]M����\�5�X.��l32�m�����O�k�ft�`�8���䑟/��M(�U4�`���㟫[�YR�⋺������E�>�8޸E�Eu�4�0_1�P��tȎØ���4GD�̚#T:��='�����H�#J�5�Ul��6̔O$���tN��cynX;��>�a�Ͽ�f��=$�[4�zܧ<fzQ�5�J�&�Z	j1�7\�=
˗��	�x-ц�H0����j�}w��'�+�;�!�}�8x"�*�>$zH��(Ԇ�[ѳ|:�P���t�S��	����Gg�K�>ն���db���3(�6?C�5��F(��<i���G��El+m<�5�VYY�	�4��'�!��-��}����fQ�4��DtY�|�%� �Ύ
6f�d^���m��^D_W�b'F����9Թ��y�6�!|���R�U�s����{ˊV�cQ�֢mZ ���NWl`*��x�|��-z�N�1dԈe>�k����\�p[�b� >���G�5��@���#�>F���(�3��}v��k@m��]r��xO*/�gu�reϯ�x�f5[�^��:�����(��u~4]p�����uL~�2��ĳ����<#ldR��$�	�)20�$�GWǼ�vO$*��teeϤ�'�T�����-��]��!˯�9l��M�{}�C�X(��U|0�I�_���gA� �Ԍ'�ɎHm���,�t]�rsQ!�۾�tZA��Ʒ��~$vڶ�G�mG�AeH�;�P5���@�t�2C1�1�#Y����)�Mi�:2[g�9��R�����2����`2�x��Uٰ�Sz�s̙d��G��F�3�*EU?#�V��H�ݞX���?�^�r'9��O�����\*(�a�*�q����d@���y%�z�hM�-�$�
������ľw�����sܵz҈���
;W�%~"a/�4��!�;s��F4�#-e�ty��V���/h"�V��z��r�[�T�E:��9(�ܦYoB�Vx�d3�z8x�v]4��]�ZM�S�-�A��Y���&Y�?�?�aN�ӝOg&=@	����?��4k!�����οp�q�q���i'���)��2J7ِ��[���.~�
~~�^0
U�̎��U�m���u����,!F�0tQ�4��M�r3�eݘC]���+�9)�����b�k�U��c��N*���d�9����μ����!Ev*�����no�of�^��{=����F"�m��7nrFrG	 ��*�j@3M��H���z#g��"�MV���\8$w��>�e8��L�W���ib�S=�CCU8��I�s�,��_b�+�%&�|'[��̚,?Lm�9I=L��	*��xXX�[�3��Y=t�7d�͈��������Gx��g�t(y��[�o`N7��)	G���tc,�,�9l�[e[�$j;?�q�P�����.�W��`���y�O����i��E������h-.�jLU�:�_iN�i�|J_[��M 0ţ��A�������8*��<G�E{�B�m�/7�a
m	*|tXT[�Vg�7/���ޙ���[��UΕ*�] ��Ӄ��>��R�m�}��a=�����Т��C�2�c_t�KX�_m����!��(y�>�0���8���m*ȡTUĠt�S�Z\�	=.�c��ki�`�٧�@X0���'�s�&9v�ch����5��~���ߙ�Mq���(S�������\t�P��_�����ϡ(�_��`����*j�/����S�ω�P���P��t0HF�I�Հ]�:	ڇ�^j���>��Z}Mxy�q�\�&�h��U����9(��{p�>f 8�c��}�\Z���j���PӢ������Ye��pKR�d��<B����8O��=�!��Е��!� ᐌ�	_��p�����Ź^(C��V�wj��l�B���e�ag��S\�90��ٹ����;��W�
���KH���r���g=��jX���Vz� =��;���Q��
h6�� (�0Fs�\���İϜ��MK����ɚ�7�t�|>�����k8f7�3q������T���S��_eS��t�Q�\p�����������j</�G���M����<��Q
J�b�/�u�Н%�������3n1Ή�LsJOhF:���s�'�-\_�nCz��6��<��z�25V=4r�? 9p�FV�d	�G��yo�t��s�\�wUD����X����9��L(j��{��,ޒ̺W~Xt�{벚��e���J�0۔[e�] 8�\&�N�]�ߛ��:9�������Op?�t�1`/UrMt�#�T/�;��^�T3O�@��z�2�N�����ǂ~ ���+rO��U$�<6V�T�+��⌘
���LL�2���ߪWYI{����IE�iC��9����-M��a����S\�Y��8td:��R�)���Hk`�2�~tN��q1Փ[�2p��b�8�Lg��_����E&�9�ϵsS�;���.$%���RC��[��84��4_B$4��d�(V"u.���q�˾\�Q,o$,�v���w$��l��f'��TWr먒�<x�o�[�bQ��StK}.����H>!J����	�U���ܘ��93�����E�c���-b"[��.�	>�m�r[��;1e`�� �(Y���Pe�#ᘎ[�KV�-mv^�r-1j&#_�X��!Gy��,�-iQ���P��aN�!`�,������IlJ���P�C�ȳb ��dg�����w"Yy�i6u.���U��6}���\����K�z
�?o�;�pl�M��eΒ���:�J�й���;S��s���utd��R�� %M�QC����=�a�u�7;���A]�1d�M�K���k�$�{e��	�ji��;גt/y£�ob��K���1���Ǖ߳�1�����U0�K��ǧ+,PZNó�2��+�zL3��}��͉��懎\N���p�LƽSة$��UጃԞrK:Ҿ�?��H@v˚)�̴#�ׁc����]�Z�)�%4��*E��H�^{�����H�T���X���y��ԙ�k��s�=Z�qE���P\�4M�M��0.��Ӻ1%����,���Ps䯚˱י�dK�*�<-@o/���|�� T�|u��U#'���Ĝ/V��E��*���"���"(�% Ga/���a��m+�*T>v�ݑV���2t=��o�	�`�u����ϻ�1���fS�$���x(��-XF����ɴ4����̧;i�gw��� �3��#p��_)9;���"�Y��|H�sh�����2���B=Y�����#�ߊ��hq����Cc1f���8�G���=�rRfL�+^#܂ �hO;n]��o��&�S=���v^I!����6=d��o0��Q9@pA�Zu�Y2*��Y3���yv�Ē�SW�O 4ᣰ8�N�]���f�D=<.�Yx�̃o+y�E�a�y�S1k�(:m����{<K�>��7ؽ0O��B%[��-��i��;C'�J�j����bM�ZS$�`�^�Ә����>���x�^G�|�!*9ˬ�f>��j�Q�¸�_	�o�|�<��C��[<k��5p��%	n�9!2�s�*�_I-�5����i��w�����!��I�bw�L�V@I�?��\��m����r���椵�;Y6�Kxe^Z@��	F7���#��1���G�K=B��1��.x	+��OTu8݆�.]������g����h�P��r�s���(I���3��M��O*�{�w�L�N���~ƥ'����~��,�0���\x��1�L�2�ɺ���l �)��3����ې�j�Α��A�E����B3�3��6Dɢ(�����!��(�%yalB�1V@���Zu�������#�ɷ�c���R�j�[s�	6����G����5�G,�=V�����]po��C�sS�5��07��^!���K���8=�7��|� F�`j���:�tNn�,�2���&1(�L-��Q� |G�_a(8�\Vj�b��7VY�^��il�2��.�u��"����R{���M��fE�BŤn*� QK�ǌ>m%I�0�������\|��-)����a-�rS��ѯ(7��Zm���S�ț�(�1DK#O(��1E1��/4����g�J���B��I���"�_�)� �
��y��@��}ƞө���Ai�}6��+���=ɼ�+�3���H���/}{\��Z�-m�8�K���m	��T(�k2�b45�L�*s�%y�D,��*��Ĵ�A�d-w0Fz��5�D'L2��%crк
F��~z�*��a73p����T��2��XR0��E T9�i�lU��d�@�W�:��`'��B�&�����)�V�X��W�uc�C��B 4_7��=�A�8��ޣ�.�E6�j}�ǣ��yf�C ,�E������+�At�l<���7�R��KS-��-wKNF4i�9�RI����ɡ��Y���Z�i���i�b�_�fPj�M� 'G�8"�W�s�;g�%x5!ƵV~�n:�e�N!��>cc�7kG�o�xf���e�
�i;��͡;������q�5*Eq�l����Ά�������m�J��K�p�ԭ�g>��ҾզZ|
� ���"��	�F��}5�^�����P̨��+BF8�BSkY����z��$a�E��pS�"7�;�:�]�-��n�7�I�R
��l�R��ҹ6ˋ���s�U����A�^�X[Xݹ&E�g'Գ���y!S{9�'���#e;k�ԁ�E���^��yT�����S�(���dh2@�DܒIn���!��v�rw���>�1��%�-f�Rbr�b���6����Vֵ²:�.�K;���>��sZe�-�V��xb&4t��ZD��_�;�4]3&�<�����1@�X<��MlyՇ�^0�޴�BU�s��XG���ߠd���J�+_Om��ڣA�%0Pn�S��Z��+BFI��s��1ĲEam��lAR>�[
\̀lĝ.-�k�U�S��-�[&{K*@�#�]D�M��k���{�QX%��T������@�rؽ!"V�2�����L�j�\����	M�#-M/|&�/�E�t�o$�e�bW��Ԑ�/��-�����w�l��з�-y�&U���s�a�\n�W����O9��ձ��E>В��ah4ec��[0e:�щ�z�e���XE(zW�i�ݗ×pRC��[�Ț@�͎z\#U��6D��ܜ�2�v1�:؅�T��L�����m��:$��%,��~r��b.�	a�z�7�ݞ�W"T����S�� :&�Ω���A3����r���^P�S��Z��)�)sd������4�r���t�I�L�9�5��1�;K��~���H`��������{g>cD;���c8��V_U�3.��t�*�E�k2t/,�c��d'Y'���)�H�e�l��}��>�+<�'����E��ɑf�#�(��Y��.i`��$������Z��6#�/�^�"�/�
�P24=��IM�q~�99%<Y#E��WmzEǶ�#�<�]J��*9N#FQ�Bm�#�ӜqMu� 9�s�#�[�Ldz'�ed�e,�9�Z外$�?�Ǆ��=D��ͣ�{�l�=�2f��<�8U)����3�^�W�@=\q/��4(���ή?�u�ǃ26�����G_|kF�$��6�dd%���^���3N��e$�0�b	R�Nئyi2� s["<�|lT�XO��)C�H�����NX��������\	���C���H��8���-�[��Y'2z��W�����?5L������#�y