��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�3,ESA ���7@B�h��ϖO��lHa��&�˸�ɮ��Z�]�V����7"Gt3�>S�P,3Z)�~��1Y��\TF��;�$��l�:�����&�{/�ڨ:?X���:�/�>A����Q��3�ꉐe�%�����O������w�9�c���i`��S�����n(b@G�Udh��+�����l��S���_�Н�M��[n���%t����aPNl��&H8��<PNw4�H.���U
�ԜؓD��	���d��<	zi���3ϯ:o!f��f%
���K+�l�^>�s�ȣQX�'���v���x��4�������M������'�!�LH�xh��7�Fۦ�ѩj���Pz�����4�|_�彞Dqm��{��'� �r9�w<�?c�
&1�_�~�t��Vf�[1�v����;4��|���
2�ŭ*T���]	,�N��h�ڽ��	Ȩ{A��F��P�]~ԭ"�C�a���gN����	b�������4E�h��[�t��K9n����u�nH4���w�6�b*-=�ϼ%R��A}�����l�{'��,�:6EZJW��[��=�!?x��]�LT�i��������у0��K �Yu�bJ� ���l�dP��9���Fᡭ�9N�O�3�.�����5s4~[\h@�)hS�V*�%��;:�[�X�]��=K c���r��>,P��7��OI���2���l0a'� ��ng ��&AE?��+�f&
���s�j��Z���)�3��,̫� �F�/�	���Zܐ�o%�h�A�t�Ǥ	���[-�����AR��5��޶��	�Iz�ra��4��w)�i�9:g���PY����~G�]P�x]�q��).м�ԽbC48���(~Z�@e�N���|q1�� ��_���������J'� &��#��(�|(�*��[��Sv,�V�N]s��\��C��&��c"�*)fj�c�2d
P��-	Ӊ��j�彋�"������!��O����1Αg�^
|'�q�p�Ձ�kZ䄶;Ӿ?��W+vX2�l0���h��}K�Q���-�,�)�|�@�0(l��]�����l�J������/�A��w��%�Qbr4_)�Y��^�q�ۄ�4��)౾�e��~�	�x޻��VDЯ�$F��J��WX�m����NZ}��( ؞�X�����lW����3��;{�_��6�ho4��痤�*caT�I?M��j!`<G$e�C����{����W�S�3#7�?	DI�i��Vu[��d8h5�q�?�͡6J�4�'��>�6��kroʩ��K&!P	g��d��(��U�S�qi�#l�xӠW��4�!��N����-����g��ԞZ��~�@�}�>��kqw��]��Z9?��w��'�I�:�glq{FQ�� 6�G�hr�>��DaLG�Ѫ8���G��V�'巛7���&��k�����Q��N����J�"�k�;<�����
�Acpq�L~�F�͎ p淏PƐѥ����B	:��DRJ]����1Y����P��DO)���ڱ�0�_�"��G	���a�u_��� �1�����Y���3nV%`/��cY�I��@�)t���i��_hWg�L�7�q�����m��c Ϫф�}��^�E�W��Oz���e��) �	����4�P�.��A�����~�K�~��/c)��� �W>�cӺ	E4�#;2�2�Ǆ�̏OK�9��}s��g�y�D��̑��c�[� ߇��n3?.�~�T����t��}��X�&qs���K�s'���ȥ탈uqN3���Z�Ӷ��j�r�L�ЧC���
8�p�YF�ˁ�����	d'�=	z�[W)+�>���BJk��5����ݷJ��S�B����4Pv�I����kԥ���<��FgǕ��`/���.a�6[	I��VW����ڢr�GT���r������̶���&@��av��f�&�#f#�u�]	ƛ��z}\),��[�W������~��Z-1��]]]Ar���K�P�L���"X���0��t��Z�����I!P��5B%�2g<��;�d�<�$Qb7e.��j)d�=��ޫؽ��A�AT�&�Z��˵ 3w��5�&�$ϝ��բx�YY�aȚ�w%�q�� �M���n�9���`j�H����;∡��R�U匧�j��G��)g,:Z�k�,�%z�?�<�PO���\�s�Pf(��@����1)��|Q��r�r��Wq�B1�Og��
�j�F�@ʎ�d�����Z�M�e�O0R��2K(�4�!	*��Q\��0���Pj:��
ֳ�7dq�,J��m9Mjk���I�<�6`�� FD�||�<�Z�W~�l�u��i����_�Ej3�ҚY��Tt�b@��EM��e)kl�Bx�ʫ�㔐P������+\���ο�V�1t�\|��۩�ہ��D���r.m�Q/V�A��r��cLѝ� vk���W��cO s������X.����$��ŕ�N��j��._��B�M(��y�!�0��Z�K��32�+�l�i�ul^c���oJ���qI�q]�?�n�ʡfJ]����Ѻ|n�D�?m ~I\T>���e���,{�Hs��`G3	'�!�`�|�^3�$"3�6 cc�t�/<�I ����ťÊx��y�k  ��O�'���V>����nퟬ���q��;��zI�phlL��n'_��ԮW�A yC�L�kY� 1�����q�����@�Ƽ���_:�3ǧ4�|W�����:k$1R=bxJl��yc���{���\nB ��!�%=
�Ϟ�a����E���d�c��� �CI1:BJ;�NΥ����2�@R<���jpb��$e�����e��^�>N}�L�a��vJ�����f� �.޼Y#�˗8� ��H6���{��*mTi�Y3�sv�!U�g�,/Ο.�|��)�%��1�Y��B �V�X��X7�D4������iý4h��o!�U��xz��#�*bg�8hc�'B�̕�D���Z �J��ly����%��pҘO}�N��j��/����Qw2�c�����&> QV�]�g���V�ׅ��	������ I� �4�E_�s��s�(%#�% ��1̜�î#|U�U�_�����n)�ռ�N�x��y�%�]�)��䬉�qmH�L�$9�� ~F�S�Y����b��a��o�e{d̼��tOjۿ��w� j�َvawǩ0��(�u[�ZCܣ�T��������4C1.�{>�|ƥW�x���ؼ(��֗Q?�9yГ"ĉY�Y^w��g&��R�e�Wٯ���1XA��x�<�SN���W�k�whq��ӣ�}�X_6�l�k�tJX��.��N�~�ˢ��:���\� ��4�޻WȖ����Wdo��T&�n����7���p����HGC�Ǩ��\z�R��U�$7nWi&��Tfu��j�Eƥ,�pP�@3�G��:�t�s�������<4a��l?Z��0^���B f�2�]|�7�S�b#kڜ�A3 �fЎ ��@�q��f��ou���nUHU�44�wI%�8:N���լ��%�8����@q>N�jG�.��l�
���2������a�r��J�p�V�Ą�xUۯ�٢uqD�bGo�),����"`V� b��+��~$��	߮���]��\ w̤��^P�D&2͸6�7.C֊����G>G�1%ʻ9;9r�����<��	���G��",��d���/
��U����a��ɺ�}�۴h�8#.��F��Du��L%T�)q�{�x/����2�w�ɗ�O��.6�=;
>�M#�N�hv��[��V�c��x��
 ��_�R:�;jOP\�d7Um����A~�-�%m�E�Pke�Ե���v�'����\z=s�J����R�o\M��T��7��ʣ�t��� CÐy�-��;��8�S �˕H;v��9�5bb�(R�gȒ3�%�E�����!��~辔nj"��1���� ����ue�7��ٿ��2Oc�;fx��X�k�/��ׇ��Oax����w��*���W��\�#��9pI.�B�%�S�Z��G�t���ʁ�y�?��r��}�ϛ찭����$�G1s��:@��
�����z�w�d1��k-�QkfK��:�b{1��}�B��TO0)A�j5ł^��^����v\Ls���m*wv`^�Ȍ{�X|]�C��$UBP��rb˗V�g\P� r1+Z�u�K�)(�����pſO�L ;ߊV�B�B�n�?%#V��E^��>(��|k�1�x
�_.҅��o惆��(m���8��ܴm�R��{uW$i��Sp�҉Sڗ]Z�Ȥz:��:���ou�0N�R�[ru,F��dw �M�o��1�M���~E|\�P���6��f�9n@�M�eR��7VT���V~����$�¶��GX�o��������]�h��s�ؐ�9�Ur�|����*����H�E)zw��Y*&�y����q���K��C� fOQ����n�hW�P~���߭>���&l�"tr1'_!�^��M���v���(#�dK�FOG$��rxzq}�q�;�wʒ�+��b�*�TK*�V����JTJ�?�[����.��A����W (')l'a0�}|N�ѣ��@�ˁ�5J��Tޫ��P�6t���$�!J_�J"9�(On���qs�:˱��W���5�w�ϰ/ Ӓ��Ҩ��즴�#f��.��u�oO%:%	��)K.�=2qh���i?���,E]=D.�T��$�VǄ_�_�n�Ȝ� .`�T�̠c��դ�æ��Ņ=S���	�R"ZM���[�$�j��i��(՗��v���%5��,��b�vŷǵ�#�˕~?AoF������kEPCLoe�Ml*��ﴱbO-!$�zx�'�Zf&Mz#R/�ұvl.�6��n藘ikU.���]����������a��J,#���O,�	;�v�2v5��nIl;�+��(Rvv��j�Fx��ͿZ'm ��3Si�L��⬺�O�Mܮ&��K.��j�>���P�G�b���g���ʙ_��i������"m��(�t��#��#ӗa1DK�/�+Q,���ћ�̚[K���$������1~�\�� �AYN3��"oo�/L��@ٳ[���Uq�NR�rk���{7	h���<�Q����
��U:%�Φǘ�^�)�x��� ����|2�j;?+��)a�uS}���mE� ����K�׽6&�4��MÞ!�.$���h������O���̥:!�T��f��7���4��� 
P=�j5h�䦕�³զK~g<��&%�^��1���,1%�LԴj7���LJO��έ�J��_����!��%n�
�'6��6�(�xU����.�����[/� M�PyR�v��U<���x�c\��?U�/\��dۅ	_+u�܇Q`�Y�'��>�wFbK����]U�c����0d�V
"�
j,��/�X��'2�&C�MO���T�̝5�݋J��KfJʹ��@ī�|�N7�+�y��9IJu^{Bˈ+c�y�o��2�kD/~
��'���9B���4��d�������Zt�E�,e�&v�ث�m̾���6�vO|����D��W��qs��a5ƚIi��m�ѩ�)"Lh�5���4�py|�=��F[5���Z$��@_ր5�����?�r�m�?�B��P�2a��&�W��K��B��I�)��r�F�����Z����+Kl�,QvL�z=��8ɨv'�|R:c��rWI��|�jN���Y8	NR�������%�W��F��5V��F�Y����#�j���
$rğ��9���`�{�;���l'h��W!���i���ƍ����E�H�0���lr 4Fc����������z�j��͠��74�Ƴ(7���FZju^����%�o� �M5y`���j���07bp�����A�5?��dv�O�˿3�^0���$��`� "Rd�'o�C 6)2Q��wNə1K�-��#W������=�-��TbL���>a�m"{�7_X�!��%��ֈf440����o�l�*�(� |����h��c}�owJGo��6X�q0�� �c2Ӥ3�~�	�8Xi�%��/�B�yqM&�"ڑ�F���H�.��n���0���@�!�W6�){�*��~��� ��	�1ѕeb�3V5cs�k�a�/�[5}o+H�!�C0�U~xi�*�H��*��Թ��\s]=�JV�.Āy��/N�@<���P��� �TDOWM��[�+z�/�����cJ�w�15�i��<�w'h�0ᕦԆHr�r�3��"�z���3k-�W��U�TN�k���܌����j*I�(��p=��S��9`�:�:�>>��w,�V�J.���tK��@*:\_A%�[��Ŧ��G�?�8&�>:�N{��I��r����R|�ޱ P���>C�U7pYK����)�T��H3ٻd��v��R8� W(���@,�A$����t�Ip�,�7A��`�NP��$�fD����'[{�H��.ɐ��9A�P�g�ٷݣ`��=�}x�����T��s��x�Cސx΄�gRc��U�?VF���uEaCxNs�g��i�������J,�C�6+є:��B#��E�����ǡ��bW�!�4r��!�L F�yެf���E-�R�j� �������b�?���K��1���=)�Ps�yV���6��E�8������b�f#��]���{y�����Q�r!z�.'�Ut"�D�/�����wU���",�����f�2m���|P�U<�+ �R���	�텐r�U��$a�R��h�:Po�xP�PN��4Ø'g�K���ԗ6��j=�,�T�݈��1�χ$׌�sZj�@�ΩL���+�sI��(p������fAV��S��t��oۡ{-�
iη���'���M�OE�ͧ90R{q��*��EPpl�1��fY��L����+�B��I��l
3�ՉO����3�Q+�PV'��N
�+k��Ǵ���I7�]�=}-~t�nBX'2&>��fS#�s��Q.|@.�<��fYfuǴ���G���-n�>ݛU�q�wm4�uy�bPT�XV�:�9�	lM;[��ܹ��:x������������) C5 yi�n��b3|�׿��I-%�?�d4\���-kF+��Hb�*��G��ok��
Y���o+����C���֫��n�=ɮdo�R/�N����q��0%TЄG�S*���c����Rr*�N<�i�y���0Lڎ�,��j�	8�Gt�V��zd4��D�ҋ"?,�`6䓝,�N)o$?�!-�5�¸uFn{TE��h���oBB�݃,șη����۱,aHeqxf�/�`D�L��D�}bO0$�M�a*\�V�S��^��K�_���a҈`YR�`C,v�9S:�q,��%�>䉎r+QJ߿��.���R��Q��L3����c��	e��E�+�9��M�?j8���+�B�dk��
�n!��t<Kn*��t]�g�t�	_�u���3�|���3��i�F�O�4��wM�x~/��̸�s�7�RP���EX���8`�n���#���y'����i�O�˥#�^�-�
{�};�oo���r��F����_s����1��������\��3��D�D��/a�ڝ_�V��Ni3��Ƨ_�5�E5���SoDyxˎ��N�(7x�{a�&��7`k��r���!k�����t��^�����H)z �h�>׉Un��=f�1~���s0A�Jv��r��0'9�Djh�-��MUlw.웈N:N-Cț�
_,��|�iI����y�嘽�Q	7
��s�Ip2�⚐(!en2U+ Xg�)m	�����-���O��ϳ���8������Ʈd;��\��&�KS�)X�T=j	Z�r�0�R̬���՛eQ8���N�X���"�OН�N�֮��W��z9�a���sW���Te��B}A��	>^����N��GT��z�����ň�ʓ (�T�|��EMe�T��,=��T���gu�}hMT�l�ŧ�<u��P���o�n'����I��Ş��γ���~��_� D�&޶n��zhT�2����1�o3�����4��&�,	����B<�:z�G[�H�bX�f���~`)d�Q2�T�[���Tm��FҰR�W.�r���raF��*ݥ0sZ�с�ٕ��٘�;�*r}3̨㽷�sY)U��Y(��4W!3�<Dzj�#G-�nT�HwO=�(~W�
)Ԝ��o�L��G�x�X���B�<�$�?�5��kW2��cc9�l�C�?b����Ċ�6���[4"���p_H��?�����w��6Z��e$��"���&c?���6�a���mM��U��&�c�6E���Y{�:n��cW������!Q(�H�P�!`j�(�i$�4���q8��,H݂���M�UʬO_���b��:��-)���T�	�U����q�1*�{�pîix�W/R�"�P=�곤�[�
9��B��*���V���[p���(��F�<?�DOc�~ҹ4o��Av��ݢK�[�C!�'�c�@&�k��U;Oc�}�D=,c��HL��2
#|VO�-N��o��7t(s�N�R�>���O�U��+���e�6)^��|{��T���w"��� )�o��	��ا�ǘ�¡�&F���M_���2RSX��Z�H��A�fQQTǻ�1KH�vZ,lxc����ǃ�?�Jq(1�S��[W(��[��n	�6	����mdU���Z�']��k��|�+1z�ù��1�inm�/i��9]_nZz���z��d����Y7B/��C2e�O&
R��a~��bR���f�V��h�?�&_h��q;L�0/�9�r;��Q�vA����K�~(�1�rI�� ����	V~^_���[*��Ϫ�=�缝�A7m��4��(�OX�BV�,�cn^��a�?M-Lm�N��im�s�I���=x�Lu�x�q<��M�\;١�5Ú�+JJ�ӺtW �C	Ġ����z��'dw�V���
�t>ra j�u�7�É '�)͝�q�Ǚ�n�m�J�7��h��vb�T尦wpA|��|g2��-'�kHW��G�-�����HO��t'�Ư��::xϳVA���!����hef6f�n]�t9�i�6�.۩���^0�6U&ܛ�� ��iDD�Ñ!�u"n��;'�v��H?�a�s��ũ�,!��l)u F_�+_����/��Id9�j݊�M$I&��Scr�?���YZ��Ll_�Ν�@s<�p�{աt��*5��S���q|��"eB[t��ͬi"��E&DsP������@rP�[�����3dݨr�֚�1����䟀N_��2e���UM!U��$�f�$0���0��5]U�w}o��G�V��E��gǶ�&�����FO:I.��W9lc��� ��+L��U��0���2��8�]q���?�$	��x)g�;���ė�;.y�x�<�����_���^q�Ե�x�R׋��|�q܋�4�v����|����"�t��zJ6S^ÄΜ�gW�K��7�"G�0��x����5�[�2�n@q�$��/�4��Aִ��w^B�$J3g�̐�݃yI�׶�)�>xW��ѫCO��Bgԋ5Y��Ti�ʶ>l��L9Mmߖ�|�ɧ�	x��9��_��:
䴼3�,�o0��a���i�)F	�QPί��m��KT�7�/��_x�vMB&����)P�^U1<��#���E�v2�讥擤�FK��S��C����~Ԓ@��4�>�����Wx�8q 3Q����� �������85Y�\×l�p�B�M*T a¢�+ $\�g?�,Ա��23吿7cb�cާ��ft����F�3����ZܿV�uCٯ6؆��\j$j�ۮZb5��Kg��ɢ8U(���:����٫M�\�'���f�_h֟I�M��C[������1�R�C*	^���Y�_���]on�t�}��h���{;FA�.��\�|j*-#�٠K��֩�EaS��u��f!V���h;�*�����
�VgDx.�lc?��u+�EG#Ľƌ�w;8��1k���=,Q���S5?\~{0[����FOv��JR#Nw{��/�ݖHM RR�{ќ�i3�geN�d�1� ����1�\Ӧ8��X�&�7�9�e&w@�����&�	�/N����������
����7�|�i�|eO\�C�WRr�p�?g ߝy'�}�'�0	�/��h���r�c�� �[�����L\��1([�#��4\$�|�tw���Ƕ�o��r5��J����2`������/l���`��r��c��O,���O��Ҫ��H7g�K7��=\MZ���[��M���UL�x��UO(K��M�-��<�_Ve�����i�}���}K�i`&��FcS�԰��o�c��-c�n���XAS]8�h�4PWs�圚u�|��M�]Of�񩱂G��^3�������Z� �#u��\�k�h$>�p�p�3�y��]����q����ȳ�cɔa���[@'����\9���k��]v��Sw4�� ���U�U��d�1s�׎�%�M�D1��ʝM�f*X��
9�$�%P!3�D�C��%؅A�_�[3ی�	�L����s�
�ﶜ�/CG�ew]6��{�d_q���F�(s�+:�3R���J�r�I��|����S���^H~Z=0��{��P�����,�4���ű"�Kj*x b�ɹ�"��D� 6R� z�2�aV0r�*�%��^�|?�+5Z���ۺ(�8S�#���\s�[A��C�sw��|��z��2�t|��<U����A��fNl�x���j�ͥ'�hK�
c���g�C��9ʱz�y�>z��%�z�*��R�,���[���k�[��\�����}@�+�&��.Cb����}Sy�%Ν
��^��r��DFMù5��\	��"J�PTu4]|Mc��f���I?�4��O����l��W-�,7��������R��[UŖY�)�Mu|}!���12Dm����M��J/PU�]ޚ�1��߿J$���i�.Dڟ�s�_Q�Nb�"+)�!H3�D�����6i��2�+�ނ�H Z��91�=B `_UWm��2:���<�因�E�v�����&��>�%����SM?ܬ$�\+�葆S�#Hs��K:,�2+9y�A�k���)\�{��s�ЕJ,��E���	��Q@�]�0�;hvl��5��DZ��Di��>���)?���U�-3�ދ�����O �akq5������̚n�ٙ�vԧ���E���urXC�Bc�Vp�GW/�QL��7
_�V�;lk��L�`��ʑ[;�?�?�F�����/�)�,�����K���*��-z�	<D>���n�^��Nw�B ��Q�.)G�����ʏJ(����V�pC�i�0��8�JmJ������Կ���h~�����a���)�]�D�B���
2�>�=6i ��b@d:`��
�?���lǼMn"��{�D�)����$7���yZHl��0�N������آ��oa��A<0AM��z�_O�"�FT��jPV6nGX�sx�?B�K�|*X�w?���'�z�g�"�8Z^H�Y9���� �[#Jpɮ�@�Q�LRڝ����HпZ�����ħ A���<38}W�J?�� R�?����%�t�ߠ����h����� @Eg]JL�:?*&Y����2K��7n�x�͘��#*��u}�R�A�L�������2%�CN��A�[ W�K�P����ȅI|�aj�Q��ϕ�עG2P=Ll��/���J��m�2 4z1�D��x�>2J8�0��yL�rs�xȄ�뀑���)��5���zv������
9'��r5���1�1	��r�*���&�E���K��_SO�6�pL%���I�4�79�H�+&&�dv��$��{�͔͆����>�O����'2K��N7 u�T�~NȇA�7*o�P�Z�Ϸ�E�=�'o<O�K�v���pjjw����OĘK��@͵��r������0<8�TD�G��,���>�T~����������Rl�9 A]I*�Q5)=�S�E8&��ѲO#	ZM\iv���U'Z�n�x.�����r���>/<�$�]��6vpR9<���e��#�^�S�ф��KJ<"�zC�:����s��{�ؙ��NG�Co$P�F��a^���ߓ�(e��4�+]�`j8H�	t;ŭ�Jl�̃+n��+��`�w��IFxc��W�0N�R�^��3U��U�w�"�]�p)ڮ�D���iB}���A����&����9[|�b	�w��HF����~���u9ͫG��s��E��|+�-�X�E%b͎4Bz����Ѕ�FAȉs��-�n�v��%����Պ�EA�/��ʇ���g5�R/����GK���
��]��<�֋>���O�j��E��=�,g6:��~�R� ��u<�N6:����ǂxuё�`��S��F�epbH��$�]f*܅�j_ Sl�|)�&��#��؎��4�#�k��Ո#�J��K蠵R�[���gQ��#��nC����]`	�ҝ��k �F}���V;��}�ܢ��n;�<�c�'��h�W�┱���� c]��d�9;�:~m�H�������N�<$�������/��%\ ��&��$���'�xn}�����a�Z	���<활���_�(~�oo�+o���i���y��cB��Cq��c��OY-�I�T�{'5D	һ��JiJ��i(U��7��v�C�Hm ����~f���6���-��t`��u�>�Ѐ�TW"xT)��_3����*|����}���_LD`?{��~y�f�g2�c��F@�ǒ${#s�q�`�����7S;�o<��"�>LLȁ??��[�É�*�b�^��V���˘QP�7���B�FJg��_k۶Z��{.`�h�8��u�k��񖁐;&|}�ke�bYv��nKV�h��L�崢��aB�qtL�Z�z9�P�ZH��;����Ic~���2�z�X�K�s�i2s[�۔Q񐚗���h�nt?��\Q�h�^��<
m�^z��
;�xj��dp]�O��$j��ˎ)j��f�զ�a���h��L�%?�"��#V�73Z�'��3
�'�yl���z�1t�4����ھ�e��/�KFo��Kb��K)ڧ��� �>d�7��0��ui���������ȥ�eMP�a��"�r�v|�6�#A��J���+�hL����(�{�/].��I�A�L�QW��Ζ��a�ݸ�h�fBF:�,��WP���h�H�d��C4���Ȣ�>����U�%�J�t�=2�&Y:����ˣ��?*q�_�i�o��W�iL����i�h��3/��o$��E�s�ښ�UJAQY[����g3�f�Er&Y�K�C�VP�Z�ǹ�t����ѯh!"$�_���P��#�4lb��E ��!�h����ϛ{�w{��<3�آ4�{�����<bl
��.4��`�2�N���Ҟh:-�r��3F�8�aSvF��Pߍ������������IS��s������۶�6�o�H�$�xQ�V`�fR����� \����Lҽ:�H����c�٪��X�s	���_�*S��qn~��0!o��-��*���+���p��Ya��}H����^"�4pv��WЮ��k��5.�絪r����@�K�/T*A-���M�6��/vX������r����E����-��{P��լ�`~\r���[��H���
�A76%V��
e��H�����Sԟ�#�N_����<[0�xŝ��"(x�7�y�q梐���Wb���as����ʞ�*�'��z�~�P���ݍw�J�.�B�q�I\Q��/�^ɷ����\	9�ul���&�t;�Ҩy�'b]2?(c�K���yt����+�J�ɟK��$Pa�#�K^��2k�lK@)_|-m
̮�����E�`�*���r(�Zy��?|"�����ek"��A��TvO��ie�Vӿ���Sˉj*�!`�j&z
�ǥ/�c)�����P�O�f7 ���y�0��D���6A@̋�ul-!"�߫G�����{�P�#�K��.M�"7RԴ�}����H9�:��,Y�'���`Ѵ7)k��Fq�I T��	l�\�9����,K����������`�x���7E��\w�E�(�~f�(=O#��J��x,r MsH�b�eѾ�t�CǊj�y���!M��E��C-N����n邂�s�T�WE��:�DiJ6lfE5�:Nt��:��)z�s���ݤ�����]��E��kP�`IVZM��&u?��-+���:cWQ�O�����W0p��6��W�U~�P\>�ƿ�)bX�kb`9ƥ�g��y%V=�*8b]�"2ш�[�B��;pe�Q��u��7 �:�y�2��У�Ik�C�՜����(~Ia��1�#Ȳ���:Fh��{b�Ȳs
�`}yr ��jUa�UK��ӑ��^t�6��K���h[�[��4��@L|I����Q��MOw}����N�Hd�6|U�'C�+|�L?����s.1�ڟ��� @C=a뎾e�C:�'@A�����}�C_G�J5��}�9�Ԝ��-I��4��ȕǖBs�&����"X:\,:~z��c�GK�n�&Hl�(!Y������xIQ���'���냻X�ô]W�P1hS�\x�!��yr:b�ӎz9I��f���� �a���x��FaOC?����UC9��������@D2,:��ϡ������-+d�,�)�����L��ܹw{�������в�3��c��JP^�)�E��ׁ !&7���*�/��h(��a��)����dD�>�|+����Q�hN�B�Ϝ��+3M��;�Iw��E���M����;�d�f��`���"^��m�?�)|GȲv�Q�TҞQK��� y�v�K渹2b���r�h;���{܁�Q��3�B�D}�',��<d(����C�8�˓�z�;�F8�Lf&����9�!
��v�-���lwK�x0lI#ܮ�'|����r�k7f
���S�S�I��9f؂:���J�/�=���z���<��?L��Z����Z�x�$8Ɉb]�N�,�n��؊<z�a�B�I��ޭ�*0��H���إ&U��Bb���Խ�T�$�5����2'P��[�d$���[W�(ew�pO; ����?��]�����3i�+��?X9���D?,آ9��Q�����&�>�N���\���h'g�����\�~�B^�}�s���rS�H<ŷ����5"�x�ղGZ��歇��7Q���ӯ� ��O�u�#2����em��[��\g�>0!��h9�C
R�+�Q�%ID=���!���(hQ��� ��mL�L`YDn�5S�q�d%�����=��=�)������Xz�}.5�Q�����-]�"��ᙧr�~I���P���Q>7;uL��E���9E9#�E\`5%E�7�?�)���H�4�� �X�p�����-<�Lpfp<ǿ��[�]l��m�H'�ʴ(? ��v�����"ʿ�~��s�ك�>:�4d�0l�>p�f�:)�/���V22�v"sl_�[�(J�w�.��`���f�N���qa��~�NW���z0�^����-h1�w-wS�["� ���%�˶^�{I%K�1�W{=>�#���lIoԐ��>^�(�.s�bA��^u��V�
��&z�$*:�>=�i�FM�N���)I�Ϸ-��J	"���N‑�PD��VV�c�}����uI�h�ZCԓHW�R���b�v�&]/!����V�o5P>`T��$Ğ��o�Ƨ���3�z�~P)q�����шy�h��T�A���4Q���I�|��5)1�q������
����A��b��!� ?�7�?���t��Y�N�jFe
�\��Jb�9
o~��y�8bL��":z�C=U���A����V�oR�rϘM�_��x��"�!����['{].�pN���f9Xڟ`Ǣ�����sl/^���D�nl)��O��0�M�3�/�R>�8zT"�� C����n�	X���u���T*`T���ܙ��v&}ɃC���NG���ž���j�)]h�{	e�@9'w3Qkf��F�	���ؽ�HY�v��k�E@���֡�1���跕�Ҵ.�����wR�,�j�$�h�� &�<NS�V�e���z�io{�7�?�����?�nL�*��T^���c�8�rf62����c U��\�Hԉ�1Ϋq��v?�隘b�{a֖��;������彴�8�{�>4H�2��e���e�����O���>tٷ8��.�.����[=W�̾t��1���A�L#ł�T
����Ӆ�$�{��7OU�-���Pf��S�-)
7���n_J6���d#��!8<����6�)L�@n>�5����疑ۿ=g b�0�?��Q8FSǆJ%����3��n����+�\j �L]R_\\���J�}ϓŅ�M�����9�7�(4?3
�!�g�|���)�+4ncI��:I_� 4���Uq����ҞH��u"�а���&��5_�ϑ��F��H,G� 0e����.�Qj�R���G^,�}��`��r7v���@�Y:�.�
���~8��p�(M�� a�#Q?2B��`X�l�������!�
K��v�8��{�XB�/P�h��8� ���I�?LO�8w;0��J���Q�F�w��m�
�"��ͭ�g�7��2W]0����8��l_�D2v��-Դ��W��Ճ�lH�]d8	��X��M��@��6eyE�q�Pk7q���٢������G�#��JK�2�~:�r~�H�� R�,��,�BϾ��s�ω�|T'�a���'W���s���;�)�ן��$G������.�+���I��;�s5�L���4��td|(x^�#}�����em��x�u��y#@k�0�G�Q��m���_�!�i��]
r,�sR�K��֑��W#C��,_,�;�S��iN�����+�v��լ�pZD�� �~����N!�E�̻�Xo�M_�n���a<p#F�+��z���2�V�"!6��+8l���es��z�����4T~TçxZ�r>S�3�]��gMl�P{&�7�gx�HP�g�fVsGf� ��4[��j~0��+h�0]ǰ󫋚0�X;���y����{a�X�J�h=h-��.o�o�)�����`���~�����o�o�9Q�(�(sd����D)G�1jX�ʦW�T6Y��	�~��������}$�E�H#B,>ZrD�6=���_ݲ�W�3	a��>lc'FaE��I���H���|�T$�<ڌ>�5�HbD�����3j~e��Ƃ'��ss��Z��qj^S��nl��Z�={h��)�)�*&�dw�Z�EN3\���>;����K*LV\��Q�]F�:~F�m�$G]CU�ɷS���qb~^\�r.�ͦ֬=a��N�M��=�#��Sq�B�_�!�>��%��7�mn�tý1�	$�7{>q��G�)����Wr�;�k��9��t�=�Q[e?�p��O�� Q����
X&;f(�@���?@�/�83����h&�oI4?`�G����eE���V��n�m>�'c��-E�]ܗ�3���d�8��	RpS�Ua?F��H��<���D۾N�-��O�27���[�� 3�.i`��4��S9��ܶ[���Hs.ʈ�Q#o�~�����IU�*��94G���η�!�������C�n�DXL7n����U�Z�ƻ��|�C�Sy�v������M}��T/�[	��q����E��,�$̋D�#�����å���z�]�"	^a�6Q9��G:��3O�*z`J!�05����HM����F׭"*
7A�5��!O���N�T������AM��P!�+j9&�{;@�v6PP%��j0=�6���E�J���}�\���Ѥ��+\Í *=0���/x/���t�O��%�M��B�n^���ge�פxy(+cq�\.	���D��NN6H�=]�M+D�%_���w8��1��5�-�n>B*܌7�(	&�Ί"���*c�m��F�
��]�K��;�M�QUwY9�;q�����7��G�Ú�Ze�ꦻ�}/�`�-��y��|c�>`'�e�E"������V��.��f����2D�y���D�U��[K �׿�c�{lϕ�Mڮ��.�
�?����[d�[Ro�b/q�KH��#����v�)�B��1����T�Q�G��� �l��oG2VEݨ�x�#r*!�0���S�������Ӳ���J��O��5v���|�"��7 ��߭2��KV����f�*�7��`��ꋰ�$- ������!dxE��Z~�v!�e?A��ub�Us�w.����9��k�
�J��������S�Jsb&��k����y
�� �"vB�9�Q�)�9�:��E��?�l�;���$��6�����a\���xaG�����S{-f�b�Zf�薋i}������h2QX��XU�53�H�e��%>Ȗ�������Û���Co�/��:_�����=)n�mv+�Rj�b.
(ϸD�����[����l�*��e����:풤�V}�[![�2������E�0���L����#J�_����ө�9���o����\�Xh��\y�Np��x^oWi�n�/X�7��=�[>��XN�=<��S�ɳ��)!)�x�j�Pz�D| �I�;��Pj�iЬA���Za^��Q��j��)7���6s>6�sM*�D'���K׫o��ր
����t��R���$1D���t���Τ�ל�����1� �O�7iBakͳ�0FCa7	I0<��V��8?8k���fK0◘b��Л������M�:��\���r(ť��_��`���C'��A�ҋA*{ý����s�����M�	�RV>���b\�7%D_8)J@��l��	�?�2�.�� 셨c��Pf4�3_-�
�d$@Ȗw1��� DK�w0��-	����H�N�.�  ܮ�����v𖉠*������ԴXL<9��l`�l�d�71��5P�#�7r��*bD*�� ����M�h�Q��Ǹ��_]��]��Ι�4��lԌ�Y���PYV�f�V������_a���:���^���֛�����p�X>�pyAN�Ohg�����|��M���"�!����\Ҧ�9`\����O����$;�?O��:�,,)����5�d��� �g��_���X��B[Ý�������/#CT��@F�����~�`��8�E�
أ2Bɖ1?Ü���j�꘨�2�J�hc"�X4��̭ai�w���D��0���ѳ�g�"��'"6W���]r���uY���&fi1��y�������U]�
�7��.�`�ӡ5��m�"�e�c�6���N����6˃F�Vǌ���g�n�V�R��\%f�،��]�Rw���mB��c�����L��i�����&b,lD��\z�(1?���5��Qh�!���ux�Ģ�ȴk��~����" /��&r���;R�r83k�$���XK��e��T�7�z�e�Q���y��]u]�R��l�U*kt+�y:���B��{�{q� ��Mmx��t2y�$l�w|l�"k,����<.��YRZ'�D��9�_/sMxB���xm��.�C�0�nZ���U�q�G�'���>��D��-^��ׇ��}�M��`�m�uKе���w�(� jH�-'F��S��;#J؋3�&c��U�(5ZPjK�%%�j�.DM��yKM�ArQ5� x�T`��"�p
!��Q���K��$4����&�	�@���㏇p���íG����|���(�EyX(��d9���+xEM�m�s�U6�>��Dy��ɽ�V�2v�tu:�I`�E���dѽճ�^x �U37Ѽ���[�vEI�P�&�쉐1�'���˞	��&�$�Xy����=q����O�	g��n[Xv-�N�����#b��"��.�B�k�}#�꘾�'�^a��Q�#5��3�B�>Ր�E��y�F;�:����)0�I��;��A7�w�T�5iD��ыk�:�������Z	�RރA ��^{��Y������I���`�H���A���L >R���v�������^��Ĕ�<!�`����� k��U�IɟZV��jfؿ��	`!�iq��?|^V��/M	��Miҵ�H���8�,7l��Ʋ� veA�:&Z(qh��5h��-/0-�tJL��u�ێ�ua?#�y	�<�w����t*,���x^�XB��!����OW��<��!�H� ���f�5��@i�`�7�b��+�8'$���,J.`�W�+>C�s�UO�5^ �6:�e�(wn�^3�V��A���V��7_�E��yt��IH�)����[�#>�g1:�<M�����S�⚲Ar(xL2�.���oC�{��1���4�\0d�wP#3���A/��;_,�愬i�fo���>���TNd�������耝!���J�>��S�����ĨUL!b5U�XiO��~�qh����8]�IW����^������.;������Gdv'��B���h�욓T����r���P�SR������3�ocVeT�`<���1��Y?�8�^��\Vy0��ik�ħ�ޗ��3�H:��r^���m(+�WĆG��3	�A'qn��6Y<�#w�66?/���u=�!�����4e�{��7PQ��J;�kv�L���C��e�B1`��k�~�u�C�����{��Gm�QJ�0��[9ZYCu:�Z9a
:k���S(�-��r.:6l'�켌/��kM8�db�쓃~\W�6T���c��w��vC縢�`j��^˖ʐ4\�F�g ݘ�R=�:��~�޺a3�Ģ���K��|ڂ�������D%��ig�eў��ц_��}������=�6��jM-"G�wQ�����[p;��k�CD۞�j����\䞙�Y4v��l��x���ӡ�����r!��..�H���zI��^	�WI&IjC�Ɵ�����s$|���,<�H��Ё0��vQ��ކ(XA%�<?3�	�$ y~hS�le��N�+���9�/� ��؛aӞ��#&m�����vuZ�&n�>,����d�/��^��lͧe�1?I���U`27q�H����G̽�_v�a9}��X�Ac�!Jh���O	��#>`�"Q�EÈ�\�����[���@n��x���{wU�~)�:H];���ҵMF:�E�R��u_eX�����I^��Kd�A�H	Z��:����z��$ș�=d:ʋ!#�So=�a�^~�^��Uhݦ�J��h5�)�.�����>�g������\�J1����yA�G�������/���K}�N����w�0=��o㱬��i_��9HD������UN#�b�m*<W�/��5fu�*�ވ�rb��@%�@;�J��h�/�ua��_Yp��PK�4|�gC���=:F�H� �<�]��
H�#�z�F���A�<�� �!U��(O��o�񏦵i��[���Wͧmw�ӿ���6�>�O^����<�c��0��H/� Gq�/{����+�)�w񄠨���'0�	��>�G����<��I!$��rJ�SM�s2O��$���ԅ�,����dҸ	��6/7a|k�����p���W񣉢+7m�u����e�SEݜW
��[��bPv!�Iy�%bi����;TF���SyG�{��L���� (�2bd/�ϱPߞx���a�v��z���BˑW�����kXF\Ïcx�P�p�x����X���n;	�N{
kK2l�Y�mX�0�!��@��/N�wrUqh1x|��GqJ�-|o�V�u	�FiR�C$��Z$��x
&Y��4���#A��q:x-1��_^��S�lT�d��
�+8O�.��^ʷ�&�̀4|:C�N1W"���O��+��&��-�������f!L�=� g��Ý)��B�~�?qB����3���_�mdL7蘠l�p�<X6CXcޭvÐ⁴�
���]P�x������qlg��ah�	�5�ۡh�F+|X�4��k��M�hy:�ݠ��'��K8��$QU��������fOn:C~�����|��ե(�k*
�u�g5凔�L'}�aHm���!Q�xz����ʕ�� ����E�w��S���Ua���Ɂ����R��o&~պ�H�w�!�,����-�x��"���{
�E�0T�S|؊M�@e��E��3�zF��:����El�'����B�0�u=���JC{�V���*�I˧R(���3j!,�p1�o�i���I�=��-/w���@���C|��H����avDl&�U�8W!z�;����ow%F�z�^ȋL�r|Lʸ���#��2�|X��,D'M���4��d�n)h9�bO������e1$$�T����l��-����mT�5�7Y�'t�:}�Y�-W��S}�J2��#s�/�YƤ����&z	�&h %W��"��C���䁤k��;�`�-M	~ Eԛ��a��j���H-�Y3L&%����Hp��~'�y�7vu���7�G�\D����_�3���e�+�x��#|,�Ǫ��C���ԏx��3�/~��e�L$ǯ��Wen@�j�Z����_�,D��5��X�~LZ"�$�FF�g:�
<�^Wa��3,��)(D��'' 3�ҝ	'�e�ᩖg�x>|p�D;�k�)�πfIj�;�"z!�ep�b�M}�U��Z���~��TC�㗚8���}����p��$8I�5l�l�����g������AE��zL����f�3oS���U����w
M�O��D==ȗG�>�9n h7����u���U�&����a��16_�amiX��@dY�<Va��A<1���������p�Jx<�X�b���Ps�c%�<x2��`����|�FF��yB��A�'R"Q� }��2�+�[ �����E;~���m�n-����w9�d�C_Q�r���mq�R�ax��E��|ua
�G��군�:���ДzWj�1��4؉����X���</��]X���-0��n>�4����^�͎�v~Y2xW��������a1�ua�7����0ĐA�/���[:Ӂ���+��y�ņm`�g��7h�
`�=[*nKxɂAm��qB�1�Hc��Z�T������)�n"�%�ʎ��dvo��ۤ�yq���)�;��&��Y��sXTcG�,�Υp&�^��u<C�I��qv��e���M+h'�b/���>�Q����ʷ��Q�*��Ȁ�}2�$��
�y�����B�}K�k�Ġ��`��TYs�6m�l��ʅr�q�_�%��s�9Xp�/����$�Q�&��?{����S7/�&W�Hݔ���E:^�]u%�`7�ƻ/U�1� 
0�U�����Τ&�������%1�Q��b�������EVvP���/NJm��� p���:k7?C7F ڵ�c��j #Q��.�R�8G�ɢjkK29	�~���תNF���ixM)rQm��і>��W��$+Z�����y"����ػ��nc��@�� ��:�_lœo�\\ڼ��'9��>I����T�͆&RL}D�Rv�P	N�+�ū�S�F9.���WNV��oӦ��XDQ����kE�F���ws.D"֐ߘw!��o����>k�w<$е�@�^���cS����d�%�� �� �R�[��#�Q��Y�c��c�wjꈺe>t�b}0ָ��k.����`NcE4��pc��d.
k�{��iu��ް��G����*��AA�-bt ��d�D��j�x��[zl���34�;��s���)PsI՜?v����/MtR����nVd,����	�_Jѥ ʗ[FF��py��6�t��sz �F"B�-洀�ŐT�;�>~6�I�,��j�m������%�>���*V�=�K�_�:�[�����&�H"��+]�?l8� 2���4���S��cS�"��@٢0���b�Q"�%m��m�@7=h�L�`1l��eţ��ߙ��Ԯ�R�#��[ ��CG��ĂH��s�!��X�.�ߪ'W�Y��'_&ww�%�χ��z�z�n��f��b��f�E�VN��{aIZ��+ډS�^ǌ������Ke��r���q�\ٌ����ܧ�Ǐ'�l�h1��0�^�'��r�t�v*V����א�c	6��K���'����.��ʵ�9����4���/�{��s�}����� G��Q1�'&͢�&#�"`ѣ�ݤNsI�b��A�A�Dh���po��9iqvLPpa|������o˖*O�t�B_Iu��f���.�~��r(6&�`o� ��C�i.���|��U�T��2�;��5��آ�g����7��Q�� l&�A<P�EuҕcE���A�hp܊��Yq�%��{X褒��t�Jg�~6�����7.�����U��/'7��`����dK@'-��Wu�@��k�s#��8�uԣҖ.�
��L[�)�(5i頓��ظ*U�u��Uc�ܼ���ʹI]�/�?�3��_�
�� �mIc]������=W�@��e���mL���>�SD���������
8Y�-c�;M�,tl�̟���x(=:F�P:H[�͡��.�/�<꺢��2�QEL@�4&L�Z3��'�'�s�N�+ш��e�B0�H�ã��Ry��{�/�}�NѸ���q?,r������hK�t�A�Č7������X#wG+�-����4_�uY6'�3tK_���q�����<�7p��|��[ZU~;7u�KG���[&���n4���;T
�	Jt�38�ca\V{��N7�@�|��)���ak�)Oؾ �Z��CMy� n��ķ�?Wb*:[�!�?U��)��'zj*�pGLEY��ar,X^�����9c�e%�����K�I�(��\4��A��Ր��0��gCX^ #�#� <3D���C����s�������,����# yu�X�l>7�X��)�~�-���On�H'9CbGG���6��
5�n�o_ Z�kdD����j	�~}��,��d�\����ݛ3}�JD�\?�D ��,��r�"�j���t���`�1JZ�\8"R�|`��-��<\+��%�f�5�������A�ƭ�ٛ��/�#C�MZ�s�r�O0:��̣'�΋�2�w�b{��ίݹ�1Z �}�žbj��)H<Уa"D�dٶ��S�l��7��W6-�^�`�<ehS'�Nn���Ȳ�iܩ�j��W�R�O��v�/y�(�?{�%ss����Lmz;�Z桮�q��1�,�`�.�3�ڗ�8K����}$�.���0�;��RRU'��v�t�C�E	�
8q��i�w��׀�b{�X��l]o@9�������Cۄy�1f�7*��+��N�V& 6���ς�#SU�uNI搩��v �G�E�,p��Ѐ�ި;ߒT�_�c�~ť�Z�W��O�h=S��猐�B�~�l�Cu};~V�Żޞ�V��DaA�Z%mA�%�4EH"�X�<GQR~҉�s�(���Î��:J���ʛ�g���T���c0*�܉�:�ȉj<}Y�Ԯ%	N.�&h_�{�!g߄�۪�}z:�@[��O<�V.|1��g_���� �0�35�E�u^��;t��m�p��?�=gJ�v�,�s�
��
8��o���	�S+�(��gE'd>��L[Ѕ�w�G_�6�8���ŵ�v�%��5�5����B�EM�Erq�T���V�,st��f��)'��m��<��,F6�׀(W�T���H��2B_O���@��V��>k���P��w�q)�<�i!��M_��O�B���ø�ڤ���Kh�E\�5\�s����j?rx��<�ހ~i���_Rp����d��3s�h���*:�FOYtN[Q{%�[r� y+���|,��{���F��cH�6\�D�m�H���_��`�@ �T�L3�xH��d�[Ɵ��@�`����?3za̓d횷�t�S�˳��kٙ!��~��K��`Ŏ�A U��gM�ZKDX�r�9p�_Ϩ���S��W�U�g�Y(�(�ƛ���)�"^]���\8��9��1��̽�Rjl'��\��DCk���YK��Ff���F�bkO~�T��u��F[�N�.mr����*M�
?�=X�� xWxߓ�^��>͔��l��t���2`�'t�[�L��r���\|Pi�^�X��l\�z9�!.e�k��o�;-���� 7���A�9#~S�G�Y����RH{���*����(H���V)���&:��@����)h��s���5�� �R���p�z�G�=����i'Nǲ{l�E���^���苖�C�	��S+g�D�w�|s��_ .��44��Vol-����u�a�+i�@����\gǁ(+�xcK�4���s�1��_1�Y�<�Z�4���Y!�W��0\[Ɩ�@gxS���E�"��o�u/��.��F�#ZD��r���T�>��������d|��(�{�k���E�_3��� ����u
�@�A-.�o=[̦L�e�D%͍��`�@N��cEKJ�Ŧ]\����Cm�]��{cvF����AL|
��������|�������g]�P�4�9_3Vv�,��z�i����F4%B�a��+��ȳY5TU4I�.����" �I��,�2[����E{l���4��{I��Ux%s�;Sk�(����!�%xc)�4���B1)��xmr���s*)GX�3����n�KH�
��!m���ili�І��0�Y ��h��Vqb��d�F�6 �'��1�k-���pkj#�W�s�<9k%o��~��>0�RdzYfo�P�m1�Zթ ��C�U0e&6ޮ@��FH�^/+���_+�d��<Ӽ�S�r�k��>�ժY��P�i g��CdYĎ|\�^9���BB�<��l��YW��{�0�ma@�����V�2���R^�#���\��Q��L���m����*�!l)9�dw>�3��Ӿ,<l�0����������˓O�:�[�n��������{� ��d�V7�ԛ�L�.�\pδg�ٲ���q 7xt0�kQ�6�]���W�\�=�%�Z��l'LW�X�b$񽜆����W�H����#���UЄ�P����l}x�r�+Q^~��5�}#�Qj�?�of�f���$d�mz	����H�ɳh��#� j�\���؀ת��\�Ĩ��fgA�Nxuۋ0��G�b�	�3�������Qm&�k��*��Bu5 �%���'7 ��Ʈj�QBuz`� ���t�h��ԂO����[��)���hxՖ뒆���əs����b��Rq�����԰��%O䁏��3h��d~���
��7�}m'��e�S���3L�*�r=�O+U~e�#Z��Z�^A�����V�nRuV�I�;A &@��]�}O[�Ԝ!�f��!�j��yK�][��G�u>K|��)�T�]�a�Tx��G�"8��6�*����`��21KR-ql됣2Y�7�������C��w�#���;d��/m�Z	���vJ�鈯D/	�˘-_���X}ϮV��lG��>;��
Lp�k�v%闟�j$�tG�մ�"��O�ZK���`0�)��y��z�*
��9�-"�7��R�nm���k�\ʾ�8�����>z�
�]�]P�+���4u�_jhu�1��_h���p�4����T�IQ�Z��{:HI�Ȋo��}=A���܁��kI���c|��$(Xt>�Z��qL�j3�jݎ� -(2�ǫ1��iN^�ؼI�U�'c�ub=s��)�"{��`�i����g|�>�)za�(���������a����5�Eg1 ��,i9�^Vcs�U�O19͝��H�F��w�c���:s����5s B���\�8R�� mx8IR�ES~(}:���[O���B|>[<"m������Л����+����M潕�1�l�	O�#I�h���+]g�^ ĨM��$S�	��	��
�Q�s�&&��;-�$h!&�����AR$̄Q�*9����4���U��!l������XM�%�n5��A�L�)A�}+8�E� �<�C��c��ʧ��'l��������8��pkd��s�e�V��^d��F 1���@`V�!��)�&vr�J�Qy�~��qLÿO}y��b�z��Ag1�z; ��~����Q��$#�����A���|���I�h:�jPv�H�N���{*���	�(�Q��i�U���Ս2f_��[ۤ�������&��ZK���[���q�]c�b�@P�?"�f�>�5��c��w��� 4�R�AC���b�]�2U�[�}zե��������\���ZQ)��CY�(���K�kޯ����+T#:�7��;?�~�������HO�����4�q��U�oW��E��E(��w��}e�x�m���Lr;x��+oBiB�=�v�%��}��?j0��S�eь�Y�2�a��>aA�ASeϻ��^����������f�6�*3B'�*]��#��V�9\o�
�O��<�`R�+���|Q���S���g �n1F��$�q�hm|�9}p%�s����c_d�=G0Q��j�K����eӍ���sm��bJeݏ�X���ŦU(�$���b/�8�V�|獫C�}�r'C� k�0����d����BP�<v�}{n�IČg���g�R��3�ZDLlg���&���ܿ`��7�k��/��I�B���~ӏ�W��KLBR�eR�G���0�ɇe���E��;[J;6ϲ �r���M���PB��_�i��H���pھ7��+��Ɉ%����\�]f��̴$~Oa��3uB�o0��W=zեS�!A�+4+P�//σ�S)�soi��o+�X��Y_�v��\�8�tc|�xV�vhO;��ͮ�5�$c�?���=�C����s�2t�����5�8�� �g�B�a�Z�fi��t�~��R��\�%/����8�EO��1�я�]ڪ>�x�v}�ȃ���5��	-~=T5��w�p�'l�-%F{:����hF�Hh��4�l��K�����텤s���:�5��-C��c�W���{�5��@ǟ�BI;d"��զ��K���x�*K>gх�g�뵯�.�-ή�Y2.���V�=Z%')�'����d�üqהּ-y�a�'�h@Z�
��$-���.�*	��0���U>Y��zP@!��L�\D�������61�&����#ˌ&�$��X�Ԓp���Sa�)J1�_6�ew2�[`��J�2�>��	��0�)]��G�OMc�d�Q0M~:bpb���#������\�h�c�
�r2e���Zf)��ߑ�3�9*+oB�򱧘�ٶ�?!R������a�i$&�.~���I
=���.���쾜^ح�2?��Zk\r���,���4��t��L��M>�ޏ��KV����4I�i]�ص��N
�T#�6�;cuX5kGmw�]��Vb����j��ś�vV$&94Y��bP�Ȼ�wc�!L0�ϝ��A�E��T@�X5�;3i�E��	�M`��P��sC U�N�z����~�z/t�0�}��X��~�ݯr�YQؖ"�K��3t��԰�}�|��Ps]��e��T6?Gd��9�,����y@̘,�%߉����;ͦu��
�͍�5d���l" �C"�Yo��,"�!%���� 
���#�3����1ԩ��8��Ӌ"1ڵܡpX���������YXfiw�r��B�h�Bp	T�q|￑����ޖ��n����>q�+�H1�����.'1�*�'އ� Hg驾�:����,l��:��J��f��ƿ^NS��:���f6��C7Ub�u�ovo��
2X~��(wW�1S�c ���<דg����/�_�4(�LR�|L��j8FvM�޽�ևm�vzl��v7O8�xV|�$�*�V;�ħ���Yەk����S��xx%�W�VJ��B��[o'�����Ӂ6fY�|�F���N��W�e��qg��f?!�wGR0��R"#���B?�%dM< ����f��zf����U$}^��	g�e�4jZ%���b��.��$,?�ˋcJm�w��lt�C�n��R zGW�5��mfz�6c���~�o����ٛ��K�Hg�1W�38�m�.W�:�pF���	���V��B�#�	1��"���Y�Do.,���I��,O��K#UvcyƱ7{!̥�U:����o����@�I?ɻ��;��~h��^�"�V�f��9,��A�G�ճ�B ��������>]?�"�9�N���yq��8'���٨����A���A&b�P	L_R2f/�?3>�Q�"*&�GՇ.*��:˸W����!�ץ���p'T�K��?��7�xRl���z@��Jo;�x�b�yщ�����/fS-L~-�tzg��һ_�����.a�a���К��uB�~�=�j����/֗Njآ���a�[T�m��,v�;�i�|�a�L��h���v������>�p��2k�V�>~�J������eK�8����}�C#`���!ھ�4ƕ��x}���,D	�!��("��ƬX��.:h;�H�0�4k�z�D.cc�^�N�'8:`܇gb><_ po�hm�^�A�Y�>0�8�|��s q�B7�G�!$�#jw�ض��g-9��j����p~e�hd�r���\����,9�d�>�'�B�?|�u�
�&�W}��k�[�/(�RB�6�6�q��.���u�gc�4 ܮ��!Hh���Wm�R-d�mbWW�(kה%�8�alh���D`-����w���3l���i\��W��H�J�3�����X�Q��{b�I;��ug#��͙��m�-��
�|�=���	�Л�P�;o��w�QP�A��l��G|Nm-��޴
y�Z�j�6I5r~���S#z����ɫ�^D�|�Q@�:�!��������\�@�YT�]&[�"Trֿ$��w�g���٦5q�N��c�S����aC������oT�m�8d���we@���������&:� u��İ|N_��M20G����BΈu����OYNƯGf�H��)6{�C�+C�D��*�g��Ծ�pٙ����,��O,���z��lOUő]6*^,�x��N�+x��|�o�^�CmaX���7BL��9G�~%����H"Ͷ]� �1b|Tl������xԌ��r�Gh��ߍ���d��R%+VE�E��u`�J�0hb�
3�s�m?��N�k���&2���>�W�'oڎ2 vY�r=�a��� )��P� ��5;&%�r��^	�5�>�|8y�S�P:�՝�p���Α̧[=��'x41k$��J���Չ)S}���ꯙ�< pF�ɤ�ìU�՛3��Mh�U���PH��}�.�n��8Hj�c��*#s�b<EJ���|��ܓ��wՋ~v��
d���0�΅�� ̴�o����$��Fw0������L���u���h8�"x�Q 5�E���Ή�j��%dvBm^��R�~�Μ�\��+x ��s�yr-I�P�N��i}BU��W��H��y �D]��b�����%�M����-���/��>k�G�	)zixBƓ�6�>Q��"/��ʩt���fW%��`?�������Ǣp�o)��+�9~&�ޓ���h%��B'�8ZID_�7�c2vJ�UF7���CxM�-��0�`g�D��(�}��Wg
���Qk�ʼzh[�9�3��؎/����]�׾��W�KGEQ\��m_�e�|p(��p���[�wD�	��UQ��?��ϢK����W���@Z|�k��a�$�Z�o���]~2�AS�<led�^@%Xt���u��ꢥ.;+��i�@�d x`�~/<`���qɂ�}�O���t=�m�D3��轸�-���?�/��hHƲ-��yjk�l�;��'0��U��>o�������6j�����Jq�|�z��A�V�K�Qt�����PqyV���F��Kd����,��g1^�I9Mi�Ҕ��22	��$�e����k������PY�)֔�^$R��Aq����\�3�ܧP܈��߯���~�3c�M���`"���ET=�wW�҂��E݋ݛe�@r��QAT  a5�k"_�U��eV�*�^=Gw��9h�b�����a����c�$F@�N��]�.j�<���Gn}}^k� ������Y���#�������cQa�!W� !$��:�$�*V�Y;���%���1��I*�E2t�C)�1sZ���D�� � Rk�1� �HL\
�.��#�
��
Ȇ��e��jB-�q\J�ז��^��w��a@�0X7MA�%=¹��C�0���[�������0��@�����ڸ%�3�8����KĖ 	�-��~Ok��9hc�uD�-�}�G%=|Z<S�{������b;��B�7tkg��:IR�����]�x�>��8C����:b�pn+8���o�`�8�vF�JQVv�r�Gْ�ňW6�5���\�M�&������E7o��}d��O�KCJ�˿!�z�+��҃�UL�
>N�n}q�NS%�]��!�,ԗr��!p W�/D�Um(R�>2i�kz�X���J�?1%��uZ0O�/�`�ԩ�'����mx����yӶq/��I�]�3��ZE�7�����}�uϦ\E���L5�t<��k�'�F�|rۅ�ȓ�,��8x�8�yA<4�D���z�ȇ�>�״ϴ,��EKm캎e���ř�9ُ�C-�������8�R�븘t�X��X@dͪ�,2���S��z�{<a���o�x8�a����2�v؝���d�e�冃�Bۑ�8n�Qb��G[�;�Q�2J>��&Ö�׬v)T�	�ZaT���o8 �geO�U���T���j"9��s4uN^��+���Tߐ�~À�"*VN��BK���J�`m�ތϔ�FB1f>U�2߇���V��3�s6������DQ�%���p��f�n��{n׭0��gD7V�>�����B�W5�9��M�ڴ�T�C#�:z1"�39�\(���餔�� ���>J�P�V;����c����W:�h��;N�����u�_5��}r����)�1��t��ó�{S8ڴ����v�>X7Lٌ����!���@n?�pΉ�2��px��LI�+=͠���P%�K��K� �r @�H��B�E�F�A��]'Lk@����`�2���ũi8&�v�93W@G�X��P�e��SO���Z�׻��joAbAz
5�4A�9�r��9T=�ٙ���gL���C��\?��>z��O,�[�������w%���l�U��؀��E�|�����0�+DS�<���i�c��U�~'��Ƒ���i���@���+C��Ge�&�؃|��@�I<�)�3�@�Xbk"a:�N���Q|0���!
h��r�������x��ɰ�p��8a������L���l+�@�NK����Pw�)*2�u�����\�
�b�,ٔ�qh0����bt��|v-X*�\�!�B���K�#X���\�ȻV���{�#����[��c�{�OE��G`W��>��EeL�e�3S�Ljp�R(l�͞f4����t��1��'��a�?�Xc���L�L<��'<�����tH-o�9yߒN-9��U����R�e�S���0�=�J'�b�2:�ΰeu�;|�Wq�~����ޜ?����߼~��Z|Τ��EH.�� ~}̼#��`�J+!�'�ea=���yv���`�z+�L��H��ĨC�w*bm/�X:��"�N7��eU3���g�i�)�7�D��}S����z=l���Z�u�׷��|c-n�偽c+JI�w�G&���iJ��z�����\7Q��0a��8{䉖E��j�T���>Y1L�8�
3k�^L�!�7~ ���/?P]`,.͓Np�N�k��o�K�z48諺�&�n��+�ʽ�xs����Cm!�r8u=ԗ}BV$<:j�&����V��En:G�)�⠍���8u�wt�40y#�u{P�um�wȫH�ĭ�F��3�?�O�>�B��4`AzO�#�F���MǷ���e=E��5��s�����9K���i��'K����-㏕|��E�������K��5�����Ѫ���%3�MOLa����Q:J���W_'_�/��Ipn�hgWTp��r>��� ��!�k�n�ؘ��O|��`�X�-����|�b"հ	�;A��Yw���'p8�Us�|(��L���%����/������QC��S�e�I��q��`� t9�#�����f�A��s( ��P�t˼���!3sz��܉4:]��5'��D�f����#u�r���%�
c�0(L(��s�ڇ�-�M���>ퟮ�E�M��X�l��Oh}B�*�<�SJύ�<.|�J�?�Ѷi�Y����ع}\�i�{`Z���n]��7�@TW�l>����戧ݐ�`��Q�2NJB���Ҧ�KR��
��g�>w�����l}��c]jCQ����VI;�E�?D��|�%کy���__P����g���=��w]�d��x?˯��+��k�o�����kC��g��f����t��A��I���E6�^Ջ�L���x��9L�����}_<Q�}d�O{g������kS����� "ff�Y�8}��آe����h<�T�ưN:�������3˨�m����Q�����+��7ne��c���
����ԎF�)"O��U�z���h rQ����_)\�"�d]�9�Yi�EV�|�uם
�L��Siύ&u��g�<K�A�X���1lw�ݪ]�.<����Oz�|Ӊ
����Zuvؒ~1�� $��LM��������ǩHn�p�V"aW��u���J�9�3��]H�@ҹ�-����m�]~�����x�Cvy�k,��R*
dF�z���ǟUe���X�v�"�mN\����+O��&ا�po��q�O���g�q���v��]��+v�O��n�q�����F-�3�D�-������FAW�n�����vT�@���2�5�M+�(���w!��Đ�~��C�P��k{1��J�K�����w�D�k��K#?e�`�YXɞ$T��&>� �v�����g
'���o�5�����4R�~ANFob����Q&���,�4NJ�bv�m�+�b���P=$�+�F��[���"-׾ory{��m���sr�Ω�ĽB�&��-�S\�BJl���,�
�II����V��d�u'��R�$m��Z?ቦ$��QD�w:@@��p�띦��Ф4���;�7?��3��z�Eհ?�S�I��˴H8Y����0��� !�{���WK]�F��-`����I�8�#�ν4��}2xJ2o��A���J�.��,']:�Qh5mi��L+O��:v�.���*o����y4S�]ȹn]f��.���&�_t��pb�A�J���&��_�p� �6����y��17�W����֨����/�X^��#�lHm'kYa�ך�� \�(��/8��5�]n�N �a�GK����T���y�z8�4A?)$/WQ�����:/����?Q{���t����R��ύ���3��V��}23J]k 1讏a���<�Sb5���0Y�f0�ѻ%з��T��~��;�Ĝ[��5Z��y�A��{?flW�AIb���&`@�"�@��NT�Ty`/@�'�d���JY��T����,U��� Ai�̟ߒ��%աC�őz�إk��X� #� Ie�e"�Kt\�z�M�C�:Sl��J�3�գF::�Wa�^qr�����p^�;-�-B�	D�0QF����!�H�����ƻ��~D0�5���	ZF���d<e�����K���ۤۙ�� dOn����Q����~>;ށB����7["t�[�?�
T
�y��aV�X�[/�<ϖ���[�1�, ']ͱ��)akf4M��%3�I7�y���;��ђ���n5�=�N��1ZW��p"������X�U� ^,�
S�N����y�UJu�n�S��������#	�k��F�����n�% 7F��P�~����t��|�����_1=}K���XB�����e�zם�ߨW��?��`I_h�A�a�S��T,�I��fy� v:�P(�5���B+Ա����5�*��r㟓׏lr>[o3���.��9@����7�%{>�����VLG��&d���NMF��Q��@�̜�0b��袏 M!�*�.Dў�Ot[�Nc�sQ?�7�w���W���GhۘwG�������{T^��u�L�^�l��Nks�B?(�P�v�G���,�F73q,ZǕg�0;�8 �M阻��/N�����룅�P����ԫ)�;�h��)9����.�fއ��%���v����yNx\�0H]��sU���������=�q��v��;��r�W�z-�YK�O3G�*y_��ttw,��'���p��MѬ9�a�r��2Vͼ|�����0�]*Z�E΂��_���y���v��#9'���Ks	�XW�y�U��,^�|��|�N�&_��P���{9�0�,�Yap[�e�� QU��gE��Ʃ�4�(��7�{�ç1���Ă@'K���8�u��ŉX[����-���W�X�p�=S�w:�ڔ,}N�v ���+]�j�F�ۉ�|y�p1"��l@򦡣�}ɠ�����x�����"��U\(����C�FJn���6�c�O`��w`�骏�M�����<F^]����`mh�ۣ�V���dm��x��iM�i�,����ȉ�6V����L�oݔ�*T4f��;��<V��?	p�#�u���>��s�-6��w�5-ܶ�'����X��:�<�Ƚ�� C��0^vJ�N��vn[y�e��I0t����-Ҁ4o�1����P��e򵀉i�9)r6(�	Q-O�l ��|��a;��晠'Tf+"��ki@'r�U�[0;���i��E�JD������QZ
Q�y	�<�*�,�+{���*�/$�p��X�D�k�0��
(��ԑ��ŌM���?���@�.Ψd��b	>����´wZنX_��Q�D�x�͕�"�� �b�?E���_M�� �/���_��}���eL��p˕*�5�V_��)�є�W���f������Dω��W�)�'0�~�X><q�k������	�^	�i�*��m���V�j�}$��
eb	Z7�����r����9x�P���γ4e��+B���L$��<�@�3E����ؒ��,U�J ���/1r��@�$�-Bs)k���^����uN�T��Pdox��z����̮��Q���M�(o��Ӥ�E��a�2y��ć)��_I �	kX��F�S���q��_�{��P{�m�|V
��М��0ȥ�p�Y�d���l���dӐL�0�n�#X~��=����Oe�̇���0%�j���ↀ�Zns(��۱b楒��~�����E6R̟�$۰�P�Ϊ�o���,B:����N֢'�����a�:JŨ�R��r�}x�c����Y�
�i���+�E��:��H�GbWtdU� �y!���+M[��A��"�%�X��v�o+l�'v��vd�����b��{ǲ�ꄭv@�ۛ�m�)V�׷�(u��	��W��0�U$K���cr�jsU]n	��hl%++:�#���6T���s1�<mTJ�v�P�M����gi�N�B�c~Z���Q��m�5t��K������K�����ҹ2�mc1��������Yt�0�p����a�"b!��UZcZ�,��_p�Y0h�	�j��ʶ� K;m���,�鵟���{��ڙ�L�&��&���)�3��^�cLi���Y�T4.��0x���967v�
��0��A^P3������꧘[�u��dC�3b��*�(}i������W�LQz_�$�#�B��d]�`�}&Wi�(��e��"C�b����	`n%�@�䕍v釟͔���BFK�H�IF����2t-qv5	�	��}m,t[����Օ[V��������`C��z��ű/��P9����	mwK�OJ�E+�����aLhMĳ�ͪ�����؍��W3��9�c<��LI(`Ea��(��M"�ggD��0j�����\}7Z^
��s�&?�d����J�%����XP��?9��Bjʠ\�q#��I���\F�����/I��5�tw�N�N�<�T�G���&�n�DE�!?KϚeRwW�E伩���w�]_p��>T�i)i��G*��G��E�����ӛ��q���X��U�/Ԧ����IH�N��[�HN՜x�\%�L���NC�Qg�LYK.](�S��1��+�ĳRw`0+Tw�Ob�P�(xc}���_��[*]Q�5�BЖ�+���a-��"�sX|�#�?��"4 �~��b�0���j�|<�������28˭�����ۅ�m� ��離	��u�u��+�.
�m�/��U�j؟R���A3�^�m>J�ɚ���7�Δȱ�r{�,��+�l �����ˇ3"�՗D��@)i.uŌ�h]��hq�ُY_5%�>��Ĩ�ԕ�.��HT1!JtHY�	ૺ4�0n
�������v��Q�GsSp�ȶH�����S��5�C^�γ�79?9�k�����{�`���	��u��ˣ_��g|W�<`��Za�=�~�?��)K�r�Eld�Ay�.����&G�ia�5e�ѕ�x���G,� f�6�䫿*uۃ�y(�Ă
gD5��!{GR�N�YV�q�Ui���4H�p5�i��<�ۇ��,ikt%���_��c�۶�a�
�>�����tW��;V
_j��[�_�\��X���@}v��aa<��}��\l����|�,֏>ʤ)x�%�O7�b�őG
-�Čt�-R����+g����typ.��JT2j
J4�#)'�T]\q����00�"���2c��9h1�0���xx��V1(8&MY�d*�9Vh�� 	E��D�������d����5��c)c�3~�0�Ѽn���x��@GXR��f�'��|և�o�t��֨!����I늛Ǯ�@5��ۭ}�ǃ�@%e����.�]Y�3P�����^�5ww������[�i6�G����Ν/YT#0O<P����cϹ�Bg"�RU�>?��
}	.�`Юq<d��.��1�>�{xp�ׯ'a^ˎ�}Tx����f�C7/B��!P�}�ɘgZG���p��[\�oƞlE_�\���4�"3&�6�O�S���uKtk4p4� �o	��t���˒�������q����`2m�������wa/�������՗K�%`�4.R�|�X��?�[�?�-�c�\�Å�ߗ2�)�V���!�T�n0GֱOU�Z�	l�UŊ����*���������v��C�~؎n��.��yE*96�}9
C���^,�	�k��W���<K���D�%��J�fJ*g�M&A[�} VGZ���8:OB�{���K��&'x��Tf+�L�v����B�^rK���ν�/OݝR#�a-�j��tݥ%�ν/�c�������̞�Q��L�q���\�\;h�v%	�3��㢪��x���:�=� Բ����X�CCl���|���	y1R����5L��w��c�~�>t#S<��b�h����]H��2���z>�bͥ@����v�` ����2e�2�����6�����Y���gn�*]ݕ�hУ�Y�F@�W񟑡��]��;�Aʫ�t?����v�Z
���5����|��U-��%8�����ћ#E�b�V
�y�Ӂr�)_Y��#�� |�~�26��B��s��(���ǆo�Z;z���\'(��#�0lt� ZHq6�è���̚A��)b�yR{��|zf!��B�U��M���d̝T'RÆ�����ycٗ���g,�v$^90E�%ۤ�k���tbd�"_�,�QE-��xYƍ�:.5��j4�Q��^j.���{u�����`��S�����~Q�ʚ���Â�ѕ�)�܎J@��z�&��T���/��s ��۵.r���eW�p�Tɓl�x�9T���PV�����鯣�=����Rz.͗�*Lp����e3S�k��QAU���Bs�d�ge�Z��|�l�l߫�i�+�' L�s�#i=*���n�*��n`��xAeXI����c�'���5��1��\�q���GQ-(��?k�I$vr�,�O�ɂ��b�%fD0��3(�N֋ ���ݥ�T�/]��=�`-!��;��1\����ճX�
����-/�>7VL�Gz_W�rX��n!V�l��۸XG��k+T�vwPg����n͜�̦S_c��0�b�|[q����B�5��/��S�=E����	-���<�.�h0�w�w�	t8Պ{��!e�����x���ıV[kw,?I|D�����F����e�՘_(Yr�hWX��S){^�<,R�\��|=��X$F���/����cM�k��y_E�]���p��B�%#+
u��w���Qޯ[ό���i�8�<�!���|�xyuT>SF�Z+A��!M�|�Jd^ٯB�pn��3���������A��kS��e=��v~�YN��n��U���H����F�~9���4���R1����/Ε��W���t��!����g�$J�?{�o���Nۭ�>þ�x�5�7��'��h�\�g��E[�>y�]P���zG��>Q��O�m���՘�v�������i�z�bL��C�er{W4<���	�~^����{╻pV����P�A���cK_��Й�"�>f���,,�3ςN�n�OV$t%�=^�j�@��%��f2x���aDy.(3%'��\NR[��ņ�P�CW�+�V�f����O��w��c�AJʐ���X�~�+��A�y�ٗ{��~�O�ȟI��|�s�o�ؽT�f�m��ŋVI�	s�GK�Rɦ||�?v���LQM�>�h��W��W�'U���?cZW �&�J Ob�Q*2	ɞ4�xHo���2|���z�b�����\"�yVBͰrNEܖ�	�;�_�]l�w����L�R	��؏{�J=𖩐ꨜ����a�A����*�	�}A#s9AC��@�����R��j�Ӌ㮶ǚq����+���ϰ_��o��8G^{��Pm*��@?��5� ��M��D�|��ʫ���u�ҽ�����fPE�v��	������w�`�w]�Ƃ8�#�r��__�z`���e�S8&����~LII�,��>.%�#�(F�U���0���B}�r}an�2����uRi�r�v�25�b�a�1V�	_�F^	��b�u��ݸ��ҥ���w��e������1�����@�<�>5�RpA++�5�u�b��뜓h?6�ۑP���$�{�-��Q��2��T^F�/p�|���ށ��L���,�C.t(�h�Y��t�K�����5<B��Jѵ�V[�V���F�)��p�*���i9��U&;6����b�R��.@r�8;5��|.��t0��#K���|��iҊ�k|H�S&�F~�FN�����	l������~�1bs&$�/���A!�7_�'N��x=����� ��$�5���A�U�t艰�jw3P��ކ~�0P��4%��~�:�����^&�C"G5U���ڡʖ�tb��I��5I�Eh�����ڛ,�_��6H�>�!fBݠ��2Q�14��:&�dR�1�T�E �&׼�������=}��T��H%+�hs	��p3�_�\�;3���; �����H���6N}�R����Q���]a4��19na
��[SE�}��i]��s�<5�A��`��繬?)��Ð���B����{�|�|fz�hd��8JGF�"�wjP/�/
�8B�2�h�qJ�

)��^��V�hʜ!� ���O�Na��?zKЬ�ݫ������I&	תi��@ʹdoqg�_Q����R�~���V.� ��G%÷*y�Y�P4�����}��Po�_�(��% ��%�c&63�gT�F0�2Zpu?S�}�pZ�"裚����E�g�!��g��&Y8huW��A�ȁ*Ӈ%�4�/�"��P�g�Sd�mP�@��T���hIL����|J��0���UVh����78z�\7ݸ)4I�|�&U�4+�)9ZD�q��L��N�Z�5҆Rc8�xɜ\x���5--���H�'�dIu�.�1i��:n�U�C��X�k��]Ф��yrj�S�)�����mJ��n�S_&Kq�|8��9d2�a�g��ֈ��wK�`��p�"ɱOY~�6��d��'�a�uS��@ZZ�^��#�5�����S�����������A��i�N���0$s��x�,�SjQ��6�G ��ǼECy�s
�|�N@�?>��nQF�&`��3{�l���q�tm��Y��(�26��K쯿���>�PW�!��<C_� �Bt�������r�J��a�@�.�SbcNr���A\i�)�Z�:��O�lb��d��X��vUYd"_�fJ�!^{[L�����D�J�Ѣ�"�/�,�?I������M�� *�f��T�d��y�g�4��U^�E?�~'�[A��56��ʣ��GK�U#T�W�3����k�3�?v�3��*9U��(,Ea�N�-��b�3;�-�^-nBwh�]�-6�!�e����!�Y#H}�Z��&["��Gc�������)ր���v#@����q0; ��JD�H��>���5�2?��(E�u�
�~���@�BF)�����}sI�T͎Edp4+gL�B"�ā��A�HR�Svm+��DH;vMs�4q�eq��s�^Q!��kC* E�Ԣ(-8�þe+j�`Pq�T��O1̟�r�^�&lc�i�V��Y���x��-�$K�6 bJ�
i��x�fl��Z����-+<�ސ*��m������-ߦ+"A�qɭ�֣J��!�/W���ۃ�¨Љ����jAPy�_��$��P��W%�Ă$4��v)r�xfb�zz������։i����kn�~9�	%���Q������;��!ۻ`�|���������]s"�QB�7�	?[٠����Ɯ���<�{S'���lE>|GD@"��X��{��?��,p�Cn�%u�˅�0�,�Ш����s��b{�m�7 m �=yB�jT�\3I����82!��CŻu(�t����db�����?�,�)<���I��7�\^<���0�����˞BS�s�ϛ�K#=��lIy��Ӎb�]�����PAEo�_ڡV�%b263�����ă�_��e��Ρ�uB�z��I, 	~�3> ��*����Q5��~���w�(؎$��x+�C(���F���m.��ߔ(�C�a�Rz�ىB9�!�q�����uG��t4���C��Y=�&!+�$��k�V�7�-���x�uVڋ��2�GXO�1<\0h�v�<����8��Ͼ�P��GE>��\�U����>l�|�VkQ����R�4����TVS(�%L^\��L��N��E�.<���1��>A��O#�������(� �:0�u���6��Z�h�]��-��Է �2�a
`0���~�o(��з��w,<���Gu�sy���}�eHw�LUs���P���6Ԣ[	��[8�:6p�(��۳O�Y�~������_pĈ�͆X�.���8z ��Un�1����՘�/ Қ��G�+װ���e��-#W6�W��M�$�T<9��+:���n�c]j��!J�Ǐ�/)�����ə�O0St��C�p���4F���-���\��G��ڴ��k'A��z�ο:���,'Mhq���ݙ��S!����܊�B'ݽ���?PO��|m�mô�����Se:Ȋj�ψ&qc��3��8S$�x�y�AP�
�4������UY��ۙ�XL��(?�5�BWV)��YRsϱ鏄>I�Cb���;gm�W,�Z�ޖ�j�`,��ڃܶi��9��	�~�!|J��	"���9�4�i�*����l�P�8�u�u��?��;X��p�~���~{�E���J�m�݇|;�C�gTz�&��KRz�ѱO��� ���M����b�I��)�J ���-�����aۀ����:"�T*��F�.(>
p�+�-V��)��x��h�c	�)<���C���ej�:�G����׵SFǺϛ⠁sN�uaoq���`R��(lX<*��=���C�����l�����ӡW��Ǡ����{�ݘ"���j��>����`�s���5�*h�1��C�1=?��V8��=�k1%B%F����f�I�u��6��L��_g�ۧ�%q��C	���]:�<pV=?���a���!��
Y���~"��V֬/�d�{�꜎h�h�On�m���=c['��{��Ŝ5�c��]�F:���/�����i��m�a�l�r��K{Y�4GO��+Ӧ���f�,W�"$J?�������lſ�8���<�b/O���M��`��{۳P��,_")��u'�e�� WFK]���z�u6�-���^���<
�Gs�����'�����������˪P3��1[�-<-�#3۽��3�6��g��}�|�z�������iO��M0<�h����nI�/F'�R�W��!7���o�}]�f \���6�qftF�CY�*A-§�᱋n4�t,e2� =4��� ��&��������ꙺ%(%&���hs����z�@�d��N���c��?Ti{$��n|XR%���O��B�-S��%�Jq�6���1�F�*�O���~����Т8V�iU�'W5�A��91�B�YyRyFMӪ�z��T�@fZ`����ڱ�4T],�|�ڐͥ��(~��B1��T���)����|hd�����������G,u����Eq�$�)��������HIY��.X]���7+�ȶ�NFP��[�!�x2(�������'d7�
4uk�=7�f�_�{tO~u�z�݊�?��uE�Ig�Ȗ��QZD���X�d!N��bdy��z���/�݄��%)�����˺�OTc��!��� �:5��hn��A�t��H�X�o�;�c!ʝح�U���`��$��|$*�
f���z��[��(�i� ����g�W���i�2�����=��	f��G�����K�D�5���zc�����R������Q=x���9�C��}��[ ����t��2�Kg� ������ !t@����2w�N�����`5m}
W��eiL�*T��݉�8�y��"U������\�yF�,6���ۺ6�doPkFpeVK���QUBd�T!+��Z�����pL�N�M�#r����W����0*�@��=��U���u�9t�����
�"���A��{�����j�C�_��k�7Q;�v�Jh�+�̍jxJ�NMl�����	P�a��&��9sF��+�"����qi׳��k�r�Վma �0�&�+������T��Du��&-�`�g��B����:T�F�4,1��za�R|�����B���U�ӓ�˒ŝ�y�7��w.��<�W��07�����J�L#[:eZ�0B'ˉ�E3��~(�Y~5z��
>������S�o��AU)r9�ؤ�@�c?���T�h  5���|���)��作��:{�,��@e�}��(��V:��;�yz�10�J?�
خ$J�8�k�.���w�sm���.�V��b1�(�)�Ņ�C�@v`Q�\@ݓ}��ҽ^s�>��?��B��g�|�r?@���q)B��Йa��4�&(�QI���Rj���6��@�h'�	w�=e�4�#��SV}�`�Z�\�(hR�Y�84������x�*�PᆗT]�P��K;�[��3@���h;k�$�Y�I;�Zƹ��*�"A�R���Ʃ�V?�1��	��~��_ܽ
܍ �ئ&��4�)r����ާ�2b�+��/h����֞ϻ!2��O�:�XMW���#i�l���B7K��鲢[6�9=1 �W%C�)U�+�b�r��hDfAqB�����G3���)��9op�ͩ����57�K��39�U�������̂�i�����h�[&#��ޠ!`#+�ĀY�s��t�6�-h/��!\�p���7F-����b�ȥ�ĩ�HESP���1sS%I:��h١�� 
^��-]3����
ٺR�}Dj�,?氦�����nT#���	�,@q^�H8O���:mT,S%H��a��93�2FO��hy����uϸ��V����@�.�t�orӿ�k��sN��Ԍ5��b1�E$S���l�Y���B��f���&J����ҧ���@�#.��4��֌�6�w�(t��������zs �M��"&7riL�^Z�D8?��6��,�*&Ñ�	�׌���r;��f8T�RH���&ѽ��YZ#9�o�Cf�?/�|
9W3��1��3��j�e��������l|�F�6�:�L/	~d/��G��h;����<I���[�gi�ij�Ȇ�O�,��BN�=�
�b��:Y��k��B�'QoKu�E<�̜_���h�4��g��ܸ��}��y'�mބ�%{�^$5�E���	���c�bqVT�������{t�u��?�GS�%�����5��/�7-�f�Ez��H�
Q-M�<T���b�G6]eS��$�[<�^�;����h��V���P�nw��a� ���.��@�/�����u)uHV,L�!�4���_��P�81dX -$5��ƻ���P���ڿ���RʊA������V�:������M���[�?`�.-�S�0
}<������6N�M�g�X
�^�D&@Vk������j
6�ԯ��d���R�ݮ��t�Yl�V- ����J (��[1��W�i=L1n�2�t��s˻�T릳�yLP(ub��ःp[���\��gT`�����Ă��~�m��S=,8���D/�s4V��6"�@c�%�?q�ɵUJ���\Ǆ�n?������ߎ�B_{9�ȴ�<]�m�\9���UB]�G#h��)d%����?2C�5�"�bډ�N�qP�:����:eaδc4����#AjY��q��]���Sc�� �-��Ք�]�p,38�4W�.r��s�' 3Q,��ۀ�1���82%5%C��nY�Jm���h_B�_���?�&7n���겭�����ݳ�{cҜ�fn��|D�o�g[mk`���!~�'?�2I�G=/��vk������Ý"�d�&"8��L=7�����?[���A�fo^�_Q+�_R�<��8Ѡ��R����jrJ+��r|���}3b)�nor� <,��;dH�q����>����?��q��h���j�n�J�������atg����'Eb���=%�5P	�EA'G�(w�/����M�&)-!5 �57h;��J��ʶyb��n�i��46�c�%5C��r��T�����\韝���� m�@�p�5�����=+�ZP���R��&�G�د�(-�
~<^zo��KQ�Ć��Ry֯��R�ʇ�:Æ�����9D]Tf�F6��!��1c�_��z��
w���B���q�m��.o�Mw���&�љ4�Kq��G�o#S%�]6�^��;'2[Mz	��:��ځ{�y����JU&���;�	A��<ڷ�Z���o\14�g�~����1���^��1ܻ���Ϝ&����@]�=`>��iN�����K�.r�Yfd�Cu�PZ�r"o�׵���&I���.<^�vݴ�4�l�������꜕�m%�Ĝӊ;�~�4ѩj�����=�G&T��������#︽G�,��y�n��Yhq]��P�l#uB�Ċ�����r�i�c�W���\�.�؝G���=�6�eƸ����ҙ��殂t+��1�7�����>���\ <!��5��'�ڐn��%9H��!�	ޥ}V��,1#����4FF3�H�po�Z�fΐ��$��a�i��t+�#�d`Q=Yuƃd0SO�a>�;S��ej~L�	D3�UĄ��U�W?4�/(����Ģ��\N#�,���k�u(Z, 7�&�;��?'D��!g� ;9"H��B|���z�Ԩ��9IsIwY�:�j"{�nֽ\j�����3ϯ����7��ΆM�(Y�O�5+����Cϸ̱���A��t�ҭ�9DK<�J�����R�B��l�N�ۤ.Ь 2:Ck�m�{>Gb0 �s薎��x���ַG<���� `Ӱ���V�a�j�+�ŋ���Q ��6G�Zp���H�X�4���b���O���di�L�[�q{�l6��
���k���s�Y`���#�r��ۯ��>�������ZQ�~,U��>��'N6�'�[Y���'}�
"Έ뱂�\�{�:yfu�DRC}峥g�~S�(�J��  ��[���):�����i���ٜk)Η_o�aI���e@�&`�1��7�=�����ڕ�M[����*�X�E��u_�J+2S���\���yР����͐�;�ϠP�lLt�^�F�(��F���� �o�����^A[��O��� �����cS,��樕1r�۞�B��������p��R��7ޟ*F>��s�ej��JS��O
 E.����A�)EH����?L���]C1�^m����[�f	y�d�©O{��ş�C�1R?U��akȎNV	6�Q^ʫ~�'���A��[.8S͘������~�T�4a9�|�}�%v}/p1]3sy2׈d��P�¿���=�5��L�e(�&@zv�9��n�Z���*�ۧ};}�����d�4�q�8���8GP�L�����NezB�1)�E�O��ٖS"рf�4`�����~(���*k�e|$�$�"ɫ����/���+�n6���@�Pʯ����f_��UːU r 9WD9���xGf|ٵ'���V��p��V��<���/z�s��t�g���������oX	��Ի/�L�uA֙F�ň|-��՘r�&Vl�����G^�H�'+{͍�F-�{U�'o8�F�Y��kV=}{#�A���(u�ďng�wQ��L�!��4=� ��l0׈���ǹ�N�^������pAٮz��(�7���d���
^o���Zr�rIW1'�?Y�_He�bY�Jڮ"�a����s[��['�_Y��T�l��<y~-u*�pIۓ�I>�3����/\c4�_��nas�� ,׳�OH ���a�]���[Ăq2Cj�ϖ�Q�QAyH"��x��*N��V�[u~�x`u��@�R>�=��qg�![� ��3+�Ng�l�Է�m�:В4���W9��F�KAɘx�3��z#CCʵD�&i��RbnD�ڧ�m"]�ȩ=� ~�*5i@d��a��H���^5��qh��6����R����`I�b׍�q����sxҕ��a]�,��	T=�s/ry����D���\{L����,R���i?j�2cR�5�1��@m9}�u�2�r���Ws���m�f^��wU	�z�b�#w�Tɤ��udz��/c��ҟp��Q��9�n}�ٚ���<`�Pwa�5���K�GEm���{��)N�Uea�W�!j��a�Ё�8?!oBtp�l5qA��A�S�^�
Lqۗ�ڎq�
�ޤ�= &���^�\��B�.M~����Q]ev*k�ݾ���0#.�B!�Z�ag-�T�#�|iN��O暽>W�ܦBp�_����H�9C]���0�w[��^���/A�]��d�ͨ�"B�����)����߬��H��%?ͷ�0ܘ�G��ҥ<�.����N��d�#�9"V��Xe�.m���9C���sz�����Qu �~a��Z��X���l�C�F�r?FK���D�Cw����q6�Ls�h8�1fl��E�(!��$B��ь8=lx���e�@4"����E�RWk|�Y{��ƌX��ԁQ�}{�Yo���+vu��s��<�3J��дo��CP�K�C_io����?z�%�_g�CӦ�*Ni��Wu��1�B`�J� ��0˭�4�ߎ��{h�z�Q.$@�}�7ט���0��!�vz�
s���&S�:�7��� (��F�N�N������ӭn��G�sh�ȭ�^%�6�R
�;5i�c�+�#�˳�0�&0�CP�����;<�V�q���	㍫�в��\�ڿ��U~��K�x0�D�:hk�	�����R�J;�����~�G*	!RP�������c|W{�|g��F%ٮ���}i�ʱv]?����8蘙Zڳ�fa��g�떬Xc��I �+�5=�K(,�"���V&X�U_��tb�sI&M/��������Q��-�@��d�<��PI����;dY<f��?�,���j��_�N �-a2`�t/��iT���KL�8�IֿAs���}�a�;N P����юp�;��Y:�D�%�}=�β�^�ɚ\1l[8�r!�]�g2���'�,g����u�I�E�K�'	`^@�0jCۢ���Id�&P��t<Uq|h]wCPզ`7����wh�����������P���n�?m��m�np\��#��2/e��\N��*#�AZ��!&�:�F��QA�6n��;i�yD���p1ص����B1p�A��pv�S�'�a\��AK��3�f����g���uY��H�x������.+͞�7����i��0ɕ��;�.�j|���̴sE�u���($�����߯D�3���ExK�X>�����jvz��mh8����y]��'�Eq�9xp�Mz�xe<]�q'=�KO3�E h#����+�m�-��׫�>8��ȕ{�܆�=�o�-Ң*c�ep���_�	���m� [5��㜚�C#~��Y5|H��ZQ�E�<���%Y�<?,˟P o�N[Mq���?��<m�eɴ�,܉�*��*�O��O��Ke��$� (SlM���ܟ݁�i32�·S�Pl餈�S���g2!i�K�x��h�� �M-
�~v.���L!2����Y����㳰���Z�f�,��-D�߁��~���:U�H,L~5�63���#���e_��W�X�sXQ��p0��,�Z��J^����H�%��*�Í����Ktun[ ��(I�� �k�^%#YG�����ͼ�� W�)?�������NM�Np­
�5���(:�9q��~jޢZ:��tx���+�G{�@mB� ��\�g�r� 5G��T�y����X�fb�����q�R.�����`7En�� 	.-�Ծ�uI�u��4�[k���Rv&s$~�6I�S����)c�c�6:3���}HB=l¼����]d$D�nFɄ�7�r~�,� 2YM8�~��Ө?٠��u�Kg���E\��h���)7>%3R'�Ru��#��@���r��d�v8?�.��ш�J����,��\�T��/���^>/0��(!/�m��:Z��b�5���}D:�<����}| j�A�|�d�辯f�BŸ��"X����,�p���?ݞI+r�ūB#�<Ā
}���Zf�武(��ra�.�����l1ե��,�F�Rg�\�S�����;8�����'�Pʁ�:���WSa��,�J�W����0�#����S硭���w�z�,;<#k	l�{�K�2�@"Y��OP���+�*��p�yGnj������Hr��z�iCg���E[��@��[X���9�-�Màd��m*X{.�;�ѽ}�T~H]Wy���+w�x�<�)

E0ի�iz�;W�U�����_��/��2s���-d*]p*�����_��ج�
H�	n��R�1NI��i��"��1�=��J!x�q�¦������|G8J��5a�6��C���>)�한�!��<�؃�M�Ǜ��|��OM�2�fC��M�4B"e+��]�o��t�fE������Ԫ�!5����'Y@��L������a��ogvk}��k�4���%2.�
�y���;�t� ΰ��	�7���\6Rj�';߾����M)�d�v�|xp�^Wu�O@M8��9BN(1��o_G���q�9~N��|N�Nw�������`��`�)�SO��t6��Pމ#�tfk����i���!��6��/�H�_n_M��-W�ɋ��D�x�35L��"w�����#��>V�*�����kGC'��:�(j���p� G�I&�q���l+hX��cCxb���Ҵ۰0� �w|���$�h��8����Y;���@h<��uӪς$����7i�����Ȍ̏w�&���˫�Zm���JQ��U1{���Py��33$s!,���x
_���	�V��Z� �m�"5��	���W��<����I@(����ٮ9.D�аm�U���Y��ҫ`�R4�����{�ߦ/`�Jbo�����#m��Z�D����]��F�K��P��TCzxhФ�jӾGn
{ۻt�?�+)�X�d�0�'D��A9�e��5]�� ��nO�o�F����0
��[�|��?eUM�>��Z,��\�<�y�������wbF�8GB��H�z�.|Td9��Fuc�D		*�_�����~�I��K<J$�꛴J��x�\Yt,�$ �+�|W�i�%��;Rb�^�"ȧM.}F��2���af),;�в{��>!�:[��9�
��;�я��	_��O>�yiV6��x��ck8)T�"��qH%I��(/�|�PV��⪹GF,����/�*l��%��_�P*e�ԅx7h�{��cb��Pu���g�}?sϖ�A�#$�y����x"��	+dD�uW�Ż�w���Ji��@�W�a_�m�'(�b��4�&@��bӾ��sԁ(�).~���͠JÇH�F�Z�d���Z�{���,WKX�V�N2��o[�\�*LP��ݒ�}��j@��F��&������*��)��ڗ� �<��<wT
��X�!�xn�V��d��9�d���7A��(t�5����V"̧�U��^��LE�4�5�c���E�E85�G��� #�Fv]Fg��ֆ��/^V��^/�gv�Z|/1v����R���F��X����(��P�_�ݻ��ܹg�4D��b���B��R7�d�f�;��Yt��:�1f��fv4X	<��~��ݟ�ˠ��>F⮵��g[�`�L�y�g�ݷ��A;���6���e5p��tF2�q:�c��n�m�h<��Z_�v7;�@w�ԕ`���Zm�^�:$w������G��_m��E���b�P�\�G�	C ͟
ތi]���o,Zk�F���V�\��Z��v��3T�Đ�(�8�g~�̎
�4h�L�R�~�$�]���<�C�ɺ_�79���-U|�F�`<6�oUjr}񉋺j�Nc%��_&@%1#�v�j�M�N�����@aȪ��P&r��?l�b'�Nj�Ed�R��A�xFê{4��1��Ê.�|�׈��9r�$���8rRne�]����-K!�M|����
�-W���A���Z�����o�JQ9�4:�D��L�M����밣6�I�nkaJ꯶���]��LaѫX���g�'�g봚i����I�'4��1�{,�X`A���Ax�b1�L�O��r$&�������2��+���>�]A�8��1
.UD��fF���]�>j���y�ʫ��@��璺f��y�+�?'}�u>��|���p����&�=U��*_ߍG�K�^����'��½l�Y��~���wk�����,��!��\�.-���B�K�}1Nפ�\'�K�8�g*teW	#�W��eʑBw:��'�f=�����i(������͏G�(�5��wD����i�����x�a��z�4��m��-�
�'�R�2oY ��<(y�{���F/����`�S x�P�ҼWQ�#�v$��YdX�C�{<�,z��+
�H�K��^+�g!�3��eъ����\�t�b�*��{�YC�I��py	7���y,�+�%Kj�n�޶d���oK|-[��u�/ݦ/r��&[�+fr�J�̚A�s��_Qى�O%��%"���1���\0���~O1���O���ƞ
�^��苼�
�,���3i/�ܖ��.I�4��tb[���j^P�R=?����*]�|"�Ac��E4߬c�iHV����!��`A<wxko�R0i�F�;��aX����3�qO��7DtG�c>~0�����I�e�2QJS��Wg��g'H�/î<T���Wjo�\뉨<Pu��%��nN��:��@�Y��A�H^�#���;Q����_��0ǁd6�f�a�c�聦{ċ�w���C�b��9�~Ɔ/2�TO�����?�T��#��6;$���lb�"� �˪��p�rF��j��x�+5zP��ԫ$eҏ����T�s�U�n��Ԟ�H�v�����=����� Wb_�;o��Bn�+\E~�������s_`j��z�7�=������{,���,0̢B���0^Bi5{���_r�֞�K'�ى�]�2��c�L��(>ru&���J~�)����<���(����:
 v[AA�z  �,!�TQ��aѢ��/��dV�^x҂�S�JEs<1݊o�fH��Jߢ���Cﵭ���_6#�T��O�1�W*��� F��1�㪡{!��3�h5QƜFB^e���OcN]u?�m�TS�}O��Y����m���2�لu��"�1}�޹��f.z��T+�H��
��a�/���si�>��om�JΑ���6���6=�,W�\{�-Y���~��/�;����}r���v�]� )��@v�;��#	��� &�
7�-<�S�-,;J���R
��7G2Ǳ�H��9f�M�O�y�(��pP�bXk���L���a��
.��#���� ��]h��@+��t���5�&xɧ���(SR�$����Ɇs��:-70��@���fo��G�1�8-���;t��(Ǚ�55s��~�i�G���A�.��=��g�#M�=�-��Z��Kf��A+�h�I�@Y�������X�7�c��7�i��ݴN�y���u�W7��~æ�T�Un��%���y~��cé�L0ͭ+ت�2͑��?�&3|���om��~-<����R�|W��LQr�L��P��z�+}���wՀ.���f��MϦދ�"m�����:	WY�|�(ܸ=$��yׯ�B��h(_u����s��ڲ�d���;�T>
/���e����6��5�M��:�uOUI�Ƕ���@��tg��07� y*���������9��U�VR����p2���]����l[@��4A�2'T�Ed�t��7�J#%)�#Ek��R�iO%��u?��ؘ��O�������ca��4^ikG����>��N;]Qo�3��}1}�b4�K'���Nv=q���/Ԗ���7�<���������������l����oq`�U�?BK�7�?�X�=�@�I�5~J(C�X��ߗ\����%q�	�9��Q���J�Y���b)��[�m��[�op��um}!B{�w�cb"g�|$�j2^[?����?��'��-ڡ(�W�;�քh�l��t�����6�X[��������Ҹ������G|�2)l���]��L�}n��v<� H�C���ڰP_>�V�a�����D'yt*|�H2�=/�5����8x�N���Yb�! �ӆ�@q�=%�k������O�ϧ��@}{kuז;���1���R�1T����)Ap�F�Q�R��wL�8�4z`��/�x�n1LI^����\�k6u��B)*��������}.)l"��K���S!q�ַ兜?m�X%U����5Gjjߜ(w�=tv��R/@�]V2����a���Ō�y��l��(�H��BT�Vm1n+Oh���A#��f|q��C�%�}""�k��E%Er��ޡ�Ӻk���Z���qw��s��9��}�~|,q)���"���t���2�^�ê|W`Qe�2p8�8.��pξ�/��6s��J^K2V�;�	>�K�R�r%kGj�xq�q�(^:6�0.��B�J�\�ʇB�{�$;%T~�W(0Ub�0��E��*�ql�WO������aY�n��_�*��p`��BIo���+�#Mŏ�n��-O�:�Xky�'xtq�qQ<u" D�Zӟh$ ��d����d�EF �P�.W�c���2Ͻ�$���ᰧD��	"���s�l�	����{">B�jc��O<ԫf�4�ˡ,��P��8��� ���.K���ԯ�N�1�Y����G��ɒ5u����}��%�r�O��-��Ȼ`��`�z��ޫB���	}3�r��CZK�I���6��\:���$���'ǵ[�E�w�a\�$В6��N�+q����
|.9T�+qY�خ-���M�������+�K%��o���t�F��8�((MuA�f�����\Kֆ�GP�RG��=��!�ӛ�ѐ�]?�ƶ�hb�� 4����x)c���.sTi�x�v}*�2Lz�w��������d�\h�=���N�*���Kt#��r��_�9��W�Eۓ�����x��)��Jꅥ+M�m��-C�3Hbh�0*�%������ŵ�+�b- ��q
m�����%ض����nh�=�!�VU�;�Z<bo����J;2F�bo�3Z>��&���.�X9�~�(�5�SK�Fh�$dN@}zAw�i,k��x�:�B"��	e�<-�H��S9���Җ�-�V�l0A���?��a\���	k68T�%��һ߶���x!�r<�u��ؗrt" i��"��Zv�������E�"����*,�U�������v�gy����̛�_a
Σ
�q6<]>�~�aGńt˜ ��2�������P �5����M�B*è���f �ڇ��9D&�X���)-�|�4�u�
08*�k12�w��5�N��=Tٖ)KgG]i��-sw�j����M*m��Ȟ1<���T��e B༆J��c2�	���hLZ�$�vC �M66���N4-9�=>42˙�W���bo�kR.���,8��b������_ҹ����4��nγ��:�D2�����a6��'֭�W���|o�7}�b�<�C ����ѣ�[��M(mkQ�qoA���Y	V1T���-��*��P�KJ��nP3�.�HA��
�0�	�({���vM�;�� }�7���f,�u��m5�����#��׈��$�Êy�6yє�K2���E+��؅�Ja��u�Y�{�9e/6���Ƒ�B64?$�	�̊�Λ�A�5�A��L���c���)>�pk{2(6I��
�P阠t�p�~�!.o���N� ��C�����H4<D�����"(�Pm�XA|v�-H,�r�5��3̾��-,}� ��Fu�ˈJ�-���h��@��WcF�)�F�!D}
����$���L�� "�>޵>��{�ظ��b� ��!��(��o���[��ftĺ���|y��IV�����n������ٌ_�*`9W�E��gF��&k�j�
7d`�RL��nJ���hPH�}�ʞ�ڨ\��^,9��k/�=K��14V��lY�������U. E��C$u@�x�b��-Zw$(􀏴q�h�焌�ۣ�Ϥ/l4'�t϶n6s�T(P�14�4���Nؕ��ŋ2�l<���� 	���e��֪u����QT'�c�. �F��Q��y��pv��Ƕ�
�]'⎵ׁ��,�����ۈc��y�l��T3`/ֹ�
�	S���f?�D��Cן�6�J�����qb��k��W&���ǖ��Ԁ��ڏ�@�h�L�8Ӝ�g���~�Z$3��I���Y�as�\;���)��!h.���mC��$E0����aBj�Oyym�9q��_����~P�4N�	��W��%�a®��*�;hG"$���~�����-;Ƽ����}4C�Dz��k���3�̍�)Y5��
���å��	�t8�W��Ხ�G�(SK���nט�S��:��7���Pxe���b⤻���/LiG����*ӝ�b�Tػn�D��%\�L��}� ���N�Z�%9+^A2l�a���`�L������8����p��<�����A�k�wS�Z_�<$}H4�N6�+(p���HW��"V+�l�5'b�H�-��%�z;>Kc��O���_\ى=��t	���M��jD-G�U��u|�H�ă\m�}Y���ג�TgQ\Ìx��_��)z��6�z��uu�?w�e?,�;��̏���^������]9+�J����
g=2P�]�7vM�J�EX��[��:�@L�DA�7JIB`��D�]Z�4 dO���#o����:L9��ۂ��N���6�2p���WF��V�Í* ����t
��>s��\�^<����,�ktXM�[�Jv�f�����'&i����O;�aNta���h�����9�5 r��5�E%��pQfM��<]bg)�[h�C��.
� ��%`��|%�p� L-������@.-(,�YyL�?k�鵲��^�W�)
������5<"]�����r��5ƕ��b�d��1߆�$,���L�ol���Hd(�Fԩ<�N���8�8�y�(G�LH%��H�,���L2	]E��Б��O���}��뮅�4����{��݁�
PX�`)Ǔ���M�C݅�NS�W��G�a�2�9�Xc��ҏ��رa�o�PT� ���\�x��ݥE�IVi��m�o���0q����/Rv+�MS�6�JX�O�	$R���>���Ʒ+l�է�Q�h�v;����_��;:ml@g�?��F�O'��.UF�i�ꄵ�q6��*Z&���bya��.@�`������\�!�HL��ϻ�A��@d~uN���ƛP�u)Ӕ+�u�P(���nO�+G�7��*m@�@�Qi7��R"(@����%�͈�T��l�����[��8>d�9�&�5飂���A��y9�͝#�.��*e*c�ʊ7�bFqv�9�g=e��c�ٙ��N��_-q��T�l��/�RRSA��Z
�͝X+5�RC��/-@q�݆��&�tl�[�hg��P���?
[��8�?C�\�����B�� �:m�>����6� g.ǧ���b�GeP�xC�8�nҔD>���X*<�QFY {��Uj�J��!Q����<x�B �x���=.�$�3�^�F�nbm%w�B��*���n� ��b��{+%A ����w���In)QX��� �I ���v:��Vل�ډ�&S�h],ޣ�{8�l飩�7���t��, �p�;��K�-���N�a-���٭����}D��[�MO�A�PGʐ���'�� <i�)<�%1�~��P�=��u�Q@O���w��rf9qQ�q�״!T�����*�����s��K���7ܫ:�`w����^:qN7k���jFOm&_a^ �qR;�)<S�Tp�x���t�
N���н�����P�<�����07��jI�&��iŹ��0�ܼ���Mڎ��+r��8K�L���N@Xl;�ˮ������#���Ҫ��������V��pӏ�\9���0Qڮ�{��ɉN]���T�wl狠�c������� �M�{ �	��т��;�k�1WP�]A�p���IvH|���r]_Q `����ל*l�4���_5!m�/�.����#S��P�wa0=(o�����K��C�����4J^z�l<���WLS��P�g�h�׍�og!4��|C�2U);#�pȓ�z���gE���z�,H��\0��)��UD]�	&��׸.Zi�Ǫ7�A��<"y�Ec�.^pCI���fq��4_����E�Rc�ɚ�o�2@�v���+٧f�x����$oU�m��ϐ�>Ϫ��LHj�3>�A���y[}S|�Y�)�%�C�fp]%p��?#�E�a���R�*��I7\ �a�b:£��{�漇���n%������^��]�����OrnQh� �|8ќ�pr�hHb(���(G��S�x<ծ�����Tb��z�s{0�+PP3���k�Q
�qM �����a#�H���>�˗�=�7�G���}��l��!?�P�D��;r����5{��eHi� �w�@R��(�NP(N�g �	���"͎�1m.#<�)�ſ�!���#�~-,a��Z���28���H�k�`�q�0��#|�\i2DYP�ha\-����JDoh�E�h�1^��4�rR��L9U�Ǭ����I����%ƣ/�%DHy`i�A؀�}��T-���ϥ��6KSv���A�=YN721��X�k���W?�0��)_O�箓.���d�*J����D��ar^�� 9l�N/� r����jap�'x��ؑ>���ck�!˨�m|p<��?�|�Os��,uJ�_�v5n�سV`	:C�O����x�C<ʗuW�Q3�$��_��g%�u�h�j&ꋓ����;Һ5�1o�|jY5�'4�|`)��R'�A�٢ŭ�7��0M#���jbŞ��?76�R�9_m�`�� �������S3�ڪ����M^����m���Sz��N����U�V�x���:���5wZ�8�FN~��_��Xt����^]WuTw4l�|�I^8 �4���IoVN��L��� 8J�k�`S�q�7{�(����T,�qX�w�ĻIҥ.kb�Ԯ�W^�Z��Y�/ً�E��zkń��!M&�Vh�#�o��ا�J�U��5HO�"�d9�ܑ��<���["/�ռ���'Ӥ�~ V�&W�B��=�tL�.�n#n��\�z�;X���T�yL����N���� 
�^e�V��~�{Y�o�2��h"������c*���WL���DP�Fw�!�^S����4^z�|��@�'�O�| ��^f��5=${}��k��\�No�4��X� U<.�j����i<79O%;ݬ赚�_Mw�� C4�(�3Y�U	D��H[\��V���"�h���������X��VU��A>�g0�(J�T���U���������&�ŧ5�@gۨ}�؂�Y��6̮���"����������Ҫw��&�~y	e���e�|b���q����"��SI����5���4��(�OQ+�c�+]�q��fd���D`�����q�3^��g�x�{����a�rΘ�I�P�'qD�:b\w`D��u-���R	�0<��Cq?aٿ���;Qi����?�uA�[zO:�Q���=f��Ѹ2�!9�����Ȅ�C�˲�Va>.R\r�X�3���fq��dX i_|6���+�UΣ;�o��UNiso�;�ʰ�Y��]yɑZݗ��IX�QlL�7����p�[qz�/-�>��[�ұW�ߢT.[sU���=R�O�CO>�[#�0�'�{��ۯ�t� �(�LC��qc��Ju�D�hG�R?+�*��j����b��g��F�e��'oNQ݈�+��m�� II��̓`�DXlh�B����gF�hZ-�C����3M�/ϡOy*k���N��[q	u~.�߀E�ZYu[%+1�~���q�ls���W����'3�
�,��%g;'�[b�%�]=���/BJ��\gJ$5oig�mv���#$�?ԧCWМ�)���N�g���I�����ӏ���XVV���,; R�T ��v�S�����ܓϩ��B\{�Y�AJ�_������;�i8a5M�U�<Q)v=���e��Z�X�NT��&�Y�EB���̆ rv��Rr�T;�:�5!���L��T~��s�e� Ɖ��j�57�M���q�ƻ�{:�&p�bǇ�����L��{�/��TC�PS�|��#]����ė��:�¿J��tQ��5'�:Q
�)r}������n�ip��Z�r�>q%%���li2z�B�j	�C���]��^�2^ĐL��#����"2r��]��3bsV�ݧ�Od�x�	+�������hJ�n���/M\��R(�������ܼ)�?C��лw���r��h��>_F�$�$e�F�8[{7���E{ꭻ+Fh�#y���%'K�(�0��������m�R�gE�W�OLբ��}�0��)�����F��vPP�����]��r2�c�?j�"�X`l��Y�;ñ��꧲�נ��/{u�M�Bֲm�����t�K��q��4j�e�r��f�z�� Er�]Z�si���Q����7��ƕ�3����6���`��?`;�'��~��[�}�v)��\miph�Th�Tk�-��s9�9��
}�F f<�_Wܢ]�h�;ۚ��	�Aq������T�a��kcT�P���:���	b���B��$q7���ýk�9��Iq��sT�AX;��ԅd/���d%L�􏬃���
��~^�ب�,/�K:�.V���I+8- O�Uv�'m�^П��ߓ�[��6�m�# `��1��Ǣ�ϰ6�4�d��*�mu�Vm�W�,n�/�gyp��D�98�K7��^��i�}�΅A�ҫ�+�CR~�O���g�H)�U����Ś�!ѝ}����#�e�>f  ���xz1����^��Dw%�_�����oMU�km��|�V���o��%�y����4���b=��|�b��G]��<@OϋO.R�ˠ�-,HN��S�̯�����>�wʙ�˚�8����m�sZu��zH���r]m��e�o�ζ��<�Voj��OEC	NWח8,2��U1c�5���3%�=D��X�ݿ����Q={��+e>�8�<G'��H\�F�;cC�ܱ��P��.P)�N+�~�D�Ɣ3@�����4���Vp���b�`�����5��L�+��)�����a�J�������Cg�;�D�2�""7f]H?�Ĺ)���SC�X�>���)���eT�D�ma�����ڙ38�7���Q#[դ���-D(�K���s�^����x��04��[s��[���4�!D�t:i/��|��@w&i�Y��W'2'�Fٙai�5F�d���E�-7��7	H�' G��5(��c���+Eʾa���jo�j)�L_X{�M��q�s���Ig0�������H���o�x�n-�H����}�=�t:cad�	Yv�b56���^�wu��jx�r����X�?��LE��p�8��
T�n�z����C�8:\ƞ�Et��Vv��6����{pzQ�/B�[p�ƅ��:��dѶ�H�?�>x�v^P��[�o}uy�qC�8�H��aш�C�+ф@��,�;�(7=(/bg�z�8�����1�jH�9N�ȁB/�E�M�Q�vC��s��dFn���j#�\�Xx��S�Rt�M`9<@��5?�_6_(�=���5���t����83����+��5�+Σ����ق��@��Ō�q��lo�B����)|�m2�eJX�/��x�vٶ9>�u&�r-KI�U����u7|9"�Q�?�8�����l��yVFb�Փ�R�e�N�i��%t�OA�5"�1tD%p����d��X����,�l����;3ܕVJ�i�����-������~�!Y�׶��TfQ�#�m0x8���~�~/���1"fsh�PO3)� �/�/���L��9�;Z/1t���-ɍ7�%p{����j�O��V)��s���A��i�T���A�T�ٱ��|Y�v%Yc��
:��V����V�p�������T�������DrΤ�юP�*nc�*���`�O�l�XvGn��$𾽘/�)��O��ԫ�?ܪв�GUǳE�,�x<e�N����T��0�R��k���t�_�x�'�$�)��
!�9Y��R�"��������Xhv@���hx^�CTp"]���,����='��Nt�������Sm� m�ӗ���3�=�	�
�#�S��m|�$��_�S�[`��g�	��6Q]*OK!����˂�S��zQ�����0u�ܲ/���8�PDƦ�yQ#��<�C&E��J�7�,���l7���,����}�\��6��ӝ�il����� &�^�|�P�/�o�i�N��l(;m�Q#t'Q�?OE�TGͳ6�+��j�u����fԙ<�ίPU1 ��zl�|g��h-�@�}r|9��E����S�|e�H6`_A���L���=�_��'�������TL�^X!�O�y9V@�T�Q�Y��=�\ƨRTbH+���9��3�^�W[p�rjg���K6��U�T��O�5�'�k@���V�J����М�|rbf�c��a��L��Į���0}����x��Nߜ�7p�T<�>|0�5r
�O�A�t�M�$���=�b�a���7uM������<�k�Ʋ�*k$7䣤/f��l3���m����3����l��@N�a���~����Le��ǒo���:U�6����!����(I�Y{��c��ڂ ���^��+�x	<���g.���I]]� ��f��x��y�Oon���?��w_�o}�j�#���;��BL/�$[RF�&1��=�K����W��&��Ƴlw&�C�?���3�(1c�>�o� �%	���=�}á:��t�B����ڋ�y.B�	����I.b��3���mŤ�d�/��Ϗ*&ǲ�#|���t"��,py;��?�4_�`(5��_�>��h���2TUDs��y��8r}>l�xDĭ�UR*/�P���<���zG����څ��SMN��d8�>0�����$XLNe7Dz�[�.�t3���c�� ��าe�yd��~����&h��r�
�ޯl6H�xkVv��yU��Ə7���b�4���
���N�qn��k���Y��S/�'��+�fP��Z�gj'���F��T%�UYk�2P��e��xh��wg�ǰ�r��Vx�Yx"55��<�K��<���!K<�������PT�_;�_W^bQl,m�l1P��� �*xX&D����^�^����G�7J	8��@U���d��00�z-�NO�`~si�!.!�
˓ʇ^�w{u�7cU��������'��.bi�|�)�z�O�����m��N�}�]�9e�ΐŵ��I���8�,̈�\� UX���V��(N�X@�@@��K/�wo�0n��7	�=����q0
s:b�>���R�Պ�d��\��7�)|	�)N"lK�2�HI2.�]g�~�3Xa�a���]ܘ���W?���K�7�]\L�GK��5��2���N�DAFސ���/\`��G�]�=��qg�yH<L,��D� X㤷�9�4,$Ë0Pfc�i�î8��:�5��z�v~��$[��(�D��$z��*�I����yw��S3��kryg��1��%�#}m�S'E4(�X��+!pe���^���oU�sdه����`f���j}"~Y���StD6%ǅH`�����m� -�^�Oz��o=B5�����؈)�I�;ِ�ǌ=7�p�g(p{�{�oG�t%l�^(MϱR��y���Tvp]�>q�
����nj[��(/�����K_�;��+N���Y,GEU��%l���)a��]��ގwV������~[�m-S�W!-z��������¥�|6~'vcV�,����2��{���n��W�k(��� q�҃��jX�;A��qx�NN|�rO��>*c���J���Z�C�~m4��?�J!N�	�M~v�����='���c�t�Q��=`��0$��vD�Y���޺��/����MN�|�80#w��L�[�h�8/|��&�F�j����|jK������$��q.����ĽC�Ux۹ ��1q���;Z�Z��O�,ؕ���m�d6���`fc˸C4����ЊQ��>��������/e�/���j��(�O��=�e�xY��ǂ2/���k����Ly��e�@�[�Q�l���!]��\���i�n�!�f�(,������m�h՟��r��AR>~�Q�7	i5�&�י�6���}g�4�"Lt�ա����W�;�w��l���[�BM�0n56�i�"��P(��x�+���Jٯt�mi��PV�Fk�#f��{*�7)ב�+��� �6,�B�����)��?�o�fMV|�x:�]��&h����&*�D���	k� Ε�qE�e"��LgڍJht�������X_��k���