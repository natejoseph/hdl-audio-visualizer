��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N����lĝRFĹfn�m'Ɗ-֎<Cɹ��k�M����u�ܾI���0
�Ѽ�$1u>���d�e�$;�P��U�i���}����ڞ ��%%7�0�{ԜA琪�\�:���j��'�h�A��J�7G}Դ	p̆�ؑ��7�=�5D�^~����8y�$U��`?
��P'�n�������3~����E,h�Y"�'!Kkok
����	�3��I\?��&p�ip������\]���n�J����E�+{�Dl����o$��P�Qk�������E;�Y	-�v`�Nϩ�j�|?�D��r_���;ͬ��;wXo3m�)�ҴS RS��Y�3��=;o���p��kx�&&nR�!�j7�S�:nX=���p������F}��˘�YW�0��RJ<�%R�+U�|��I������4�G6��V�e�m6%�+�$�4@Xp)�{�+��kNg�[�Gv��I���1v��.vN1O5aǟXz���I��[3`�Q�;Q�yC�=C��@Ń�=��9���T%�w��;�Q�YOt� �dz�f��Im����l�LIa�Z�x��d���ho��<r�7��1]��p\�1�;Gxy�VK���e������7������TA��J�9@��"Z������(p	�W��h�2X߈�J���;���1���[{TDgT���� �%��\�S��|l%�x\�}�h�J��k����/���y3r�0���yT�E�{������^�BM>�x�����њ�mj�����<��خq��>���S�5�}8l#��6i���Q�!ܱ�Y>��0�+����>Rlx��q�괼�{l���������B���vmTu�22b�
jb{h3#�گC6�3�30���볘�� �m�X�Q �Լ���)\��/��c�V��YK�Vi�4���3!Z�嗚~f�oD��?8���n1��R�]�t8�n������g`c��а{��Qk�.����jf/3?��.��B��ef�_�<J�"T�]��_S�Љ�(d5�~q�% _�H��//�2_��\��/�SN�}���=o��l,d��A�e
3��s��F�=D���� �l"ad]fZ?p$�E�_L�i�NV�[x�2#�d����q7���<K15�BbG	?�<��"�C��oݰY��~��4�9t�y�X���2����Jি�nSD5:��YB,�fa.�@������0�)���:*�D�����N׾�V���(����j���.y�	���r�� ��B�"��k��"�d��]hUo��1h�,���D�����Sj�q$�;�����Q0��RBƄN�ڎ�3����@�za�R����#�k{�U���@k��c��aa-� 8�%�߃����b
o"([���������:��.�Ϫ�bD8füS �z;��lݒnX̾�n���f"�Vi/�%�o��jר�j�j��J���L\z����ݛ�)ܠ��Ϫ��x'��,̂���)�r�Q@_#Q31�sJ����JVԝ���72�Ϳ]~Da,��p����Z���z-�&|\���踎�>��N�%m>�6�E�R\���G���#��*�\�n0V�.0�:b��䋢'���ä��ǝ��DJ�
Gkz���������;�Ge�u|��~�J�գ-�����;�r�|�yl}j���H��tgu�!�ஹ\��I8t�\��{�e���ΈYB�\7:��w���d#�)�?~�ňi�^�8���e��ѯ���*1[ٵ�t��%a7�-�?r�ɡ<y/A�q��eӬg��g��C�U����;	s5��dղv�lo��j��5��)y'Yx��[5e}$����m%�,��k( y_����!C4���V��K?�����7�WU@����Y{�ش�aMHSN���׉_0#���RS����5=��3)S�=\t8u?>i�:.k�5ʲ��7m��f��+�->[���C��h���6h幚_�oB*�L�> �%<�/�S��ɩxha�>�R3mJM���H��9���>�"���2����x���<;�֯��h
1����'xi MmK[(�Ѳn�*��M�;��3���#W��ޫ��S���/�.�5��Ca���(Y��!b=�bOm�op�>�xc���I�GDc�}�4�ʤ���̗j r*�|�N4�[�I�;�wĩ)7JBث���^O�W~}�~�$�c~{~��7t��D���Q ÜG���\���m`2�x5>��^V�]���������aCF���T�JDd[�l�����-�n��W|h��
)�ܠ�kj(�X��{n���v��''�L�w����IX���ļ}��J"��)����k�M0Q/�N�w.POl�d #��M(^7���N�ȃ�0����=S�{����hk_�� �� �����l���@��+���^£5<ˋ����
�h4�yY�9���P��3��Q���c�uf��Fq%���5��ɇ������S+-�� Ă�%{E�~�(e���%�{�#o�^*A��%���/�:@��u2�ߘ�ܦ��z�0��"��Ǐ�;%�>1�=M�B�S �c�g7y�#H��{��0,R�:#���yU���[\̑�[��X�ԐB8�"���Ìq�k�=��lj1�9ý�`"�����-���&E��8��1�s�J:6�Op�tUAF �ȃ�W�����)@R���L�L,Д	��¿��X��w��5xq������5�%2w�-[��`��%���qTj�L`���X��C���vP���!߾���x	w@�ۺw3  =/���8r��~��Tv��;��L�[iX���q�3[��5/-�G2�XP7İ}i9���z���������y���9T�����E��¯ �`	8��Z�����\7��X�`�*l�t�?�0�����1s�OBF�Q-�T&n�b��c�r~<�hu�ev���$em�Ѝ����k�I����������Sj ����s���?6� �}׺���~��ƃ����\eq�P縜q�~�Z�f���'r�D֭Y�ㆉ��ӆ�{�?S�꼩)�3rWv���0��a�x�D
wX��~`�~7��c��Z�F4:L"�w�LZ�!���g���,g�P�	ڨu�+{c���+�+���]�}8@3&�`M|Hop[:�/!������u/b!���87y1�m#Nں�Z�-����ps�W�q�HpgƬ?U��ŗh`I�ݦ����&򯛪�E%���"�-bѥF�h�;��D{���_�lס�i���� �(�gi�p��M��Q��GRF^/Yr�zp�?�l���(�C�v*M'����V�����ٽ�V�9�p7�%��oB�@AM�2�	��r�Ƈ����m���K���B7�p�+���v9��qP�)��>���W�H`�=A��F���%oW@)hw�|00$|k3Xuku���֙�/{�/T��F�3[���ȏElʈ�o(�<��8�9P��J�ͨL|"��'��@�gr��|��I�w��th0A�h�5 �<9�������a�h@R#�h���SV��e�D'H���u��������Ǻ���^�{%�]2k��wrmu��3���;YWi�#�(�!��l&�1�9Y��_%&�i�[�Ks7�JS�UΧ�N�X�$�a����x��i?b�2g��s��}�D�>��_�}�sI�q�ݓ6a���9<�7r����d
0N܄��F����OW۔
ߓ�-�S7�"O���4`=C<+�Xa��n�T�͈r"S�4Tn�\8�K+���8��f���Be18��4B4ht=Es����?P˺/��P����ݓ<�BY�Q�Ą|�hNYm���j�N���uĒF�=xI�Bh���Uc��M��K�v� ��w96[�CA�mc�_ Z�2�a&��V��KXB]��]Lh(�NI��b8|yܿ|N�T�.tpsZ�@��o͂"�zq�w���u_��1�Aq�{��< ���I�o7ȭ���� iB���Hȅz�륒u[XO��i�X�ȼ�8}i�7�ff*��M�,J%��G�^�*X�$;�Zڸ@M���r�)�8��S�I���,*#�PS��7��_)-��I'�R/NC�tz(��E�)?9�e⩁ 'z���۪���vYU��� ��NcE��,�H�#��xgG�Zښ�������V�����<F\�`Q���Y��0�����ni�UCi���_$�E�4�����.�-�-�%��}��%}���m�\�=�<M�ء�A�A��,@�`��6�QZ�0��� �k�ZzF1:Q2�d��稁�rB��ʮ{���*45"<���Kdd�O*�wᕿ�a��[hb/���]�c5eco~Ԋ��Hi����-y?��Fp���\ ��pw��Z��A�����:�~�L'�yV�d�%@�'�KD��H8l'�w�|Z�Ȳ�Wq�
s��?�9� -�����:͊�	c]Г8�r�G%���� �w���}J���[=����@�0���#aA��R�.#ޥ<��xF!ޣ,��N�`_��ѧ���^���G�t���F������X���w�[ꢜ���8=�h��j;44�/������'sJ�&��8��[CQ���p�¾��%Ǆp��ڋP�ke��ռ�]�$�ἨV�<}�V���Bx㗜k3')� 1:����D�v���Z��-ۈ�op�_������B���EJ��Y]ie*&��P�S�GȺ��;�t�k�����̛7�x���Z��tU,P�HN��΅($���rf�ßj`k�Y��D�y���;)$�v|�U0v�6b���T�W=���i���]>�l8��dzo?�p6j�u�1����6"������)�ִx�IC�������K�aʎ|U��^x0|l�����׷��`���h=iB�*�q��\�Q{��ؗ���g���.�'���w6����  WX>/���-�8��Xi!x��պ�ϑ2=��ٖr��<��~��6g�N�J���C���эvqu+a��b#"���\"r���#�Z�#=�t�@g!�m�9i->��uo�G`�Q�����~�uY���&���E�+F~ Z���G�G�.}b�;Y�ˤ���33�S��"�L'�O�m��t��xPE�ý�w��T�'���G�ơ�!���o
�&<ل�t�E�zyQ�������xa��s��}�+n��k�r�?�c��l�/Wb����A�U��� ���_@M[LLV��þ��^T�D�(������]>ڪU�6��V`]��%�M�wd�׻�����'  1�y�>�AE�u�e~φjʟZ�X'�P[���b�_Ʉ&���ɎX6jV��5�6l�e���$37d�����}��-q�\�K��v��R��o9j>Me�NM��@�ɢ�d?7��Ȕ��f:�oIT^�4�?j��|�
�r��(�v���t~Ӵpkߏk\G�����/oDտ�f�ljS
:�q}�߼�v�$X�
�������k�hfF��+�Ù�6���ٷs�'<�$�����IAUfw-~�r ��,�&zX�����F���ˠ4>rC�K�[�;϶ML�-8R� Fm�!�Z��a鞸��0��7i!�q��P!���Ѻ<��+�k8���$�	�ɬdj�$���M�����?C�]�a K�W�i�Yғ>g҉5����HRd�]���c�6kl�{}��ݡ1��g�|�|�Ms����,��C0m�?�$�~qj�ㅱ��q������C�� �8jl��A�c�`�����'��6k���ƃ��>zI�iyBձ��)7o>�:t|�� /�g7����gS<C���MO	�	�G�����f��}����2;�2F�a�K�K���c~N�< -�ªy*4��M ����}��RK��2�
.����t���I��^�8g�S4az5�Jܚ�����dY�l��bԜ�M&r���L�BQFW�:��CW���(�mt#�M?tN�H��R�%�w8��7V�/iU��|{�`Q��h���ِ�ڔ�\��8�h�$
\
�bx5p'BL���D��/2v�o��b~�� ��fFrY!���<0���h�7±*��l�at�9��H�XƿgݩIDH�xH;Z=��/�\�>��Q���Y�mng�TR՗x��.��s�'ma����/Nqә^�M(1 ���뒒H�M�k?� E�,�}S�miғ��F�plI�◃�%8����W|��80��o�|]C�J����<�y���j�s^+�M*����/ ���x�^1��+�Fs��s�l�ċ����w
� Ր�vČ�(�]2w�Ӵ�>�/#R�_�r�^�����6xU��<�.���-բɇ3m;�0v.�?'T��8u�<꿂pY��E�A��БЈ.������J��ݓ,A�E^��e����	[U�x"@��f҄��n��*ބJ������?}�Գ'���aϽ벸��ƛV���>.����ַ����қlWr�u��ip�P��"�7s�i`������Y�����8)�n��%�ѦɑJۊ��S�*���Ka����A��̀Ox�yl��m���[���r�@��'؀��)>��h3�'ߛ��	�&��A���$S4а�O��3O>���jB��j*����ns�t��z;��� �I��sG�`j�������Ƅ��H6��ǫ�.\�� iR.s� o%$=1��U@
��
��d��K�py�7���Ѫ��W����^��˗_�'�~��N�F�����^z�����y��� #�� �T<_!��rm��B*֚����c�S�%�f�'}�l"�7c����$!I;�i3I8�(5Ѷ�_.����H��eA���je����XH���vʄs��������SIc�-w��@"�o�lk��3���s�}���P���L�H��/�6��F�։�h?O�J���.d��ѩ���o�E(���/��ŏt�|�5�L���?���[=�~qW!�!�����6o��K�y�Pأ��
[�3� ��X`�
�0u��^��M�>�E"�;��<�7��(%��і*w�"Nd�ͅ���r�G�%�n~Й�O株O.���a"�i*�8sE�;��Fj�/�^�Za$t�����{����-?�|,���57V��G�)}��P��.7�`G�M(c3�}��3�ڠ���h˕�	����s�����W N�er�*R��i=���0�Bf��?]ځ�_��vǎ�ǚ����<�mE/�8��`f�	�`\�t��\
�����M{2X`܍��d���԰LU���&.\�~�ʡ���8ՠL���_�G�b��MM��}p[5������I}Ɇ�^e��)hE@3�7C�)fIy�� �S�E�8Џ}J%����9vn@��;�"�:]���ކf��gѡ�#�|��SX�'�b���a �DΓ�#�����2 ��r 4r�g��=�	�I�x�����F;xy�E
���P��ɰeZ۞��B=��~Kh�P�=�_̌�MV&]L�h�Tn������1�I�
�rgB�V8���bKo<�]}2�p�_�1"�!7�ӲMm�%B�thȐ	��>�=YM�KƋ}@�P&���5�����2�=߉�J��$!)J�4@��z��Wam rhZD@oǜ?	f̢D���݋a�{�X4V�jX[F��O�V�Ftg YZ�O&�jgl��V!:�W���T���wd�-��s
Eϼ�ZL`��l|v6T+��Խ=~v�e�}S$�e��Qn�̙6F8�,�{������+��=`��v�c�H璓6FF��L5�,��,��ؔ/O~�ͦ�c�% �� �&s�@��H��S��Պ���i�mK��c�|��j�$J/��Wg������6-֘���V�UB�N���	�t#���l[�߫r�#�>5�W:J��4��G<Dk ��-^�O�6+V��c��:��,�]r�}g��|xͩ��f~��P>qXR�L�����Z(i�o�ҞG��1�P\�J磡��u��zO��k�m<�J���������y���=p+	>l�o*�.˲tW�o�2���zjcC�����|�6\�����,�����2kO�T!�b����S���E~:�;��`�����P2����¢��FI8���q�,�e�S&��%���:�/��x��]�tn�ٓ�� Y��$\���Փ��q�c�+Gh]������՛��2{�U�_+i�D����<yhwʁ��/o��l`��B?�a�����J:a��ώ�p�����	�ǟ�-cn������9��+4x���5��'Q�8uk��2��9+S��!&�^�LC;�6C<�KP ���,�9��7��Z�58����] r��	<Ky�*���_�T�}pY���a	pd=˨'��jU��>��r@_.&@�t�����{��K<ra�U�^��jڿ�j+�L�6�*�X	\C�h�i�C����^�\��^��Ӈ�V�W(2�ӰT���$:�ש�Of��.���2���[���b�',鶐���Pär@���ˮL�k7�tL�=��ѝ����"�s��RXw�G�B�o������:X���ݾ�t?j��S]�:P�Zۀ�]�>��0{"	�i�([��6$w�H�u�ı�Y&����C��rp^�L7��	��=lC"C���Nt���� "�*'*q�g��?o�	ˏ=��Lz��� �z�(����u��z�FN���Ӗ���#�!ض���\��R��촑y{�P&[�����k[�
�Wh�Pz�0N����brO4�MI,XG���z!�6zv�jfk0K�E| �j�N�R�G6k���ASi�7�"���y��6W��9�j�4����><���8d���@��V׺[�:�Sj4m���|a���
��7��%{�3t��w�,����>�R�����OS���Tp����GJ�҂N�y���R��5�s׹� ��]=w6�M˿N��h\�V�V�e8dEa�P�o�=	�Ӄ���׃���GXZk���K��fzY�P�9r�` �����禳�GΛ�-V~�S����Z���Q��a���%7��>k6����e~T���5�l�K�$P��B������O$/�:}8�z�����k1�r>Mr�*L��F`����3}�`+9p�ͺ����f��Ŏ��;���v���XQ��`͘2���V H�%�Դ�%)�B2�dE`lUa�;+ڇ�'��>� �u�>}�ze �I�!o�i�ARv k��"ԻXS9z��'�\�M�8��ћ\0�7F�4���M)��Xr=פT1�"��	Τ�-�-�XJp%{AB4<��ݍ�F���o���b��LR 8x�-T�=��cfo�lP���G����g��3"[`2nʢ]b�z.�J��\�NM�s�w?�v���z��q���R!����|����y�8~��Q�Q����?|���#z�%�<1���k�M�[e)�ˆV�{�(��Pի��I��H踊��q�P{��c�.@���Ã־�ޏ�����\��!�{E��G�aY�c�Uf�ϼ՜:~e�:q�	�����*�`Z�xg���n.�+���Hs��oTVZ�5j�S�h��I��2;�Ov]KK�1l�^>Ky_��;�qS�!��~0�����\.�J�*L����e�A�@*8���Fx�]8�o0bc���c2��\!~�nK<�~DJ,��P��4��剢[7�'h�PeԀ��%p�BMIӨfW��\��HA&q%d�1��J�>�l��?+�zT4��jj*9��B��1��=[�I�%��`&U/�F�=�3��v_w����1[��4�����2G��4��?Ǝ�5Gį�X't�'���?��x���cl��N"턂�G�@N��m.�a�9��|��hX�Ŧ�9�X�FN�ڋ��_T��
Mq�С�%w��SQ����g7�_!��Բ�����=�����GT�*�ۡ�Ӵe$pGSF�(��G�ba�6�DD��/��婤�������G\���^:Nٺ-��Y�@2����-��%J=�YqN-�J�q
��(�r�:殗���?�vE���T1����Q�}�0��3���Jx��Y6;�9��.�/O����	�ئE�)���}�~."qi�Aϟީ���qG,��i�>0��pq�V��t�ӱKL��a��	-�͏�.�Qn���P	L�>m�n����Ŋnp�w����ޜT������� ��y/��o2��˖w�ֆ%�F�o�d$4j�#��^C8(,��v��_x�M�P�y�G�D�_�V��	��s@��)���J�>�.\���D���gw��ȃ*c�R��|Tu�N�KE�v�=x�c���4�!#�U�A�:����`�#��  訇P Z�iP{��$J���S);(ڳ�Fm3�?�������6����	����ZL*n����O��T�}l}'���e��lG�v�!+�h�\���].����+Y�����9�2�
[NI�XVP�L^��-�����Eш�J�7���;]�<�q�>6�l�w�r)yi7z�\9i_��87�J4�����/<^��fP��%l)ņ�������ȍ;�񎅱���-���*���p����$7���^���+}4e�X�Z�\��A2�Q��@��u��@��$?�N�T	�&�,NX���;�֒{O���>��������ٖ@ɫf3��LV�צ2�[�RL;��i��c��J�`�����3��q�B���Q��i�?���L+�C����<����k�"�Q�)g���ʆ^�^��m?�Ta�,�'�F�=�����ћ`�RV�t�ڵ�M��K�ځr��{���}��#�(<rjN�6@�GC��zst�(h��ݝa�e��D��2�$��JG��;�� %?j�����ɘ�'���M-�t�-����0)�p鱌�,>���1���vA<�6u)bl2f��J�O�R�ځϨ�Te�W�s�Os#��E�UTm ���+��]�&e�����8Vu�B�c��E��;!d/���m���q��6p���Mc6��4��%ZP��{��b*[��fk�u��q�3eG=�=���'�WNp�������J�Lc-�>�'���T�Ͽ�C���O�A��t=[���vU9xPɯY�QM�z�=���G �����n!�K'�e���(Y'C_����x�P��M���?0�E���!���آPŮh�/l7���8��j�i����X<e�?缟I�L�4#���QK(�eYS��Ec�������eT��;	�DamQ��	�SM��gi^^]y|#�����3{t�2�"G?2�Oe�G܁���4�z�5oV�:���!,ȭ�Z"0��D.cn-��ʟM� �Fg`��Xg<A_�k-�ChF�����kZ!k���s�qc&@��H5�h�6Ĝ3��/����a�B��{�7W��z�|P�bX���L�.��}*��]��%��/D�)u2V|PۃI]��9ᰄ��5Σ���?��v`9�uC���c?֠
:��c����:a���m�3����&a�ګ]�j�h;�W9�Gv��Z�+W��	�����a�vԷS������0�1�F W�"��,q2��(J�v�*���es&�Ͳ��P�J�1���}��2��s��+<Q�X}���;�u�q?K��=�I���{9�c�� �����v2�ȝ�B)	>��ܪ�4N�/p|U�>��6�j�:�}3�����;�N��X�ח�}��f�A���сg#z:�I�oГ�6���@���@?����4�fF�;gK����� B��e�Pr���׌U���їt/�E9\�i%���#�lFE�����]�-"�5��#7����	�qe�N�S{�ک�4�:�AW�XEGI��C�P#o�Q��^���T�j��BZ��3'�^���j��>1�ќF��\ڟX�e��-p��iQ'c��W����g�&��Ѧ��!ُF���?���H�EA�g����}��0���T����p���Z`�R����^N���K:Z��T1�XN<NeM�,���~��q>*�e��Md{�Jk�sD�~kK����N�gp&f���#����u����.+v.��M9u ����aշQ=5�i��I��f?�t�8ӖM�T្�ޞ�ew�x�޸5ؓ�K��|��l���Z�,l�G����Y#}�AXϡx�	!��I��?\���L���z�M��}���ܓ^���XZ<޸OVX���͐9�`i��^k��'qr6����!�&��1��fz���o)Q��C��eJ�]1Y��
�F�1��yoU��x��K;����Χ&-�po�5���fł�ۖQ��K��F�<��t�
�6K�Ut7
{7f�@E��	�+�.��2��P�{��sS��3+:��:mX@Ӄ�����=�[�mS���t�j���D�����M�v�X-���a�͵�לB5���V�#�{ڮc%�*�!\O�(
���j�'þC f����bJ!�>�����Lǽ�U:�XA�^����;�!����/V��&ث?�ne1��W^:y5!�����\8YBߤ^K$c�� a�mt#��mF����Z��Ex����*��$٥���|��>�Z�� �F�l�>U�赩S����|%x���ћ{�f�g���d�_�n5S�W�ہyi�Q�25��\�1�{pI����?�0����}���9׶�)Z}�z�(�K��+ �uc��T���ф2���l+x
A�c� /y�_rd�5:��Z)3�d�Q���BI2Pjm��e��O!=�H'�6.�N@'x��D�M��N�����	8���EN�R�đN��K���Ή�5�CK����J��ͬO
<��Ln���Z/�?&�^3>xs�1y���צ�QbB/h�_���$����!֐��>c��B"���D��է={q��ll��BYT�U��Pҹn��� �r��i��}[��>`2>j齀������C[�݌�6d���ZC��!�(����
������ա��s���l6��&����Gmx�����?j�f���$����M�ӱ�*/���<Wr�4��(~��0���mN�h9���f�6��	��vd��Al�A�Y��9���
]��c�RK{E-F6�#��?�T��||�9(�iG�삟���!}�7D�6�K{��VG�?��J�����F �p�������
�7��DTm��}���t{z�-����y��?��U%a|�c�60��O�CD���/���h�L��_p�%a�ۮ��J�Nm�X��-���M}�b�_!�q��"I�UC�e�^��hޡ��2�FG:2������r���w²�-������R�fti�l���	�5@Z�����XU���:�O���t}�B�B���d�̕�J��.��m�"	�IH31����p�����e<���[�a�bϱ�B�3� ,��c��;�[9'U���*d��T���E��6s�8c.�glSS��C�Z�����o���<��X���z�I��[���v��聹����ܕB8#=�A�,Q����P�2�tDv�A�>w:�S[R��أ�`~ܔ^H9��GK��b}8��!�=�veV<{�����6&0��"�3��u�`1���"�u�ʵQa���iX���t�Q)[=����*G;�kr�DL8"��3�I!��و�G�������ף�6��P`�D�Ŋ#��c����x��#95�E�vK�Ƒ���m�ܨ�=��P��7��h��goB�ֿ�Ao�� 3��+�.�/�6��^�7��l�hH�2.���缦�����<����sꌫZ�sI2)��t�^jQ1餇]΅��쩇���C{� N�:/���ǝt�H8�~��b�K�f����o�rM#M�}�xH�<j�n`�(.�iGZ�0��H��-x�2c�������2� �f���0&28!M���D2Q�����4��IW/,�ZMA�#�51�ΐ�����j��u���nĎ���qE͉|�Y��D�"�!�Ǩ����~z|Z�o���6{����o��S����gS�mn�VپS&���[;
�˛��Z�[��r7�S�(�0$2��ց����d�L�(���OIK�m��>��ȩ�+J��t�R}z1H�G<���{���Q�f���)S���@!=|�W�]y�۳��:�fb"�v�	.��;�y��<q���Cxg����_0�
�2��R���{�S��(>��3���\\��H����)l��
s�kM|)`$���J?�U
Z.�Q��ɂ����[�as*�H .FA]@@J�M���R~泬�ᡘ�5Έ\sY�p{:���W��C��e�<�;��m��(q�!��6ܓ�j#���'�x��!Hp���v��֚��:�j�ث���ppٯ������B�E(]8��=�K����\嬌C�<a��&"��5���N�f���za�j3֏��o���]��%�KϹ��D����ch�r�3�j*�=_��#��h����g���K���	�&�'���L���l��
����u�+�q�S���|ϓP�=p��}Hw�j�-nxr��鬧����P"�HfW��Q,��(�ކq�A4k��C���3�L��3��#dƦff��R<(E�:�R�%�Y�
ܝ�ߜnB�F�y�l��۽��
�8���4�n���]=l��0̨��{��y�]��;r�}�;x!�f�9A.�@鄅?Zi��P��.�ב�c�g�ii9��J��:�%i��XA�$Ӗ6Q�uUJf|�)>�.���AO'8��#6(���t&F�$ϪB�`D����h�7��N�l��m�^(�y�8h�S�HN��ݶ���\9��I����x��m��ɏ�;�a�aH�
��pYJ��f���������7�6zQ
�e�4���Ba�0��%�-��C��{$|:�Vz/������3�k{�k���"��\���4��U�����ȭ~�{����>#��քl���])Ta�n=���#��͜���'�X�z�Ct>ѝ�����\�2!�XhU���܉�Ik�Q���u�I�f:%����n8�R�u+o]^jJ���3GO�a�g�ӔG\���+�)-]��ӷ�ҍ�`� \�ZwHL�k� ����T\hݢ��wY)rcE�
'�i�&�V�L�ǅ���^��f��B�C��aU�*>�=��Zp+4j~�:�`LIި��k�gZ���= {q�D{n�������Ѽ(? �ow!�Z>�z_w�v���4���X��ڧc5��`j׳/U{��L�*����K�a�St�i��a=f��L�iW]y
�3�@�^`��;4�[���#v�l38�-���L�^����$���v��w��PϞ����CK�exg
Lq
��� ���7�y�2��fػ����{�-�c!�Y��T���Ϭ�s�l�8[�:�L~h����*�S����a[������3�R.�Ɔ�U�"�ܓBw����'�y	�6]@oܞl�QI>�Y�fFR5��mjY"��5ڲ�`O�Kvdd{0�?���d�hQ��S��Q���)ߩd��Q[͹���|����F�d�����b�2hu�7Ίq	��s�d=i�+� �EzoDX�+A��}�F�S�r�� ��P�B�	��1����:�� Sxk��e<"��4o��xYO/��c+Y��;|,w�f�g��<:Es��1�tF��(R��]QX�t�r�M�qȖ-tPǠ��	VyL����[���bEl����z��u8�ז
��	�g[�/B&1�:�-ވ+1�!��	�Owؼ���L��Yi��.�M���e���!�	sҔ���8� u�C��d��v'7��>����^q���`���$�z�x�0���a�98�ȏ$�6p:߰k�kf[��qL�Ϧl]�)38��X�-~o�IG黇HؒL�w��q��v^?��̍����"����*2(����������:�f+��
A�3��^A��Qz���o%Q���7p�h��ϕ^Oy�şؕl�5$U�]g#`F$�r�d��8��B�Ԉ|N|�z,	��h�����[���R1����`:_�-<IsEɶ{F��N�s�g A�1?98(���xy��ʑ�T�S�ow6��t�X��dbt����#���"c���1	��|R��o���2+�8��^N��3*�CE���L@��cn��Ͼ���y�J��
v��u�o��C����nx�Y�G8�G/�����'dy^o���/2Tw�䭔���\���o�{d?��W���F'�p�#���,S��tr' h�.-D�/���ep̽�<�5�����\�b'�,3�:Z_F�m�=\�5�1��X���o-�w:����K�jy�A�/[ƴ����h3eM�Rz�ֹ�3��R�l�����z(�,&�4um�q��8D��9�Z��7`���]�9�	:��j�U_��0�y;��،`����1&�@[Y�3[��,��g"O_ 2lkhz!u4>c2�'�Q+��V��U�*"�}�B2K;RI5�H����n�p��b�(��~*�/�����B쩞�$t�S����H�Bz[�~���4��gE h]h�4O&��l��̹`��18u�V�͋��Z�5�q����~�w���ヅ
d��|�֭���@��:��W^ݢth�0��
����5�Ee��,޺8�j$��	�|��G�_dp��_�˕_��d�S޻"��Un^���q�w/��0:�Fv}+=]v����˘;�k@wn[�vmGB�-��P7�T�Ky��7Ob5�� p}�i�.�.!~Ti� ����V��Jr�PN
�O�xi)�l�VM=���f��mG��i��鵑T(�/�y��j(/�C�\��������i�je-�[7�����ڊcS5X��c�N�:�\~�**�sځ��	6��"=/�RO���Eϒ�G�ƚ�Ou��2��]�mXm]��V��_���k{��O�-�г|�<o�\�b)�q��6�G�d�	T�睯�Wvɻ?�|���/��9�iM]��$n3P��ˌ����S�%�gdeF*+u>��`�a�����AZD�<���E��P3C�?�����lO6<�-.��c���uX,�8s=x�͛����B%�S<����r�Wlɷ����#�T�k��ўo
�ݶX�B�@�#�w��V�6X�{s��GS��؏4�P�F���\�zgMЮ��p����P,3\z��^,Ŵ�z[���XAA���U�He�a������]�`7�5��Ȏ6%�I�$���Aq�k[R�b�ݬ3*���Ì�q2��Ǹ��^�JAP?6�1�嫓e:sb��OVכ�0޷Ipk��:꼍Y�&&�o[���A�!�a������ra؟����i��΋*ˍ��J'@��J������#��;)u\B�pyu|�8E�I�������u��ւ&V͆���g�[�%N����@ᆔn��$2�LQ�A6���,�Hq����o:8�ظ�Gԑqvސ��`�'m��|4q�|����L�د�c[���f���#��^�TX�K�ai��B�?e�ķ́�4��w�r�.~�c�����`�p�K�6B��)���T����vs{����{��A��/�:�3$ȵ�#��*� d�� V6`�]�	Pc�)���n�(�"
����R{�;�G�� Z������jB���_������p,��+�dY�Ha�����`�F��v��N�';^h7�f�j���Ϲ�3ܨ��_Ѓ����6�b!�$��pJ�A*�Iˉ#������� �LBG �K�=���?h�W�.<�z������׵#�8"�2/@���5�v�\�J�Ԟ�帙�k�l�5�3A��E�Kmr�Cآs������#�	�=��cb.[������x��ȭ�H�<���4F�8��
�&/̥�����>���:�;X|��>���(���yC���Z��lmJZ��惼8�j�p�xm/���i�6�*wE#��zeA�9�2b1~;�^6=��i���6[����HD?�����'��j̲�(��w�|<�5���h�?��,�۞}�%�Z�1�2E�_��w	1Z�xm����~s�Ύ,`�ҟT�Բ�w�@�)�����ю�>�J\��d4Ɗ	��,����"����P�L2)�u��#�N�>���31m����"�s�����Ds�s�J��K���7���hR�v��ҧ�Yt���0��Tm���P�H�jk�gB��K����B�ˑ��ݳ�Qߵ ��@d`*L@6^&��y����~�˹����(y`����?+L��_)�d��W<��������$�E��/hW����[qN����W��Br��*�e!P���#�^[�T�!ǴE�u�Y��~֏�~�#'xn�2�����hl�;3x�%����P#��T�u�'Ol�2X�G@:X2��;y��e�.O7UhX�6��d2\"�ǲݼ쑽�� Hגy��n�<_��М*�@>�2ZK
�0R��(ݴq=�U����:�lW)�{U����-�$�m/'��7�v�ib�;�Ȏ�?r�z#�y�EݖYt�Ɵ�����C�-�<;�q�Xb���0cOC�o����_i�˫?�.�]|�
�3(��V�5���3�`7H�mȦ8;t,�:�<E��Q���L#���Mnz�
����{����6���'�� �".������r����^���2<�zqJ3 �%�"���@�����m��u�����8�P6	@���@�-��	��2ڌN������J���B�'h��w�ӛ҂Ch:#���x]����E���59՘�����{�-���Zs�=���&���o��H�=�#��:���k��q?ܝ���/6��%���B��244MӯU�Q!�2�4`Ѣ:D��p���
O�A�u��$�`سo�^�T�a�{E��e�չ������7YDj1p�2Q�Yx.��H�'�'W�����t6�6a�6��v�z����>�:g�&��UX��p$A�Y4���J�>� �K���/&�H���#�*�P�Kº�(=I�6*��;����QPQ
��ǃ-���Wm������{W�O�}8s������7��-�&nI��: jC�ol)�ɛ1�Ӫj��W�Ȼ�ma��̽$��7q�5�1�z 8?-�X�ȡ����I#'Ee�ڟ�߯q�ц%�����o�P���p��H�*�\b/�0D�����`{�6/�M�Z}U�m{��wS����,��2��	
�'�B3|mO��EJf�"��Uߢ�U&���*�8�\
�f�d�&��ˡ'�ˑ��K��f.7��O �e��ȶ_�1�q�?̍SEt��HL�\�����;���H�b%U4 ��&��[P��������g$ (�á�6ܽ}v�����L�� �o-�6����u��2,>�u,�u���5��F���\�^�+�M�����:������,��Ӥݤ�<1�e����U~����mkW���W��{:|��M���,Ϭ��qԭ�u%��s9�i��e���(A����!Z�2�uQ\I��[�ZXѾ�6y�^��8�%I�a�эN�����y�΃��\����.�teB���2m6ȗl��tI7�%�N�5�P��P�Q�s�@�v��;.��b�cܣ��M "?>f���h�w_�D��?T���X��O�a�}��*��6+8�V�X]��EW��Gw&��Iۍ���s�m�n�*`�߱�,^v�w���Ҳ��ڤ4�2V�A��+/�D<��ӌ�1�2����}H�^V(�&2�Op����.�[�y�h�hq1G�0�)<:T��F�t��*$�I�^��ч"�|��[֣�Y+Q��VӔ�?���R��2��,L�rlq��.��
�҄g'��R9
V�j��su��	-��a��؟�3lP�p���A����:ψ�[m2.E�?��8�.R򡩛�e��~g=�wa9RcF����������][y%t��`�M���_���H�N����b?�=���t��(;2��UЄ�w��z�#��y~x `@|��� [;ϸ��ӝ_�u�6����&��`$v%�x�/��)�D�Ts�΂�Ĵ��T����;}`@S뮶`��O�&
B<������,����2C�f1<k�O�ˏ�ً�É����+��"UV��q�=��"���a����r�eI^i8z)d�Y�*
������#�,��]���Nf��3�)�h�..x��M;Z&ql��6���G���2�sռ+.SH�V�浀���0n$7���7����n�0�9�ҁ�Y���b)� ��j� �|.RX��hA�v(���1����g�+���B�+V2"ڑ��ZJ��Q�&���n`����n�=�y���)�/���\�Y�Ӵ-��ȟ�ю(a���-/�=�9�g�/Aq��_V�!=�	��A� ��Qt�j���}56 k�,'p�9��L��@TFd~�k���1�hQ/�a��,����c�&�a�qh|��1�*z�_��C����b�+)�)�Np��H��8��g^ٲqC7A��
ե��+�VyʮF� i������`g5�y�1�6��<�֓�A2ٱ�`&��YF$Գ�@����峊�ߡ�Ѩ�Z��+W�s���6�GZ�ܐ�&�=¬�l!]�ꖾ[b#3�}�7�s��	]�ril��fQr{�N
�����ݘ�(f`�v�=j)�����,���Z�Ʋ�#��)�?M�J��(��W<��v���J��2��%��4��P���1кW�?_������%�A�n�-Jk�BK�j��N�����І�Z��0�Թ�����m�I��^�9r�_��~��O�y�	;�d̠m>>i8Ez��T��iS���Ѳ���ufs����pA���� ƈB�
O8$A�X\��N�&���1^��j�7(�J�2+rRW.1Q���j�n�feHm:p6�tAP>��i�<،�K���W吭���U�|qx{�� z������W�s�Ek!����Ob��	S��e��R���EH������/A ����K�+y*y�_��- ��m�j�>�G9mv���u,�F��!R��G��zMً֢�`n���K�Bv�eL�5ɣ��Z%4���WI���r�x�b&|��6�9�����!�X��
�i.j��P���|���W���i�WUe��<��L@G�g�t�}�WB`͹1B �!��jEc
�WAuR�q�cg���9�&�Ry�Ι�Oe����7h� E���t��:������������:�
��Ş�~i��fgA��#b�:S�e��]����]���F�2@	��~�v���5$0|i��O�z��WG��ՑH�6��x���֐�+j�s���w�1��N���|ۦ_55���xܴx��
�h��4��&Տ�rKAgK`m����aO��M"�,��Q�H.Ɂ}��J#/�f��;(���u��v�x���4�t����-)�5��q��#��@k䵡g��������qS���61Q�D������4�W����HS���@u>��n&���w�q<���$�*?U����])��?e��֢]ǭ���+�W�ݜ���gO��� x*�c �d��`�`
{�d��
�`Gp|�H�V��>!�-@0�lcZ�mw]D�T�����-���Y.Ⱦ�[�u���x�������}\�<��"z\�ѹJacٵ�i�Q10N���a����\��9!G�����0י��=�S&D�Tr�4yV��S5Q�Lr^-'�l�UVEPБ���>�~1�U͋�#[�'��9�H��ɫcS�E5$����$?V�s��6��Rq� �/��(E�u0��"\�~�:��h���w�B~���R��ֽ)m�s������M�׀�>��na8�)֡J�m��<�#���s�6R"G�,<���Q��t�����-6��jw�Lei������Y$ׄ0d�f*��*�+fV��{�_����=�[X���NH}s!�|�m�\m*>"}��ζ^��3��ߒ�5�u�]��O� Uq��T�������B���$rz��d4¤ٕ����x�Z�R�<竡=Mn��	:��l�
:0�i0�bhefxy�9�'�<��Bq�#� s�����s�Esk���^�Ķ��PQ\���q��,k�r	%�(t;]�˯�����a��N���@vb ���U�>n
�#]>A��"��)h��A��t��k���\�Y�h�3��  }#���G�`��#�gP9�ƮQ!_�f ����`w�7�b��J�(>�Yy�s핽u#$}\4��ri�t���Q�P,j�B'��f�'���0��F�mU�W���2}��\��ъ#t�fm
�ŏ����
�]��Ls�'�.G<��8j�A����F�1��I�jv^�������u�a�Wd�g�h�Q��p��F;�j��Ո�Y�n`d�Ƅ�#_S5�/+�X�,ϸGђ���Kh�QI�]�T=� L��f���g�(��$�����V�U3:��Z�F���� cE)�ks�o�n".�w��}�ۻ��w���[���Ӵ%����r��W�~S�mQES^G5v��xz��/Xkt=�}N�[����.q���n����W/��Č�K�й�Y�ܾ��bYI�k�e���Ad�_�u�>A�8+��λj��aF����QքJ���TpP�\��{h�m��y�q�J�=ؒ�o�i�})�zx� ��C_v��{�ja�$U�?�kq��Ao��JE"� ���-�+�=I+������6=��Nt��S�:�!����R�@ ���ṫX����Kj�	�i��K�1�[��e�huAI��%ӗe��dQ��|A�((�3��tu�Ǥlh��8v��U_�GrH��N'-Y�H ����U6K�+���`r��f��	��/�	��o��\r�%1�6�cT���\J�z�5��P0%�� �~v�c�0n|+�o���w ?Z�P�v���vg��s��qxf��Ľ!����ٗ�Y����X���Y��.���m��4d�nfz�qL$г��΁QQ���`&����'O��:%����@���]2��:5ͳBdQ`���R�8���:���@��>��l��0�5eeFq��m���g��}�Қ42"w_��dwga��e-���_l0�خ��Y{L 'oP���&�/�l��$sz!����0��"I`��TN�����e��R۳��5��GƼld�S����'�R�2ڍ�]�,�P��m�;c�=2�ӽ,xҺt<��nlZ
au��
ͲtA�����|����B��D�	Si5�	����f���vG�X�/�gڨ3{��.j���B���j�?+i��.��_ۙA2�n�1��j��\΄GY^�X��b�m�M��@(�[M\����k�����$�k{�e��$:��ɼ[��$��b5��[��y��w�:�I�� �8�\�R�p����^E����E����~�J>)�"��p���s�u��@��Z����}x��*�,�&|�x�� >㈻�Ipi��_��F8B�<���MA	�5(�eA�f�D��>q�GN�C)��Ȥ�;�=����*�\�Zv���e��'à��Y
��0�ki?M��GO���$�pԒ�ҳu��~k�k�C)6X)MS�Ā �����#�U�R�#ߪz�����~����%�����p�מ��b�>Y����>���C�J̙���C�`Y�XʘV~
�9ߙ��҄�zPj7h��d�t�l�EeR�Z�-{�����a°�µ{+�F���	xG=�����-q�0|[��x�61�3���:,��
>�+{�2�_�.r�T�Ȯ���"t�u����*-@  (oH�h��R��WŪ���������7�l^�)�o KL��o+� 2(���!�`;E�<�����6�:�T��`�T�U���^}3��m2@G:)M` ��'v.2
�Y�؀ra��u��NRN/���ץl���1�!��,��+��xꕊ����SשQ��Ӛ&~�vO���0��bHHO�Φ����?N���~��ۍJ�[�J�dv�pI�~��,��E�Ԯ�����e��V��OH=+!���w%�ԝl6k�����T�a��Ϸ���)�bQq`��7�V��1���[��[J�l/v7��cO��.,K6������(����;�s�NCG|�}*��K��1��? j��'0��Է���lz%{h�`,rs~�)z<�7ek"�a����Ͻ�fh�F�^�-U(T�
�)����|�ێM�]	�����أO�D��%��!�ҳ���ןq)�v:�?��	��(������+x�rc��Z�~X�l�O6zJr�K(A�)�2������6~�E�2i�D<J�����Gef{��h�(��O�ʢ��/��ل��pi8��O�@�~�˟�%�x��N��;�u�	PϦ�77��ߝ��A��Z�� }'�&B*K���6���0�cj@*�gC�5 ���33���k�.�LZ��d+)�z闁�P�У��H%���L���CBV��u��mU��?ɭ���Y�!��#�~M�`��<�X*f�A�v��D�}���D�9kh-����[i[��G�[i=VC�d��t�����|d�㲇���;Y����O�O"1�L-ۋ�_a TGYa�8�*�2,#����;��c�"n�m��r�1Ѹ����㥪6���I#ȟ�<�|{�1���+���|Q4�j�)����4+8ekGtA>��cKE�0�n�
���ՎM8����-t����� NR��W��i�o�&�6=��X��	O��y�'���^-^TI��f�Y���Zh-.�A����S�~��8�2nM;�v�mS�f4��3���kF�}�jD0�~�.#�FZ��vC`v&.����x�R���ߚt��/ ��x�ٔ;O�xB���V�6�#�AgkL�&^�Wz�a]�)�u�q==�E<	ӯ7�m8��VR˝Rx6_V���u�IY3���#��ҟ�QN��&H��g1P�mRu����p����~������ .����s�R��5D坵�_�@��̍
t�ěhL��Q�C|�E���>%��_��F�}�������k���/o�(D/�����1��!����g	,�8�@��WPճ����7��W̤����>���I�����9�_��:V�p�5�=��A���VLy-� E*���հ�ln��p��CF����D�?��V��eZ��#��~���vrI�^4D�M��t�X �����d�݊���MB_���F�(l��E�0�>�ɬߝ���ʫ2��2\���w�"T��_1~/}V��|�R��5��&.2U�~�\�k��tD�[�W�=~���Eۖ���|C�OQ#Y�W�}��]��������B2��Ĵ��Y2}����Q�%i�Z���!)�DliUǸ�&{� ���`r@OZy}Ѳ�z�,���X�y}�/���$%�Q�q�8jZ�2j.�E�ؼ)�Om�*�?+v)��a2�H�^� Lݴ���`�.!����U���|�0��ޟu5���zj���i����7� ��F���"�p� E�"�w
�A��M� ��Ѐ�5L\��s��\4bZ�eګD����9,J�������7���I��U�#���k����2�9�pz�)!��A9����Z�[2����W̢�4��Ra�O�/# �)�в��Ǹ�H46��.�S:��Vա�՗�:Z�YѢ�+�'B�ͯ��_y�h�W�og���덣��j�.o�N^{�b�z�U9�~�v�Y4���*��7?�ι�M��9aT�7˩tK��)>��0 s�!�1��J�[H�;�e�ϭ#�6�0 ��l�k2@ч�{�ZJ�c��cY�� H-��Ρ��4�b����TNl�C�R�A��k��3u�r��|�)�����K�l��l��E��߆��c�櫒?g��=G�~m��IƇ������~�M���;J���_�v�x[B�x�F�ģ3�{Ԣ-�S��nXސ�1����a�''�Uf2�)\Y�z0ɠ�%th�br-`�����]&B8�FAC�.��wlOI/A.\�
閶�O���;��n����a�/�R	ܹ�� 8�)��Z'�{;	�<��g	���Ȟ�x\h74��:F�q���Y�"��1"dF:�
��L#L|z?���%P͍��O�X|?�b��FuH���M����m|���װ@?M1�7Wr��|��� �P+�.U,V�
�)/a�!6� �~"u!����wM8�����S�0���������N�-��>�ԑ$(ܑ����ML�=;�~"5�	o\P5(������a���J����\�s����&ъ5���ZJ�ߩ�� t2O���d�������vOξ��%�7ũ�^�z�KH�@^I���@E��6���⫕/%<�d�̸���&��i��� �q�����9�DlO��r�b��+P�j��q&.���B|1�ڜm�)�]ʷ�D0����G�$^Rʨe��D��MN�%�*�W�udI@,Oq|�M�����Hdb��&C�rB/�@\�	�|Ogv��Vy꧖h.�B?�*5���B+�W(��gUy��R�.U��v���J�Y��)�`#Y�vL�����tZ-������=5�״��a�|�8�;�y=oV�ğ�۾0�̮j��C�6p5�VcˀFL����
��˓�(�~�x�Ne&�GPmT"��WS�lu��+�ˤ�G�FR=p��9\sN4��q��/ɍ�T��%?Y�9����5��2j%T��N^�fi�@ʬK>�Z��Q������twQ�1�;_W>����nā�H�K�iJ;H���z �g,��������{��q�Q��	A�����a���N�6z0�� �PE��_m� �z� �+~�g�Ȃ���KSK�M��{��IBF;�zv�m](�ḥ����HD�z��۶�b��8��� �����u�hBx��[�2i���Օ滀��A�G��r1q��=w��Z{��H��@���,�dm)ˬ��40u�-�Jy�\k�z@ !�+Vu�5�Ė�Fi�uR���Q�=�;��}��5e����g�V��%�/ ����8�U���R7���׋�������+�ˉ_�w��ó3���#�ĵɖk(��Ah���OHI3_IY(!�E��Aj��%�º� �ybQ7ln�Jf��&��ߤ������g�Y6�|�o0ieǌ���E��4�놪8x��&��_�6b�#]��q�M�SQ��?T}���S�ĪdB���_Д>�0r$�94����n2�kR �SYT��6zЧ���"��hg�"�?e��q �TbH����U��B������`M���`�\����}�m�i3D65=��Qlk�a\\�Hr&�<��w���Na�^C�����B�"���یv�	����������>v�uf��.x��|Fo��������b��R?��;��g�;�3B)�&z<�}��E2.��9���}��Oa�����eV�2/�WԾH�o�� \ߗ�ݼ��f])�S�w ��tE���9A)^s}�<���$�O�����/���B��?��Nە�]����p�fϗ{�w0=UUI��2������P��ʿ�]B�VDb�H�r_���L��1��c��nF^��'��e�V�.����2$X�Cb�Q5�8
Su�Ɋ�j]wbv��,Kڀr=u�E�0k4�6ݨ�0UՂ�BZ���^Ю�xv�&���(�B��"�<���;�ޥ��Tc@�Ǜ_�~g����T"rh��T]�0�Ӑ���7P�� V�$z������L*=�#Hϯp\Ԑt9N�[�����N�u�X����>�%�9��	lEW��N��~�q���c��K�d�E�]��rUx���۝������Շ=�<��0�u�����R�f�Ɏn�*c��(n���'ᑍ�����W�$q��O��eɉ�6�=UB�X��_Y��rN��P\����� I4��-aZܭ5x++)�%�U���;��t�S��8Ʊ�3hi)�$%���}6I����)���~t��1;��J��cI�?)7�S���g�E2�.Q)=<F�O��B����,Oi��YS
J�	U��E���yTs��S]�.�0w����z��r���i���q,�_I���z�t�A��k�;ʌQ�(�M�0B7�C��&�YlK��&jlL��� Ht���8J
W��=�g]q�SxD�>{A?_2x?��Mq�3S�`�l8�]�a���$:M�[�Nn�N������i��[>vYR�{%���sG!�itk6����:����W?��QA�E��cuT�5��+�zXi��?��{��qw7�X��":6='D؆�x�{?��$��� L�h8�%�� S{Ua� j��H�ˋ�$�~>*�ճ'�]�~F��_���(0� \z�qvL���r+A�J��5�7�#n{��AȞ�Qѽ?�nHp�*}��x�w�xc����#���Q��xC�G;Njk��ܱ�m�x@�8��67�S6�HP�����.IpjzcL%��8�X�i��A�e�uHj��2�)��:I
qs�U���u�armo]���0n�gXv�f���6��\�s�V�"����,�}���?M.���l�����R�?�U3�(�
�Ƥ�Çp�����.�A�>��P6��ao2�B�Ğ����?IR���ۻ\�W�%��0]��A�Ǯ����ϴ�VfQf�6���M�v���p�v��-�y�5���		'E�wd��ȯH�U��c.���mh���w�V����ޯ����X3��#>���xa�~��1E�w��#�����L�۬�	L2�����f�e�M529A9@��-�c������I3Ct�%��ȄH��?K��\º�}R)[�"m�oM�?2F/�\B�_��vU�ҙS�7zɇ�2�fO��O�}	R_�u�W�B�XZ��1ۯg<�Q��:�3��E���v/q"�3M�qw<~�y�z�=�ݑ
.�>y�8�M�>��\z?{3�=M���=��^A�U��#5����	��jf(��#�?�RY�	��@6v3f\؟I>ɒ�K���S}&@L���Pԕ��[�[#sa���_�Ŧ�k��� �K4��~i�"�6j%G6E�M��ۣXP'n���B#OX�>3�R>p,���|�)��w�3�֯�qH�E�r%�zH3R�١�y��GH^Hj�����Lq��a��eܫ��;�Y�Ӌ�]L�v�NjQ���XA��c�t�@��@�7��Ա�8�����Y?���d�n�Ę1�Mԫl�ԧi sǜJ|�a�'�oy�P/�]>8�5����:-9��}PI�n� ����E����Ƌ�kq��M�j6Uʙ�.�_�g	��0�q��Q
��AإK���Z������̻'
�l�����@����da��ŭ �';��Zu��U@>^�Q��)�|��x��V�o>�I3�P<3l��ј����}"d�*.��ؿ!3�����A:[}w�̲ɇ)�ȟd$�i�BN@i��@[����r-�R�>*0b�}I!�`;���v<@����I4��GE(����ή�z0�����g��w�/����큀i3-��z�'k\6��r&jN��p��g�7�9���f�uF��Q�l>�$�-5�.ϩ.L�����a�Aux2�n�ˀ��R���PjW.s�L�6�B�`��?+�+�����.��劐Z���t`u����Ȟ���`�Q�<�p,ɷu���P�M���砬�rÃ��]�l��n�����z�,��I��E]B �S����f^F��YSz�Ck���95��>���9R[������!�}V@����(K��7����|i� ���SW2��NM�U��|��0�ѓ�X���(А�Y3�H���]��T1~���bU@�[ι�R���� ��6$��:7���n�g@���f�$�c�ce�c\r�6B������Ά��7D��Zyـ���o���t�3_�w�����}ψ'����r��w���R�b��~�tKݽ���{�y�b }���y���&�3�����ǖ���N ���i���6(�׸o��e�+5�����ۏ*.�d������Vg#b�u�6�L����2 �,k'��.I5S�4����'���G-�RC���s:�*Kď �7ȩ�B��Sg��%����ȭ}����J�\�W~':2�Iw!`[��'�b�^�7Z/.�5�=�>/�=�Y�s�_Ex݇XQo�j�3��%9�K�`뭿������Ll���+ޣJ�P>��������`-���+����&�l���{�hq��.:}IK_I4���1�n�K��5j���$����Ix���	�f�Qxq�	���J��7ϐ�A���B�z�	�}�)@.�.#����T�	�&�Lᐢz�Ч��|xY��۶�&#7�n�{YR�6x��ݖܐ��-���Dk�C�EJ�I���@��!Ha�<;�=�Q��D��&���H��~)�xN��AA"JB?���Ǟ<@�	Tj��[��T�����n�+����H=�G�Z�
��xZ�9+����w�;s�J`ީ� H�:�ֵ�%"
=�;���Ḃ��#�d�/QpA7���Y�<�����&m(�0/N���DGX����R/D ����<���¢s�"F��5��ᴫ"O+~s�C%��M@�-�=��y3�&81ڷ�����:���Yrd���J�����9c�i2VB��J����H�f{E��i��y�<����b��>H�텾�2��3Ǿ��b�=� C�-b��<������^��v���'��L*TeO��%1�#� �X����9�H�Ԃ������hS������Ǥ�0��;&����pdwu�o&|\��-r����߿�R�2�h�=b�ʛf���i��rw� �P��QBd
��.7��X����d���3�di�g"C��|�_�*��>CJ{U��ߞ/#qѧ�)쁭�Q�i�s���w��;���xQ��Y�L��*���(I�z�j��3��Jy}��«��pc�l�7�����Se��Da^�~^}��0��(�)�`�m=��<��`�(�#���zS�D��lAS&����OJ&?�d���色`�?�eO/�<����uX�	6�Fs引����"��S~�D�\����Bg�A�D2�w�ڇѠk^��(�&r��!z���w��̸���zQ��2����kfx�̗<�=Z+Ë
�t-�(}�f٩�`��Vf7���R�� �l^X��f���|t��E��c��NI$$zJ��{�W۸�I�z�<������	f�1[���:+n�h!+��ߑ$}i��G7�R-���n`C��|蕠s�X�Dgu28�ȟo���2�-�A.�Lbm��%9��9��GS�5�3�ԩ��v�U�F0�'�	k��Rʔ��Wg��6�t�� ����#���a��	��Jr��]<��$�>^W��5�<J�z�E� V��8�c��<��S�"R��'Qk�"�2ɿD�y�?#zX�( [�
G/���m9>b����`r\��}��ħ�[�#�,��3�� �ٛx��9R��V�1<,��{ID{i�4��T�R�QS�g�a�'����o/�;�iT婝�p@���z��1oZ�YN�h�y�9���n�<N�6���d]���7������¼��N�j2Ͽǵ��7^� 5�LS�6��)�b�v��ş��J3g�5��5_	��2J����u=�O�#�cc��+��j�a`�M�E�ؚ�ß,K�<,GY��������N����;.#^� !�5�3���Kx�����^]�BY+Y^�Y�UN��� 0IS*ze�3�x�I��[:m(<�*�ț��N'�Q� 3-ғ@��3��CJ�$�`l��e�$U�����O�o���cƯ�z\#���A�|�&�Q�/�X�>D��[���	�F�=e�(�I�О���2xa\���Q�u=C�B������� j�v��%P}Є��$j��-�0��'N��4"��s�P���O��e��~�jR%���IOnFHV�@	��nx� ,��lf�j��x�, ֑\3n�C�y�+���[b��찶�����QҖ񹭻��t�nlx���щf�_�,Ię��?��/D[[aUWH�w~��*�kU:kY9ax3��}
���^zO����H��O}�d��2���}jxe8p<�0$i����e��P/V��V�H�\��'��m����X�/X��f�2��֯WN��S��,�B��rHd\@M9K/ݭ��|S�Ž���D2��`��2��n	mѬ��jV�Ig�s[ӪcoWDE�*��t3�#!��EƆ��8�'�=}џ6(���$ᩂ� ��d'�W"ʫ�?�/�m�.6�I�-��ϳ����A�����u�u�M��)M�8dB�߀,�J�)"72k����	�"�US=N6�4/V��� �:�X<��hQ�R��t>Ç�:��=r' ƂP/�H���275��R$>"��{ᨫ�fR��f���Y�f�*�D�#��X\�O�;}<��n�'IK��}�����ӟ��d�iiZ���Ds��\$�>�k�2Cyw-Ҕm��;�t���w<t`5aY�Rܣ�P����|5b񏂰�v��k+;]x����}N��pn��f�k�O�(��qKȌN��b������ǡ~t2*ƶ��,�w�Py��bSf��9EGU����A��ξU�kۑθX�y�l���%GǊ�ε�E��:�ᰏ���f�|������Y�J�J'�.���[^E	na;l9�������Eu���	��FZ��DG�Ξf��I����lDl$��+�"����P�M�zN��\�C�s3�	ix����Li��'Ӳ6;)�T\�Ҁ�����I�f�w���D���i�u�[?�o�zY:�Ǎ��㦙�VH�d�Ԍ����݄2����\�}�4��96؈,��[m��I􁯽�����w�ȥT�)�!����T��,:�_)a��B��E�qf�L�?+I�4 �)d%w2�7�G4�����Od\ UK����%6M������9�����%)U��y��bjm=[���'�Ct�c�&�C�L<�n`�J��c!�<xmN3���H��_[��~틁Z�Kf-����X}�� �ސ<z���ʡ��?g���\��oJ��?R����57���j���[la�����> ��w�)|Q5���}�� ���#�O"SB"�{{-8���o�ׯg]�y���7�3)��)�����*��m��VYO����w����>CkEI���r�����ƅ���J�Q�$��aTȺ �Z`�]M#3c�.u?sqvl�/�G&+8!ԎD�^���h�+^��Z��d�on�<du��\貼gK����i��8�d�u� ��~��xLY��� ��LJ��Lj�T��=�E��T��Rl��K1ǵ<�����b��÷��N�U�k�:k6��q�,%�T mݽ��j�C?�����X������n��)>	:��(0�iU)�F4�!�1EHfȶ'�m❒Z8>G(E�/	}�l=��VSe802�����Y[�P�c����Βb}OK}&�Q���[����rE��NOz���eD�>�hG�=}0��.�
��ň�u�Q+K��' �(��@4L�	W.�}�6�̈́?=*O�� m��>��:��L�-�5"�����i����i��O<���oY�7�cׄH"U@��ʊ�u��e�a��-85j7#��bl��)��C��o�l� ,|��1��f��:f�܀�M���+i�}���%�RD��AΫ��-�����D�B�� �~����V^����*�o�i��Ps�K�|��a�J�:��BM���)��k�gm���'*�&8Y85��d�RK�z�Pc�\O��I@��ٵ�i:� �����2�K���S��_�	�#�T��(�r1��̾`X�Qj[��"]�ZUk�Ƅ<s��=�]�D'��v�5���Ĵb�ㄾ?�7�gK��4&!����s��6R��_�d��ь��n3E��I�w�M\]L�M����<� b!j�