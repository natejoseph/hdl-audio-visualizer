��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C��S3x�K���á�	��)���D����V�[#i.��G靿s���o�K̋`�wD�7��d�ធo��7���Jkr�����aM�,Aݮa���|$���Tk��Ci���k��m�
�X
�φ?ժ��������x�',����K!Uǫ㸝�,}b��a%�p���
Yr�D���9��]v����������R��B����pTmUr�o����K��66IR���
�����,��u�q��O�~��ӾA����Z��k\�xy��r3�Y��܁!xb՚lHKJ�f&��=��+�r[@u�����ey/Q����r$`����#B�u�g2(!�:	�E���A2�3��>���Al�ݺ�ݑP�z�i��.x��&��ط��v��f?c9��G
R-�j�q�:8X�~�����,0~G�zF��d�4%��N�����fĵ�\܃*�sδT�cl�uѧ���[f�0`y�؍�i0�:/��t�F� V��Y���6
��뢪 w�hi�v��a�͢y�T��J������H��{�2��s�/Dˍ�IU}����-S`�msBF����6��8i�u�����@�`�#��g��9�a�A���1�O�i��_���Ue3'T��rc��z�
 �=��GRW��Wyi��Q�zO����:4Y�k/����bw|���M�P�L$�tѷ��>s+2>�VYsoÖ���h�Q'��8�泐���5�	[г�2�/@�����k=�d�X�_��Oퟶ�Q����H�b79̤tڇ2/�JԎh.��m����v3
�4qл�ۉF5��ϛ�7�����/��-1%�ւ�hl�ˮ�t�-H�B�V�lx��Uo���sK?I hZ�ѧ�����F	�k��H2e�U�!��c�Oz0dG�U=�Y�;�k��qE��?fA*�ێS���u�J<&o�t��,�� �ս���������C����K���ԛ�w~�Q�����ė������u�����%��_����wŝ]����K�c�@ɤA����a39����kY��R��	U��"�a� ]v���rp�ǃ��S���5��Y���B-r�H��U�W�~��˃�,�/���2���:=�ʙX`�	P��7���������u,����^"   ��T͒�(�G��I���{s�}��#.��x�.LU�n���c�	a�Y��b�\֎1��0<k�E&.l�Ʈ;��