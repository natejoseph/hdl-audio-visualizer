��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N���ֈ���ß]$�R��������f�n�X�+kfm^�M'f�m#$\^VV��0[H;^t�������7�c�ge�3��"L��H�F����u����t�2'�l��bV��	���*�(^JE��WwŞz(.}I�ט�D[�'�vz_i펈*�+%gs�.K���UYS%tR
�}�K� -6>E�094�����y�=ޗg\�$Ed�6W�?�t�R��1/|O+��[d$M�8�ٳ���w���'��0�z�H����^����~�� s�vǎ�(�Afa�)L[v�@e�`��
�ʃ��e ����~�u�'����}7�e�$4�������v�A��aOB�]�W����fb����K�˭8iB, E:1��gn�����M�ue��ֱ
���SK�l�*X"Pg�g�&�������^���5 �b����kb�,]��ԇ�b�@�1Z^�0�ޝ��ґq���TS��O�\_n�f�ѹ�=�=Щy���S51u�/y?�Ł1~���T4���2K���-�Y���1�#Ҩ�l���ΐS-����������nR /����(����.�����ݕ�����sg�C]X&:�]P�	>�\ �8�ǖƜX�5O�4��z�R���-G?p(Qe�۽��fũ�@S�4���`׎�/A�1rC?^�j�Y!���A{�Jj2�[e�Y���;p�p^��v@ Ƣ(e�{0����ؼM�m�8�z���(����p[��v���E�Xƭ}!;M������?ݱ.wM��`��W�K�2s	��0:�[���kj-�͞y�������0�~�TW4;�-�r�w�����tւ�s4�s.Ė&��=�	k.�~�bª��̶k����H���ߕE��9�|���&gpȆ;�N������+��_�
�j�3�l�[Z���h�@��I����hMӯb�a��e}�%ݫ�J1j�6?��.�{j�D5c�O�l�*C&<i��drǤ�wu���I��$r֓o~6^Lji1�d�T�c��Oe�v'�u��Z���oB�aK�z�$Xpv����ѨP�X2�2ӈL]��$l��YC�s0lZ�`s�+n�<θ��$����/������W���������Y�,ђ���I���W���`��+;�.k��5��w4�Y��=��;� ��lD��+���G�l:?¹�W��� -�æ6�Z��XXG���`ti��\"ۏl�`O��M��r[Q��C6�@��t�"���R�~�����p:�@|�Y�yq�5�p�dLh�X�#���[ ������锛V���r�ҋN��%�˭��+)qR�d�?"�t�L \"�����d'9���ả�b�wtvg�X�!�aU~�(Q�uDcd�&z1չ����G�G��D�놘�?��g@�(:+�(�8���EO��Z��kx����;�O	.�V<��Ȥ��T���� ��[5�*.C�&�Y�R3v��NFk���ᶑs�qA�ʣ�� ˺`d!_1S��.�IȎ�ea���+��0=�a[�5<��}ej�"�Ɓ�H%}�Y�6���q�@�UЬ��i����-7��e�"��,��%9�� +A	_d���ha���c��bA�m	�-M=C�@�X���Ӡm�AdO4O�D� ���|��I�qz�zg�v޺�R0�!�Lr"������lS�n��P��:ѿ�}�T���Z@:�h\�xF��t�ZE���lݽ�A�h�����H����*(��ͺl��(w�`�E~ .	�r!��nF�a��(�Rv�le�p�lu�%�z�t�9{&s7�&�,��Ixe��
8�:)��lԟ�#��ԃ��8�549>3���M�O,q��"U�! �����X9���!��TS�6"�vp�2�c�<+��z���1�4a).c໖2<�I�C�U��BUxjl���>�k���!A�j�w�6���gH����*��RQTEE
Fj�h|���6����9�B��<��J��d���Xr�}&Í�\�]�;�Ss�&��GPL"�BK�>�Bb6$�藓�5��f�����t�̞VB�{�ւ�$�sH�"¯���$q�D �
�B�h��u�Hl,��Tk�ɣa��t��At��9�~�Y�)�	�Ngh�!V�S�[~�}<޾��`��Y�gJF�C�0�3�� S2AI�)'��J�
��I��o���|&V�YM/�y����
��"�E+�e�!s�"�B����:�Zj�!�<voZBh����\O��zӨz���K��k~\\�Xt$: ��a�������gZ�9��u�m��<�����1`�x���)��J#@�$���c�z�d�!��x4����+'	u�&�A{���1,��PBy�����w|��S��shY|?v)��������^��Q;B�K:��2H�\&�p��	�}���[���=/v�����K!_j�l�`Z�HwW��{����s��U�:~���*�uCt����e��(���:�D�NŸ���%wOI�O,����6lS��S��lt'`ŵ�4ӅAA�Bڕ�+��`
���3=�6ξ��b��Yf���/�c4����7yZ ��4*u��������,��S ]�G��|�Ab�O�� �����ݴ�~]�h�&��^�M<k�ҙ�	O�Ӊ��r�pH>��|o���D��#�f�|,ɆEA]�%;x|�9�ڲK�T��ImQ,��CcV���F�N�+�,�����x;��4�)>���Jt޳��0�ezoW��L�S>���Qi4����NS���fa���wW��ʥ�"�� �3�m�%��ˢ�8�>�k���M�A�٥��(>>���} ��
��%ݏ6����}�� Q3�
$�󃍯�Vd�0߁&�4h��pB���V8��Pb��	�%���QJ
�iypd͊o��]sqs'�g���G����9X��7�Ͼ�o8�[{K��|�a}*��I� .�I���@�{&�A��܅��� �Q9��+�@u�/�a={��1o�H5�p�<n}�	��=e)�Q��W~���C�-T���*����*^�U�G���^���}@��|�9�c.�X`p%�c���M��m[�V�#�:�L���)dIo����1�����x���#֘�uU�љ�k��8gA��,\]���D��ȀQ��U�"�����0sr�WǏx!�(�D<�2��Q譪�Ԕ$9�_IaV�,�|������^�ŊV5|�U�|��]٨`���`V̸��(�9H�L�����ˑ	��;��;o����ûF�J� )����P��zhG���T��S�Ý� u�Ho�Y���x3>KA�~��n�-Dy�Ш���ΰzA���zF� ��aXe��ĕ�dJ��賅��;�z}W��߈ݲ�{0R�J}$j���	`��޶s��8L�ۥ��Q�t�������Ş�	���d�ľ�����z�{=W��%#%e$�����b�zju�Z��a��P�Z���p/A � y=��f�q�Q���(%l-�q9_镺4�&�tk<i;!���o��N��d,{��6��'1��f&?!��@�-B^�a��[S�(��}���Խ}��0r3������eS]��̊���	E��j��UX�}Z�j��
�)��뫧�X�a5F���2]bۣb�	�X��'��3?�����2����\^���r�v�1��ej���_Z�}�Vc4�N����|C��K�� ������7������~󠧁.yGS���	L���'4�ʁ��K�'�� ����Yn9%�9)*U�T- �y�_F�E���I=oj�h�Z��9�$���!��r���,����
3��E��?��U�ֈr-)�s�e�ނ�J��~��hvK}��j�̓?�qk�>�T�bN<�/�a�@'[�]I�S����5a��}���R�»�Ǟ��̺H&S�����Ef�}�G���&����ٵ5���-�����6�p�ͪN$�zi��l}�/���\�>X>�gRm��-V+"�iP����w��],\��f_a�v��c�>���M��D�C�Sp֨�\�k%}Ku?Яh�X�:!f�4�*�&I��C��g@���q׿N����5�y��p*2D�iٺ�d�`��G]��	^�%w$|놆��˚��uy ^(��o�V�,$<
4uO��Ϋ���Esg�qH �`Hw�5W�P]�a��B8e���P��xn��jV�Ih��`?���V#��A��#�����CdMpN��� ��ڳ@ˎ(������6v'�ʙg�=��?�0�m*>�Չ��^Q$��)#t�h�h��9e_O�n��>*��5zV�v���@SN< Ǣ�T��K�\��$�L 7�����?MLT��#%�����im(S$T
�J��Qg+���|��s��8k��X��|R�M�:��l��֊���S���-��R��1��|76Jco[W>eeC���h/)4�s'&bQ؃���)�9<��1Vd�`o�HшI޻c�RA��!,%�{wz���4�D8��P���p,����a�TO̍ROЛ�*<X�Ȋ��@��L[���D�=�t,J)K���6U<��w�љ$5{@(8�����0H��X�O�u��}~f� +�*4�=��h�0h�.���԰|�u����_�bo�wd�I����N���>��_Qz2[�����P'��ě�ء��@�d�כ���\G�S��M�%��{��Y�/n=!�Ji�ΰ�9�]�:��&i{W0�B�(j��0Üw������
���R= eTK�-��j&|y��X/�!��;�9Sʥ����UZ� Y�QVK�欀��툴=U\S+ډZ5A���X�=�wC�:�C�`���=b�M1	,���r'���{�5�ĩY�L��`yJ�ڧ�j(؜�"�^������f�'�?4�k�� Ά ��5�_�E��Ϊ�v���%1�Y��\{T��cj'?1"1��uUu��2���3{�-a�<#����~ɭO��ְ� x��^2.�6�-@v*���%��S�q�g@��c*� ��@�ߤn3�X�X��D��Rj֢�p��wL�OLN���������YXa@@�0��̥�39U�Ja��lb6߲5_E켕cJ�N]���D�>���/9�Kj���@c�tcHh�y&%H��H���ܺܔo`5vz A�ɩ1�,
����>]�g��ڔ
+����R�d����R�����L#��q>��k�<1����k�:� �_RWġ{h\z}sH��a:ڤ0� �%�x���hXǞKȱ����»J�`c�]�X�L�#Vo�������t2��	9Z��R��׌���!C��d�Op��,�����$�L]uހ$evg�s��}�.?O5h�K��xdg��w��5��+���x�}-v�3S��U���%I�R�S�
A��ʺ�w�x���R�y���2=�|F���wE�K����8�s2��E��^����Ň��2bK�Z�]	7Uq�S��<A���Ղ���,.T.�F��bG���W([�;��B�W:��!�Y����,���٪`�{�[�Q��K��8X>�K�F�	��`z�maa� ���dD��4c��[a�щ�gP����p�H����+��ʔ�,+]s�|4�$Qg�)�>a�I��ȇ�ڸ���{^�,2�^.��<��e�n �9��u�m6����4_��0���iX��!qj�r�3��~�1�:Ԇ<��tn&7J:�Q��2OnGd@f���Wsýἵ.M�,T�Ą�,^�E��e�`z�r��CŹe����J��)���=�H�<�ݥ��\N���������4xN#�"���s<�%�.��w!�lI�Y�m[���jO���^�3-T��L�r�Ӭ�d^&���g��0sC�M�%D��#è)W��M���?Ԅ$�S�'U�TWYf&�HQ�<�sb���	v@�&_��)Q.�ٍ�1*�|a�=��8��{���L����:��I��b�}�R�&�ˡ����@F�;�!���,�3ǀ�A~��1,~������N/U.�k�{�	x��'���E���$� ��30!x-�#g4�� �%�
�_���.~;,��CDi�ʋ��U�}x��>m��c��T�>��"�A�����.']�J�n����,>^#���i--���p��A�Mdk�S}l�dA�J��Ŭ�*�V�p�0B�Ї�6�������
G: ��x��%����w�ޟ͙a�]�y?5fu�^��Ҝߦ}�����u:�� Wؕ�b�(��l��3�}�1-='�� ���_~-j��Uhص�6 :籽�i�v�8��-Y��tT�E �g��|֣�KC�p�ƀ�-9�"Z��<��yM�q˃�n�f����W�3)p1|�~�U͡��]QC� ��[M�=|��-���	��`����P�p��g0���}��7� �?���hV��7+F��C�������'�J+��[m��t4�\	���6e���"���h�@M�M���uj5�.
G��ʞ���V��{�=�*�A*>����>|Ķ���7Ň�2!�_����k�)F�h�Ԡ=�5F��=k�Q��f�O?��Tk���4�^:~�ĢX �!�9��,+�����?�,�e�CRG<@Zh~ʡyY9
�#�`׋�� �Ax!�B��o@ufW"��:H ;�E��eq<1,���iU�S<�����h
S���!��Afp:BD�	�_�DN�o�vI�$Yɐ���?
'���d,�\u*�05�G����P��eL���[�6��P9S�q�xYϱ ?�4>�.(���*�f>5m�F�Ս�fi��%e���}h�S�.�J�R"E� �.���t{�:��$y~!V��V�h�I�恍n�~w;f�E1�3c��:�r&��?� ]��� C6�$�g�fE �O��8nvAu��>�+\.�+��"��k��<��b�<f�wLV~��X�KE.�bu�X����6���'s�����{\�ZKV%��4�)�6�ph�.:~@�,6Q�>���0�8�Sۼ���f ��Ϝ�n#=�2�v���G����)3ܼ��Rt�Ǩ Z����"����\�����]s'j>����^������ ��Q�8���Ǔ��`ZǕM�> �X˵ q�f\�:\n�WW��	��lk�zĿY�e{��p�ˈ��cp�ƌ1��#s�&d@�yg���ف�� �J_m߁~.|&B�&B�_3���u��d�Ht��zF�[�V�z;�3@��?~��Xb4��9�2��2��>�vZW��:�"->S[�65���;&ᯩ��:Y�zC�
� <����42�s�2j?�CO�:]ҫ1v�����/m���S �')I�ե�PL�y��z�ι}��5������BI�b�*�)��5��L�X9 S�[�Ǣ�ruW������!����A�gn�yh����%���4>��߆p����~�E�&ߛ�zq�OV`ZO�P���L)�>r�{�������+�s�w�z�Ѭ7��~nMۄ�3�7b��K8���'��}�M��UZ0;r���*�|���Fq���6��#Zn��ظ��߄r�)��L%�cUH|�e�=�;�x:N ��T���Me�2��(1�r (2$&����Y�&z_ah�)Rl�e6yי#�I�x����?�3��������X��bA���>"��1$Z{�kJK���㲢�ۖ�P�i�}:�),�m��imM51ߐ��y���;u�Z8�� 2�p6ԛ����~��צ2u�&�w���spÞʘჷU�e��Ĳt�a�1������W�+��=��SP�Y�)����3aR�jW�)��I"L��Vx(���UVv��W���%�<)�v6�u����S�"+/>��vo���������
DyH��~�y��FU���	�O��z]�h-hĠ�Ô~����}�L���a�D�u\Xw�D��x�PP�CQ���}C��WB�.9���(e�W��Ñ�n;CC��zC�L,;�`��܈Auz�V�_�Z5�S2�"��i��S�ؔ�םİj#-��2l�l�k�Q	�~`R{aȽ5^��XЧ�bS��1�2�z-���a�VW�e�_DL�	?�P15P`�@(:��o����D���@7�(�����>�)���z��SErX%��Q���	٩~�M>���F&=��B�kЬ��5`d!�#	ܧ�p3�Y�N�
{����ɥ���t!�.����\�/[�(����)n���B��e�w͸Mи��gT�Hj�^�?5�8�%�o�m�jA�xW�U��>_���.27�w<3��{��}.^R��)�k�HT��ts���Z�'��2�cÞ~���	g���g��O�f���6B2ܿg��'0(t�o-��WK�)�!��7�z���F���7D�J8�k0ħ�j�1\�fi �	�{Ĉ�k�˾�(��q��ֱ�(�W~ nZ4nT���~���%���7¿���sj�6�Z?=��6jV�l�y
�k'L�϶�np�"4T�E�c�o�擎ѻ1�n��E�vP�g���rna�3���@l.a�G��'����E���ƫ��iQo�V����U�ur�!���m3�0C)�}�z�B8�4������5'��_ޜK�S��y_���@����o5oc���|����JFQ%�N�92��mdl`6�Fj����$_��8^ʂ]�m���}����|UUq9v�ՖĎ����YZ�2��z����N����Y:�lc܏O���AW��G��ĉ���B��YO
�_��>���%�KL�-1c�z�	&B�ƀ"��'�t5w�E>lh���fE@��H�J��B�)1�"*x�C�Qj<F��~��o
 ���	�I���޶�D�� �3V�dgƝ�*�2� ��C?xƓ~�����e�N
#�v��Ua���Bfں�i�}�B�v����1-W+B��D.#=���ҍf���Ir��`,Z-�u������`�{��v�dESoO6���AӣI�­�x�|�AL��a�̷���W%��;�H�nFGH4��0�(/��,cN?O+������?�V�֌��Є~���̎a}��<Uf�W �@n�$�} ��6��GO��n�fYaZ�70,�	��Y5'���*�n�i0��v����t *1��1���8{���Z�yiK4���S>�o���иkk���'Dd{MDٴR@2|p�)4�� �Vx�Q��w�Q'��^��5
0�"��w��ԓ[�-��0q����G#AnW�ȷ��v�RM�X�o+/R�[M�7n= ��x�h���"α����3�i���ϛ��$�G1���s�m�)Oe�a*���Km3������U��c�Pj Gjc4���k<�c�����ȥ�d���c4�QH��[�Iw�����k�g��9h궸�7C�N{��N��,}�&����B���j�0E�(g%;�J]����ڦ�r��O���)I��� l$`�S� �R��	�ZO��*�,Rdp��.܌��(6A���
rg*���U5����_��2�@� ���YR�!7^�-�K�o�*H��a�H�D�YjP�<gnǺ���H�hO>��"K�U�����R��\�3�A�,ҹf��I���a�TN�ULwB��}�	�&�|p��o�6R9ӄDu�dÉ��=��,��b=R� �8���;u�.?��<�[
o��r}V��PD����0�1��kǔͨ�i�=�OK��',ŕ�"�9W<�OdO�p��r�P�lo�m��ͨA׳'1�������4>JG�4;��֒j=�g1�δ����:���0<�C���( ��!PU�0�M��RA�>��`�ߢq>[�#=���J���Q@����K�j7��{��~_��{������i���-:�����4���Ca4� ���4P'/[��d��ԵU�]۞/�0y��ō�z*X�H�E�)�]>2V�d�|O���;w:�$�sz���q�l��c�����ϻ2N������5�H՞�:�D��8��@���?��ڗ|�@Q�Ё)�&���]#B�yz�2�u ���F�&�ڡ)c���;3�X�������E�3�f�M/$�,����E(L�Qsc�hd%;��<�� sO����D�_>��E�?�$�n8��,�g���<YU,��'5PL��/ag%W|�u(w]q��J�����J�S}�)���g��������E�EYs�U+�|;Eհs�%�]����s�K�ϱ���`3����V��Q0h^��h�=�����|��b	�r,iGȧ��P�2��0{��`D&��Ј��'����R�@��l0C��T��u���,�6{u���p��(]Z ����
�p�4�&�	�Gю�s�@��R^�	Բ��d�i���4LT]��m��K6��칩��FZ�qɃ�u��!���G
Ŷ]D1����)��A�ӵ:���ID�;���\d�9�8����t��dV��gc�g9Ƙ��F�h("�8�F{�Î��m�[1&Rڈ�Z�_+���l($��C�T�pm�����������\)�K<����(��!c|���gOY��o�ڀ� 3�w�R��H�at�.�1H�!�������C�[�?�%�%�����J�lZ�� H���Jxe�������I�Ϋ�ͨ� l��m-�@q�2��R�R��v7�L.^����%��iPK#�<��Si硃���~�� |�QۺR^�,f��set?K4�E�e��V�*�Q/tt�<�ɸg�j��,H��M@ɐ~7FF1�Ͽ��3�r�V
ش�|}�yT`\��b�޵�'8�����-$���Wx�-��u��MP���ՁN����u��οƮ R!Y����:ao[;օ:���%�f�$�4l)�&�
�tp?�(�i��W��N�����:����5\!�8L���|�U͟��%��<�$C�!u�C��ʽd����w���9k�!�݌��f2|��fH��C��F�Vrf�RKm��b:yĈ�YHI���*f���G�F�/��:q��b����Zkz ��Ho�����^O�s]�(7���x�n��z5����u���U"�K�*F+	�_�W5��}+) k|xT�R���em�A��x,���G|��vz���G��낖�l��+���k�3䉬�y��ix���n�#X�4��$I�%��=۰�	�x�!\:�$j��v��o����U]���V�%���v���+�M�>�3�����#���<I�A&�����^�w�"#�b֯�A���PҖ�.�Y�c��	�D�ZȆm�����񚫢&d}(W��n��.Y����9T�
z�$1Mj�_U��s���X&%��C�Ѿ�b��t�mr���2���	�A�.G*�rUw@C�j�\x�j��k�MoP>y!��0�oh�����n���\$�m+�H��ʫ�;��n��^�5ߣ��R`��J�)���>�~键0P3bz����_)9�w� w6�R,��Lŧ��T2���V_j(Uv�6�+L\�~d������.q�
<�kMU��M���}��&�����I��i\�G3��:�ʙhI��-��N3$��V nR�� gU�&�wT�
�A��P6{2�}J]��}��4g<�q���I��R��L�q��TГ����UP\�^��[:����$e[3�ܞ�Ɂ��r<��yPO�#!H�%V�2V�w�r%����b��F" �)_~	f��E;�0t�Oږ���0��:����ݏi�R�pl2i=P�]��o�-�u�/	Vmd�|K+��O�ng<���3�r/��q�x�>d�i^�%����	��߄Mҍf@��_d�%GzdXO��P\��h�>���M��rl�T	u-��ُ��s��ih�����Z{�7�k��#ʜ2�P&�(��`..?��Cy�6\L�b�p��扶��Z�kk�ŵ�+�W��F��<{գ%U�(�^�d��ޙ+����յ��r���ЗԊ���Y/4V_�zۋ�
p���O�S+��B`���psY�|���&��&�H%1[V2�m�.�q�'��؟����5L��f�e%�^���^�����E�rW��j�ى��A�N�O/�&�q
�N�`ǔjqX��}�����S�B���
p��;7���_.�} ���Ў`���>�y�ƒ�s<�i6Yn84Θpg�4����9v8��k�:Ef���8��;���vG����N+t<z0d��X�Ə��^�6BOeq:$�>�naD2D�01�L���h��0+�i�������)�q�#N,0�ȫ�=<�����8
k������|���ә2XH
��4��{ыUz:%��������aF��B�נvd��}��F煋m���(8z��ߩ~�Y�'��c=oi�������� 8��Z8��L���wKFv�s�Uې�O֠!!N��Ufo,����R��%���8Q�6���|0�RU�Ƨ�Eo#Ûg���5Q��|LRH`S-l#J9|����b�d73P�3]�a�׋,�Eβ��m��S��[bM����w2c�E*s�E�H�n�w抎E�������� ���ߢONo4���n*2��B�4ef&/)��~��,ݏe�Zb&�|y Y���>_�o�n}Y?"[�5�:��2*s���	Jf`B�ܰ������D𼽟�;`6�@d_�c�d8��4�B��7e��S�h�8 l��g3z��K�I&�r��+�_m����VCz�y��Q~F�8"�,�����txm��(?��۱X�#T�~�ͯ_{���� |X+(D-��d�b/
O���)v�D 4Zg�_)r�|�Z�¯����@�&3$gF��@��T�0�:�eGbD�lH����ֻ˦�;�W9��ﭰ�����[B��1�\��1Y/ln� )r���7��x�� #/���C�d��F{�v����6g���!�����C��6}�����`�l�04�&�aW���Y�JS����,P���^~�����>hc�?^\�t�Oۘ�h,[�iS��v�
M��筚8C,�:m�v޳ƿ�n$1o��i�7$J�|�&4��T����^���� �%���9�lQ��A��wuN����_@Qd�_i
�h��O�΀�GZ��[!ةAn�}�1�/g>ݩ�3kNab�K��O �#�J�7-x�O�~�ǿ�l�oi5�}�2.+y�S ���0��{��C�ڸ�o�o���S�,R����D���"4�<u�	�e��ey
 �AD�!�)��p�0G��Dx������o����Z3�F�Q�i�B�����L���Xo�_�����m<��̼��F�1�$���ޝ嘻ػrz0{_Z�[�k��������HO��^�h*�O�ڒ#NdvQ�R���$@L`l�:�F"���^�4����Ƿ�P�D��^���{��}�s��r���&��6�����Thd�-٫G�FIZ2	�d�kA����'�Pcv�rk�TT#�Ʌ;7-��9ډ��4�`�FE/x�!�;k� ��� �p�<дJ����۱L�t9�q�t%�:�nƠ�"����B�Oe���|=�R���
��#�ǖ:�m���]�.oV�;����@4H'E�D��B�^���s�����ӵ�9��V���4H[�i�����G�eor��}�s����G5�j���r:_0x��'_�
�~������[dA3p�L`�Ԩ����PleE�k��{,�3��D��,%�Gw��
�ak�T�?>�Ȃ���1�@mQd=�#�|�.i� �	8��̽��6���Fjƚ���.s]�߬���/�o�񡙌�(��[[�#0�l��"����{t%�!�.?����T�[zu���JG%Ü����(�b}�%6V�!�/���M���*��(Q��c�!�`��\�$���&�L��D�P�F ˷\-��$�/��,�㟩Q����u��E�G�|��$�n+�{�vy��-��eE�9җrV=ɧ�Hs�϶OY=w��6���c�Ǜ�{GG�c-7��vb��>'�W���K[{��1#3�hQ�G���=�#�������~u�ޚ��V6��tgs�L�J�l��D�u��f�D�OZ�FL��r�6M�N	-�����A ��=O_�����y����5�X��`��U/��]mz���D�W�����K�M|���OMO�Q����6Swz�ly>��j������&`J������6�0�Sp�i���cRҠ��K��)&��b#'� U���a�R�M�;�yi����� ɮ
C�7l�˿�����.Y���t�(-b»��A��le��E^�hd,��%���Ga�ѧ.��ո%U/[�Q�[#9ګ���Qc?(���Q/[�:9��!��U�;:��gb�CG��5X>���i!��}!�Ц:�Ç4�Ѣ�ԝ�*��W�¤I.��c��A���Y��>�N��[�e����݆��(���ܸը��3p�?�b9�\O��/�:F=��^au92yBO��.�-^~���Ϫ�˚����2��$[���g�=Tz6���NiO�U/Ğ�0���|��0fԂ�6�K�d:����Ғ^��n���HI�y�z��EZ�1�h�O6n���S(S�����h,�C>���{tRo��wǟ�q���y��&邞lx$�%:�gc�<t:Ip�D%��P��n�y��.ٸ�׆�u����p	����H�^�y�]�gB(��(�߻���3�'�>>��>�E�3G�U�~�L�۳eE,FA��c�����L���e0�G��kSO�E�E��gkz�
_����/c�i���j�0i���lz��_c��b�i;�P<F�D?F�"q�D_C7�ˊ�VOj6�)!������.�Z{��o.�}�Z�r�H=�`��\_{3*�p-���0����6�ܟB��9%f}iE�"&�����߀
�|վ�TX�s����:g��g��ٳ�YzZ�\#S�L����a>����GF����c:O�N�*XT�8��y�JN2P]-��,�߉K0�+֗�Z{)�J��q�Y���󯿤o�ߚ�Jx���'��,Y-e�Ϋ�1C�5.��k�j=���!��nn�1LBaf�|S����;]����s�����t���5��j���m���8�mj+�6��V�&N �L�P����{.Sp��V`4��tK�� jF���F�k��VS	T��I�о1"���R.H��ܫ��ET<�s����5Kk �e�[���i	�`��9�;��I CV:xC�{kE���RKWX�N�l�r��)sLp�H�z���r��\�3>�"A/�{�������1g��"T�N( ����O����ڶ\r�ov���m��̯�eжs~�.�ϽxY:l�_~W���P=R��  �a�)j�lP�b��g:F�y{�r)�Z�|�is{X���B��;��r�9h�4I*{�ﰓ�d�^�+�����ɟ�ahQPO�a���b�%�3{�qQ�a��JU�].>@�y?�/�/�/<�*�G�5�;��-૕���H�{�x!����C�����]�+�KA[F��i0������xߎU��/�=��-re9��0���r�&��eg�?��sZ�k�ͺJbAC��GY8.%�Ҍe]�����R�
 aV�� M*�}� ���=h�}F�� P��˲�D��L�b(������v�q@Сp�[��?�a�1ۨİv5̫\18s��h�l�<�j�!�/���:�۶�Q`kL�)��y:����\���e�N}X����T~�>^m?a����­i��X&�՚έ/DV���� x8�G�d��C-v޿;X�����ԁ=��.�گ8��x�,�;c_�ӝ��o8���`�Z��8��+8VI��d��<�t�K��;�ա�%]w��>��^��!h7����=~��9��R�w����<Hk�����`Q�����&H|8�B1�#�_1�[p��f�V'�`}�@����Ȃ��MJӿ�D�D/�C�o	6f�YM�u��2��Б��n�%���=Ԏ�dhF�/�.���If �����yW+;z�g�-H|�h`>�O\����q�]��R'�5 d߆yfC�⮦aRM	�5���[J��2���ɢ%k<�X :|��ӻ��f���)��v���b�:)�e�K�Wn���R9��	 ���� D�Ǡ
���5��ኌ{�J��W�ut�/@�k0��2Ebe��:ž��m�ٛFz�87���Զ]X=�{��*�vg�"Ϛ�86Z��cfH���ŖUY�+p�fӗ��P�q]GLV6vԬ�*j,�؝Ç�Q*���� FO�_kPv�@M�ZĪ���B����|ov>CTڕ��6N�G ���Pt	wܱ��U�[𦃳�t���r�ll�� ���;FG�Gh*-w|��6���Z�Y�y�������h`u�:I��5 ��q���c�_�u�#���*bNL=��&�~��d�c�N�>�;s��g����竎����4��I��V�*�g�y#��E�n���Ƕ��B4Gp#����Y��C!�]Z�~�Lx/Rz�T����,����5"��������H�O��6���Ӻ�����������x��Ɇ��KUD��ٜ��e�},�AV�FBfWEʾ?-'�m�G"���#���Ǭ�����Vy��ɛP����5��5?�A�dׂ�W6��<�ss㼿��͢h��'{�)z$u<]�怒Hdo���@�\Ī�{�Od|]�����F��r�(	�a�f+��q���t�~���t�t &����Z~:�i˚��:�f}���86��ls���叨1:f��Ǽ��S!,en��/eɳc"�*_���D���5	��]�]W�Q""bq�x����a�yn�s�=D���J�햦�58�f�+�/�Ht�n �?&�nms*3\���!}�w��l�HDXv��Ğ�M$�w&�%��dƣD9jAHp���L�#��d�>b��?1,�t���N�T�]�	�=����5N$9�1�b���|櫃�d~�������-��>��!��= �b'���h՜||ח�b�,�}��+Rn����(mǵ��M��:8&�<s�L�X��Q
��Y\Y5��J3���G\�G��v����:$��[-��Q���În)Ղm�������T<�-�j~��z�f��x��Q�UI]���5FY@�	\�iӌ��]���)�gZ8�1�E���X�v��R
�ߨupѭ'����|Q��Z����ه2�ta~�,�:��&�b�1�Ω�o^?���@9����r��-8�/����$��i���'�m$?̕0zj�s�T���;�(�^��<�%̘���]���b|+]���^���.����$Z��g���f���h@�^����ff��4�@jݕ@�@���x;<�Ty���֨��
J�ջ�����^x��ɮ���Y�������Z!�>���?G�f�.]~)&2ܓ��Z�$0��_�BG<j��A�^�=�q����f2�)IêH;F���q^�Kȗҩ#�:�Be�F����Z��U�ز W����n�[NE�jAr��봓%~�ؽH�8ih�������9�g�Z;x��_�\34 n�1�ƃ!�����f �ACG�ck�NZ)uw�����(��M���p1�1R5�rb�]	e)>� �QA�:���lp��L
]�����5��|�O�鴣ؓ�v,�^Z�ZGW���y�_�}q�:)
l�jꓽ�#�o�:x;��۰k"'B��thu��7���@/vc���9�H�~bz��E�"�i��f�J^gTxDR^v�q�2�����$�qB�l\�rT��@�Y1� ����I�,���Scb����^O�br���@$ĽD;A*���b�ՀC�j������|t	��o=>-wz6飭p���O�̖�4��ݪs3Zi+l)�tҼ��")Jo/Q1P(bU�?f9�;5|�?W$���Z8��(����f���W�7������M�O(u���'$�`J �zY-!�$�z�*f锐rQ5P�$(�^��. <T/��xm�Z��ˆ�MΆ��xݱg���\�� 	H Cp�C� E�9|����_����OGTi���(
TvR��i�3F~y�s�h�����窇�x�����Q1��9>5����� c��p#�EsI3���ED&� 6����?r�>�n�^U�9hյ ��g�����\�J>�:�8o��J��{�ҁ\з �*�}�z���$Y��׃B|���bTٴ�2[Y��!
<d=8�+d�����>�V���)�,x�kt��Ѵ�l�o&��<٥�.�u����[j֔Z}lɞ��	�q�\��|sM��Ю٨�~JB1|������GR1
z�1�e���#l�_d�:�e7��7~���@T|���2�%,4�:ԫ�����0��;������c.�YU��wX՜��3��_���K����ɋM�4���ԗGp�N&��p=�����S��Կ˘x��9�T����K1'M�$];�]e���Lp��S���T�5��=�Ƈ��v	�?ƛ#J�L��#L��D�u$K������ۤa>��gg�]@He��p�W�Ѝ�}����f�BH`��DC��	�����YN�C[X�v	�)�:w�W�J)��s0�?�އ���\>3.ލƚxm=���^Ҹ��3�T�L&�oJR�y��姳y	X���Y-��X���=�."-�|dnUʾ�? �8*{�m��%����}�#�Hӊ�y��9���,d>E�Uʢ�$g�e�N�m�/�_SL!2Ҡ��� L�W4|f\�6�d�$g��F7J'���V�gIz�����2)}�6�5[�p�{W[l�P3>��>��F�-ţ���2c� y*�f�fV��(bv� ��+5��~o�cH�����Fa(���d&�π�s�pg]=_0f�#�m�l�������kR��9XW�)�JnA�҃����%���~��!!Ew����;W��8Ҿlu�N�2hPtv;�璾J�m�^�x�I����Z� ���0��&(��m�',#�Q�����J��䩣�+���OQ��@1��u��;�ē�NbØe��lj���|�*}����N�рb���'��jT&�C�b���Q���ɎиP��X}�.�g���r�;_��A�l���u��VM=C����tS���g�w�>�l�'�H�|� m~�j@V<��8�!��Pz�`fةL|���ǘء���4����u�b�zIR�F�s�ιؓ�	ɬ1r��m�;��ۿi{�凴�Ɇ� �KC1&I̸��/��(�f�Z�?03g�N8޶%e.�֡ҏ"Ѽ��Y��27�Et�I-C`��Ɛ�n��8D%�m?5��˾�詸��"���T���C��<��S�֘^z�W���\�!��Q%�QB�6���(����c���Ú�����Y����b2�#�G<[i*���V�y�^/�I
�vR��'��*OSXǒ�s_�$�<��EA�0䖲����� ���ԭ�wFc������/m5���Qc�Tc�5��[G��=��y�ߩ�m��(�i��� u����_�p(����ʪ�/��8r}�d�R���8<ɣ���5f��5��&/����.f��~4�I���� e�^ �r���@
ύ.�D�A^�<4ųB�:� ��	tQ�,�>�\�CA̰`���#�3�>�C����i'�i>�:�x�ݨ�?���d�����K���z��s��j���c�s��Y����=B0�ɧ�nU���ؒ�V
D�+��֒���=��*��׀�	���k�lvt�m#���;��
 T�:0��=0_�a#vE��d�ckK�ͺ���S��L0H�F4?6��W���w�����+!~@H���ai��7�&b���z6�R����0"�.��M�q�A������׆�fG75<��$�/?�$�Hc��Ю��2Y׾'��Eּj�1|��3N��U��	�,�������X5�n\0�8+�c'b542�Sζ/N��7�K�2wX7U�Z݊����|o4dь��g��c3}۔�کѦ�QSɱ~uY�މ���Ԛ�\�\��f/����l{�_�	�A5���p�{g�i�n,�m4p���{�i��U��
髰:�&B1��v�G�^F�N4J����(v�C��9�S�#�vcѕ�`�UW�1ծ	a�a�E2�bBA����/a���yC��S%ȣ'%�b&?�,|*9i���ו��9#�)l,j�i�܊�q>'��)��h�3�v�ė��Y�@��r�x���Q$�,�?鹤ny��1O��"��5> 5eX�SK�"GI�~x#����&<���ZݰP|;�����&Q����>$E�T�SVy
�׎�c��[{����:e/+6T���YR�R���e�6f�S�J�}<�-����^�{}�X��7s y��r�z.1�S���r�Є*@���]A��n��;~e�AC���L��f�l��^�����;=���'�}����Ī��L��� ��m�^+%KR�fDv!�|�{���.��-�5�ڱ�jX�(}�ْ*4�g�1�������r�nj!�2Rd��FӪ��A��hV���I9�*�ă
x�4����:��ƌe��Պ]J��M�+�L4hLLw�I��dЦ;٧��4�"��n�=B��`���?\'��Ö�PB�,� �v����H?1�V�3V,���tR�������'����I&&4� |b�y�j-����V��1'i�;�%K�����Z� 嫑Z��-Qo��~��+���E�,}��Usnv�E��N�M��c�o������r-0v��cܶҝM-�����(����mT����� 1���%D�L��R�<O�'E�D�;�0Y���u�x�?�ȇX_��+�1�i`JӦ���0k"b��X�)��� B��fϛz��� %(��U�;rF 2�9*��0� �?�M?�b�C����3`����Në�T��P� l,�s��\�'�d�풗9�w���7E��37�)�شkF����K3�h��1��tl��Pmp1�dg�C�*_l��� S���֙w��ݽ\��?�����\ؒ�N)���3w�d&���叹3lޜI���36�^�F�y[�R��w�E�c��u(��~s��rR
�U{����PYh� 䦦����<���q���E��Wu�Ͻ�Wr�U`�Z�ɧ�B�����Cl+�~��:����5QN�i���0���vo�B���Dt�[C��'��A������E]Xt/��Ҡ�����0�������������_����o�
� !�bY�FP�V2�������dl;_�����`f��H� �Ԣ��As�+t��]����1 mG?ʵ�ۻW��;$tq��1��(�Kwa�WX:�v�tQX9nE0�C<��k+�:Kt�T����B�c_��d��g;�9�D������ �q`A,r�~�'�t�qԑ>�W�g_g?���ޏ2܊�g����MmU�}�h;���
1��`4��'�*��N�j��;�)�ѽn>�@�x�YF M���}�*��R���	��Hq?�?�C4�#A��f�
i-�F%֗��[�{~��.l{=����IM��#6w�%�vf��
���C��V�O��,�W�\��w�э~,��+c�2���Y$��:f4��#:��?otJ9[��$�|�6B���e�*=�#��@��,Pۓr�T��[���b
m��\��Ȁ~�d]�z@��\L�Uye��?��suf�iWO�%�
��&�-�-)��4����,'�6�!�I��W����(��Ĥ����r/Qc%�g%�i(���{����e�<�$��H���p�H ��N��_	A���ŋ-(��#���c�~)����濃Μ�'jl���C�D�2��������8>��_�t`�`HZj�	@�Ŭ@b?��4�B��>F���5c�1���%r�L&t)�!���UNy>�Ǩ�<��g6������:+�����)��I��$��IJ��:��>�{��A�{�w��E;Z�/�� �k��00�1:�o�-����z�����Kn%��x�mJH�ږ�w�Yo��`@�6<pΞJ�P�9�؞����9�2=��+!p[9��"'�L�N�`�2�m�����K!=f¾&�ui~�5t�3z�+;��e6�Q�&��#T����C1C����O�\�'Q��?�ޟ)n*Ӧ��	KD*�����IF�r<�z���Х�#�NuZ�X��ܷv%*��H�~p͖��^�Է�|r���: 0;#u�"�/�fԁy5m~�vO}�����Y˰<����H�b�m�vO���*	��Ǧ�Di��j�"K�	�j���IN˩��'ج��k�'����p��cu��z�Sk����-z�B�J�F�-.糛j�@�c�uE3 O�EVW�?䁟�nx���)FR�y��^�B���D���!�B��;o(?��/��C�P��1qp�CM��/ �ȃ�A����w�qGN/]Hg���<e�v�e.�Iחr؏z��n�x�ϛ�k�2��.U��}�y�̈�-	�J��<�J� �jI���i�#
�~>k�g��}�B���/����am�D�Ѩĵ05�p� �0r;�j�ހji?��ث&��my�7.7��dװa����ƪW�	���M��,��Ft��e~�/�z�;���jln�R:��K��_$��ȵ��L>�������[��I�-i���Xd�`�4'2jf��=G����$>p���� �M>u����1N�BQQa��x� q}Y$<˙�r�d�qI�.�K�EX���f�~�,����ޖK:o���S�sp-f'u���Rd�oc�e*�Ӿ��|�,j�¬�n�^@u���Cuh�|�^%�YV�H&�X���p�B`�zQ�s8�+��쾝e��5�+IBE:{@����(��D��=���2�4}��*z�f�`�P�0�ɺ���6�`;l��+5e�wB��a�}�X��y��W�b���8���i�)�u"Qm|ü��	��¦2i7������CCW3R$(���X�9�8_���8�,��F�yDǰ�X����)�Ul��o�ѷ���LYku����m{�*��Z��s�1&������"��9��պԱF�Sv��F��p�M����$)�5B���DW�#�7�w1ATc�c�X�>Z�L�+X����fԝ;�`���id���)G"+^W��@��0s�p��$8��}�N��r6:G�m��_�G��°XFƎ�}�ݹ��E.�#q���v���c>׀B��P>`D�� �3=��C��֨^&�N�e3��ɬtƶ�;������\�X�<�HaهU�!�9�#d������e/Д�=�9]�j�nq�U��ȱ��5F�`�m��v����~���Bf5m�! �uZpN�F�A|�"�1���N��[89�'��XWr�G��|1�a�}���GW{�SH��m���U�$쬻Mj߬���T��)����$j]��?�%w®������[�0ɿ�����ʤN���.�s�Ϛ��a���Z�rp͓����9�^>=ѿvk,�@BR��a��n#��.��Mv�kl"�@�mc�`�_<��C0t�/�"(�$2'r����v�K�6�#��ĨEk�E�3�sK��P�A�D��n��t��J��}�۠�Jzqjl]P��l�+����4�~��G��~�=�:S8�C���A=�+$��?����>?�Do�bg�%���-�s��Y��ϛ���k��Ӹj(�Xr7�iE�)��,u��q�Җv�HW�G��;�V<j��l�&M����7�]�3Mp��AR���.�t������R�AL>8f��p�m���Z\V]7�W~�c��!�2a�IE*� _Nb�c�ޏeI���$nBo��k�$����/�J?���W�K,��ȹ���k�5��M юb�3PǷ�P�/]-*N��F,��>��:��v~H�ܦ!/���w��\&�F(Oytx�f���R��xj�k�������^�����jO�C3�ؓ:���$=�J�th('��h
�#!�1�
�%/�:k�U*}ri��m8� 悌J`ٍG3��L^P�M �������&H�O�[�ȴ'?����'�I�F)��Nr) �8.}�����9�|�=��8|��.�����(��>J��^N`A%�o%����{�Ԡ��&�'�	�=[k;�-��)ȯ��n"W]b$��:o��Egs�J#c��">��j��7y IlU`���o-��{�-�g�}qtPf���R�w@�L Ue�]���ώx�2^DFg��0�䆲xӔ���5�hY�����H_SB�2ea�RA�ը]��EG�C�JۊO�XX/�8*r����(5�ʜ"��5fP��2�6��uI�g=�Z%U���-���Ex~&�f�ϖ9��Is��x�w���� �(~��?BpYc3�o�-%nh��-�l����E�N{������6�x�`E,���_O��.�X^2��1�����6A�h�ڣ�MH!2�TNw��:�������K+{�?��f��g�C����Q�vćO�l"�!cH#E���ɨ�q�Č�����Xu��Q�*�ZٱVs�<NޙuP�e��|�� �M�+��/ ��4F�+E������?��ɯ�gLo����4�d"q����o�!��^r���r���LU����*�S��Eh�%v�n�X7���^�J�{q-��%�#l���o�N����Q�~�`�D�x�_|M���Bg�õ�U䅀]l���7����ޤ4Y?n۸��t"P5����:C�%'��4{���(��������ߢn&�>���?�U�SRߢ�^�����<�rg�z���䶑�X짲����Q8/n��I��53����@k�~{�з/�1����"�VT�2@NOzz(*�؂U(����+��Ƅ`JwV���8�ܫ�K���8,St4�E;<�G��iԍw�H��C*��PT܅i�&����p@[�c�0�
[�揖� &E���4�g˰����`� Ȫ��k�<���#B�o��E 3T����6ؒи��{7$ڜ��m&x�D��>^�E�1�֤�? "��1�����x��!�Qah��#��gy�H�y�k6�����z�JL�|[A���_hC�y=	K}*]od���.��iY�tVd6M�;?_m�3L��'&�6�����G^�D>�z�>����������@I`N};��lg�?4P�;M�EJH�_o������s��z�Oɕh,_�}M�.h�.*�_#�qv�^[h�:0;��T�}�>�KA��ȫB^�{O�� �H/ rq�ð�0q�5��!��u��b]�
��
w.O۲Ӆ��b�W����>k:a�R�1�����\��M�d([���Qh������Lv{f�z#����kя}R����%1�Jz#�B{О�����}L�\���՚�M�e!��h7I�b[iM퇾�$��^y�9������oG��2�~�%�m��,��,��h��T�|o	#p�+�WxTl�g � ���7ڇq�ɦWNx�$��Mƈ-^�}�?��;b9)�N��<S�����K �mL�TvGt1�H��B�%�Y=M~����W�g,�g`9�P���!��L!���&�#\`��̹���w�RSA,62��SA�l_��S��À,"����m�E�F\��]�39!�K��*�<<����p��8sq\��!��݃��<��Ɣ��5�&���sa��7ӧO�	��
)�5�kľYF��Ʀ^�f�\�@їJ�}�"=�N��=��^Հ�c�l0��|� �����9��(�>�BAH�QV�L�B������V�/X���؇�쳛$`֎�P?�5m��կZե��"�Py�H���O? ���C�l�Z]J@��U}Y \~���>R��們��m���@���i��NT�1`��9���KB\�8����}� 4�%�P��'���0c�		�G�KV�©�-2%�KҌ�W)���#>;�S�G;��C��VfBz����ǣ���u�Tހ2�����6��Б�z��0�R���������3*iٰ�s�_7nڀ�ɪ���U��N���t$%u�\I�3]
��>�*��]Xvs���.m��,~_��I~���C��fI�b��|�5�9�e8��!��=?��!���������U|_�r�D[01Ҕ��A�;��<�B\����D�f�H�((:�J�}p(X:_����Fm�O�����O�sR0Fg����6㴋�4 ���iN�/��������'⻊��sfa;�#ߔy�P���a�-ع�+k&���1�`t;�z�t��xd�3Yt@9� *�ˍ� �� �޶��:�P���	1$[�ǝ�݅���8k���̶�93����Q�M�8�,*�	)4�ad`�]�}yH�.���,T�3��;ݛ+�஑22��C�����re��`�� �!ۆ��*��_s���:}��@���غ+��c�UU�J���`=z���mp�:��r��\8[O��AX�*B��(���=?�3����[����e$?o���A�O�Rms�D��%,l\K�!�đp��D�]������CGj���O�ZO ���dЦ�����(țҴ����ι��E�����M��0; �.I�A�2���)�-��$n�E�����ۊ1I����UM�6ۘo+�����`�nď�?��#����s��|��Q�.]��a��� {	�m�0|(z���SWz�(�z8��P�L��T��Hs^[�[=�3�����ѓ�1��r�Ʃ�.|D�K�x����N��G��u~�G�=�M��~��X\���3��JjH�D�S���"��U��>F��<��Β!�3i �����;�	�b�O�l5eW��DE;����6��}�I򑞀�����������>V�ɱMa�N}�?�X��7�^�:=R���ScP0��G� \�r��Pg,�.��E�A�����d	��J�,߆����%3��hVg>��TdK����Qڬ�:��ɂ�4O��j�TJqշ�M回BZ!���Pn�p&�]�y'O�-E����܆p5=o�F�6}I�B��6Y�W�,!,��Ɂ=���w��Mz{Y�"6˕{5>�l���hS�B��t����Y�D�Ͽ��v���{P����A����t�>-B��?�ܫ"U}�sS�� t^��4��1������ն�xhN(4"Ԫ�����Z&�� H�+>�I�~Ra���ve�sC�� �ȍ?T�|�=}%@�k���i/�rG�b���Kk��ä�WU@�3�LʯM���o�.x`����u��ƹ��MvY>� �m�$�e��%��}!���d��%��F����Kg"��^d!�m�� ��X��=��0�aH�R��:5��.��@��v>�ą���>c`����#{:�an���"E�[����Ux-�B����<< (�T�$�t��u'I�Vw�AA:�\�h��L_=#�и�:�z�*|�r�_D�"ߦ퓒V�m�[J��\�G���-�Z_|ˡͩD�sl����I  Z���SK{f�&MWCu��6{qTGM����|[G�#G�z����Ri��\��7چY�Ok�(�2�ऍ��U��vwFL��힧�uk̮&���k�f�Z|o�-v�FQ�'�Z�d��k�U���%�,��[�Re3��a���/�V�w� ���J�R#,�q _���.��K�����
D[�|;�#$��S�5�lP*�&�j��o�"=dTx7Pm���j��ISRih�?��^.	b���"����u<s�&�L Ah�3KW��v�G�5/n�O�5o�;��59�AQ�1�u\I☂��3�u�x|��IO�?�ШG��$)�d��Fܢ�� L��z��)	�1�����O&��f���D���*�G��o����ۯ��D�̪���P-'�֗z�T`�L�'�F� n+�ȫ=d��2b�,kٽ�v��>��M0����!�ؙ����<U�m�׹�B���|�e���B��h\^�M9��$��	5����;�Fch�X��m����mqc^
y��8Zjf�ɱ�ܳ��Zf�+5@�Gp�Z˿�D4l����uLh��!�˄��u�Z���'|>���H%�w��J�p���)���lJ <Տ,��=�M��C�G� 7�~`�%G*Tz���6
.)�N�n��I�?и:q���ub��YK9I�2$z���6QM���D�"��ݫI5{��A���r�> )�V��+mqoO���O!����"������[��L���flx`AB����CL�q��������ߩ<�|�������tu�'�_Oa���$��h(>@����_��<�� ��-�TZ˘mͳ2w),S�e���53/fO(�F2^�(I����A!F�&9�v~LV�ûdRh�_8��/I���P1f�٤;ٱ��zy�8��aPm�i���<�š�eJ���Na���i�}�|҄�9�1G�P�gas8	|�F��S��1�eJ�.dUh�:�|���g�rc�Z�=6���������S�X�A�J�<�wkg����CW����vG�S�-yT��
��3A�th�a7SD�2]��;�Z$��hF���b@{������J�]ȓ������d��$�����7�Գ�<wL�7�4����{a:�V�~��M(6yР��rv<!������eHp��zkd���3ka1'�Q����?;��l��;P� =�	u��1�@0�z��b��ʉ���������7���	n�<b|nm��&��^s�V����*�I��<� �����l�)8��7ֻG�б�����G|f�;�s�WH�F.�*�Fx��	6���Q��o%�Ǯ_�w-��X=�&#5H0Ia<}ⵧf<�7fe誘�\�!e|�� �9��m��ڛF���	-2��͆��j��Ҿ���-���)J�~,l�Q����t�0mA5I�=z�E�i�?4�$�ayԹ'�\���d��Ԋ��5�肍���_G��u�wP���`OI]LR�&�ܙ����9�����K�����%>'ZᏙ8�hC�x&��3*H~Z�]�uA�g�לd�Y+���o�C�V��ԻM��˽H�d�O���~�����F,���ȸBK8Y qo�yCG� A��G2�\�� ���������-�*���-�;g�mΣ����¦QK��煐��R{�� M�6d^��& 6 ����xV����
8TqX�.ӥN ��7Я=�\N.�/7(
�P\�p�:�*{�25�Rp�L��#���t����t-��}���v5sԾ�t��?��@�\l4��5zq�ͬ��2�T�+��
5�lFR�>Y%�YZks�VkΟ��$���9�p,Ǜ��f�23&�����Rn��� �tZ0���N�_!�dC����=��Z���J��!�\I����������X6yM�S�LO�c@v�R�����������2��T��{�́qy�T��F���q�x�� �]�NQo�A0�!��l��鸧�<���xԩ�w/6[�(v"�{O�������h��.���N���%��%gA�}	4.G�,z��`P�6N��f��q6�gכ�E�$�v5h+yH~�9�A$�����M������4|T�̚��*�^�"�yA��u�l�d�ک��ﭽ�
�<�����+}���5�4'p��g��,��*tI�`]S~:)o� ��z3���ނ8��"���aL~��][�C3"��I����'&�o�,<L?F�N���CI��j�>�;F*�ח9*Y9������w��!�x�L�`����9��H5��k���O�	j��ZO-Io$�ձ^��D7�6�Ԏ0��^��ۿ�C<���O���Hll�B!�>o���ӱ�_w�>��Cz8�ˁ Vf�*�Kz�d�,Z��B�M	�'ؐ`)K@��e��	�0���K&6����]�R�+���+��fS,��H+�*�Omvb�t
�D���!e�]7��W�JF'tK�z�	Y?v�����8���F�!&=o��M�sL��}]�V6pt㸉L~2>�[7��)�T�:٩�WR�e57�)]�IaZ?N��v�����WAu�2)���0��	���9��.�`�h�!6�ҽ��]�U0_D�cν��wF��V
�8�eM��U��[���s�s-������e�[�����鶌3�hK[�������g�\�%��x����i���JV3�q�Uϐ]t�=�?�$귵�8qQTśJ�C֌tFI�6%U��ͤ�+P'1��cu�j"�<("*����?r�-.!E2҄E��{�{FZ���%'h1	<�Ļ_2�c��bҡ ����+L�>��[1����v�K���	�P��о	�z����>5g(��8�K�S��v���"�� �#�^ϑ�mT��m�7��4���&�U��,�,3��^�{�k�z�ل-Hy�X77E)Ճ�����-���:.�5NI<T1Q�����_��
��a�3ܓ^)\=�&������ ������h,&�U���/�܁���F��Tj�A6��Lm�ÊZ�:�7L�-���ݥ|��l^,�o�����Ƶ��MK���k_�
�KV�ftRc�5��+�(V�5��#(��6,c��'����������T�0��e�͂|�K6�"}t�Z��M�x��yW�!���w@F��Dȓ�����r&��VS�񰐷��4}���VTn:�B�F�:"��3 ��=�ǹ�W��c���8RF�C0��d�}�D��x[12�oT'v��.��z��3#k��/vxR��F��+��T$FX`�0�:�3�����:�E�北1݊�͢�*��4�(֝��,o��W��pR�����-�_3	���U���p�]�c}�`�H{=�KPS=��d7�;X6�y���?����8� M�t��Z���	T���~��z;��p[�Z�P�L��`
�e�|~�E���{6�Q��u6�_������]A{yAI��[�w]��>jZ�v��"�9���AV�1ݥ��g� (���{;�jf�,ϛ���H�32����b��4�p���]T�V��wS���df7�k���3мt�%�W��NY����wn_|�>�?�a�O�q}	(iu�6ձ�F.!���u��`7B2�e�y�u�R3��)-��䳲����Y�z��[������ִ�D��R͚}M�}{��|Gm7�G)c1R�nw3�)��"!̈́��u Ip܄�z���wFl���uKe�x:8|��
����|��*��� "o��C�s�ݖşb�0�ZWY�ßLX�H8�X�+x�;4�MX�X[�,���������)L��q��.W�![c't�O�E^ͩ�"����wyg�)xZr~Ѐ����7���(�������ӎ�'�5���M�k�a�n�����uG�+`EY��A4moq`���a�#Ȱ��u����$���He��� �P�l���cv�BM�/iJ�o��+��Fg��xH/�=c, �^�������a�4S2�+�v)d��FΫ�@��p���O�1���1�l���C"�XK��뛠��H�-��w��
�i��t��0�����hj�~h���͍��t �3��U��W4~�ȣ��A��q�F+	��LIAs!v(����u���K�o>�Tpnt�x���̑��6�j*�v�g����[(_���;��x�. #��ޒ#�K`�2m��q�(���HR�>�g�j�c��p�|Pe��un�_7wN%҃1�_�Em%u�DI���(�pc����Q�s�|�ڥ�DC�M}%���S�ۭ[1�@&�������fL��Q�5 /��\�U>�ƛS2���{"A�g��tQ�{Lߥ�&����렂�#B�vm�Ƕ���ǉ�C�U��ǽ�˒c��֯q�[kv��.zf�E~M�F+_�x�<g'�܄B�����}j��J5S����U�Ԓ#-
�w��&�F��j탇�z*3��륾`�*��S���q&��.�x�ޜ9�f���N�ws'��kO`7���(�� �#a4�❞����jg� �'�j��|1��e�p�:٬J�����%�t��3z7΅=ge�
�Z�ֈ%�P8χ�<�C��m���'bS��A-��FG!i�
����hh��u��vqE�q�1��Va=�K�R?�r��9u�)7��[el\�x�Z�z
u:�y����^�������K�����χ@ĩ?��X���O�C��Q�x5	zY�K�LBV	B��L��(�-tT�b#H=��˖ٻx���Fu(R���\�G�钾 2��Iє�ip�_�O����dM���$�!��x�n�W<�%N��\��TM�ݐ��Ϗ�f���v�p0�����]���g��a��礭�iGj+���I�ua�P�ul��N�^�W��t��R[�ɠ��-I�~7�{�-0�=}�k�p-�D��ͨ�E*�ǣ
-:� �)M�l��������I�����؞�׆�Y)�Y�n5r) ]�6Fr*�.%��=B:z�I�e�.�)s�VMq�*⒛ C⅓�2p32Q��`������qo�`�ďE���o��U=��j_�b�ƴ��E���,Ł�l[�p��;,摃M?5b�j'A�� �s�R�����4��`u	�O5��d��e�6U..*44Z,~����o��e_'�c�'3F��m�	D����X���r {��\Go�6�M��i<�A&�H�<��C8O��O\aFR+
v'ҍ�h����R7O��uSI����3<�'4��YFɠI_袊d��t��7(
$�-��+ɇQ<��x�Q��2�+���#��B�|S.�(i4�J /l�8pi�ӥ��0�[�#$�ˍ�_�6%Uv=�����z��Y7V	�'�E~�L��1�7&�Ƿ\��Z���s�p���|�n0�Ț�;�J��MH��)W?�Vy:�b���!�{���H�w���mcQ�����z�G���J	v�Ɉ9E�~�*�C�B쎮����́������H.d})C�{�&��^V">�=2�%L�*���uK�݄L�߆��R�NRV�;�B.� u�EMY�����c�,		nh�������]6���	X�i�s���n�T�kޡ��*(S�f���(�ڠ��K��"�T� �Ha.�J��q&���2��\�D�U, 3Rm[�����Y�g�Zɺ2x5���s�O܈��vXH�5����Yv[��`!��7=�w�g#��$
���D�,�D�_�o엯���K�yz���IJ��H�����E7�>�L�	�$��zxy`o��+m3D�Wi&6�����n�ڡ�_��xk��nY�:�*�����#L���	x��o��3��o�r_�P0����o��F1�k�n��/�����(�.v�uȇ���L�;F�"�38��k@�4�|�@�_~Q!�,
���H�4�r�/2Y��&>����1YN$���E����#�����}�̒܅h�n����v��sH��@�á�?���G\������g�Xj+JG1F�V����%5���Ϧ7�6*6����}��N�!��Kr8�����b�#N+�)o��-ۏ��t\�1y�5$.�0����\ģ4A��)�b�>	���_��FOp+񨦺�+s1���v酒���ԝ<ǐ�|��Ђ�/3>h/�.,���U�Q�#ո(�,Z����K���.e-���狀�)�yz鐚r����9�]l(�}3BA����!4�>�f�q��O�`]��٦׏I��8�
f�(���e��1<�m�~XN�c@��e�A?8��j��;If�J.<���d�AG�-�i8�2��<�z��9ǻ�%��D2j�h�w�ߔ)�}�6�����]7R��X��̡��i֍�V4�9���D�H��&�Q@�a@�Qw���y�|3�'����"�
�A�kQ0٤�<�;��ϊ���]�ۂO��b���.��׿-���ƛ'�d,�a~����Yz�������.��Gީm�̕Pد+�V<$}EfT�4�3Gڍ�dG#w���1vf>�5���p��)�*�/�.wE�SK�Ȱ}�=<�!8�DXkU�DȺ�	�ć�#���xi��J��k-��H�xEt�=��Ó�#[��L�t:��Lӱ��b�.�Ĳ֩�E��H�F�����K}��L{7:���D�vƯ�K�^��B����2d�)>��n.(a
�P�}:&8	�ӟ9P����=69�W�Z?�����Ε�5��]���LU#d�ȈW)@�W�u��'پ�-h�T������)=�$�3�}kK��s��|�,<���A�c �/�;\F��3�o%u��W�9A�=��6��O|�;B����#{F�-������b�y�9�S�),h#7��n}�Y <b�!����!6&�{@#�/^0��`��K�!6��JbL�,7��X�WY(	�I�b� }��Yw#�\�d�N��Ht��ƛ-���e.?�j1���5�F5��dǾ��*��3Yk�R�#�!K=�,���E� Lr�ّA���k������P�	�(܅�%'V�Z���aش�Z���#g�֓S�z$m�B�aC~x$���^���,nN^w��bLC��s{�y �����:B�ɱF��=PL;�/�u�N$�����T���u&f�ȲY���	�%k6͋�3݉?��K�8[�'\L��c��6��Ucv,ҰSH��X�2t,KՆS��-�"��+E�2�>�#�4�`sb�nj�$��G�-"N�Y�k�E�υ9��n͒���q��.H��!^%�ʪ:���TyTS1�f �H�!d��a��pƭ=�v<;�ճ�g��~�TC�h�%�R�E�)j�U�ћ�Nmx�O���sa�o<�?���]��y�9�:���PXC��rW�>-ShY�[r�/���C������Q�,~t���G���A�7OJ�>|`|��*K	+��yx�OC�#h^M��S�A�X�m����X,!����3�t-��+���e�������R��x2�a+�	��]3�e`����5tX��+���^�����?��M�C^��@�/�L�⇧w�5ێ���v��Ç�Wt����;�,;���y�gX�C��A�<DL7k�=cW^�RfF1�tF+���`7�`�H]�X=�j�]�Q>8�w1���?; P�%9px@DZ�2m�y�<������d�\g��#n��I|�lb��%<��G���I��N*S;H��z���Xʀ^�z��z�FW��Ң{~��w�1���(f*�%����`��
L��}�i�,�2!�y��G
�@��%*H�q_5��j��G��Y��	��t�^:(���Gh�L�)DF�Ho�e�"�0�Tڻ�{�P���������� 9`�ȿ�y�
x�̌U[�j�m���C)�H
�1��	eIs�iS(��XfC��`��Ǭb����"�}_o����u[e�k�AN��Gw�V4`�B����ޓ����kQ�-�V��ʪ�@��_$��v����~\#� cm(m��]��Q���9{��oV�k��(��Ꮴ0�	lE�7�jv���a����?�Q{�PwI��ꏡt=cb8��ľU�p$Ş�1�$��Q��gI:-6�Q;6Ԙ�G��La���A��=N����c�:O�"��ӔR�pq���t�V��I,#g��'�n	�w�p�΃`�&N����Qr�>薡��<v�K��Ă;�uq"��S*�J���k����*,#'���)��$��
�V^�{K��k���3��d��SU�_]T}����;��b�u6�6�.���F81��z�LR;G�l�g��O�J5��сY�=����c���yM��?����W��Ѿ����4F]/	_��*"Ӯ���|���^�|<���l�w��
��F���H"��P=�X����3���������C�.����9�Tz�jE��tl�+W v��Ƅfe����E{-�L�q�a;����3|���n?��9��^�T���ׅB5�2ժY h��
ߔ~���*�OW-y#�=lq I~��Û��b���ϣ��Py��Iٚe!�(�Z���4܊Y.wo�����Ƣ�~�KH4`G��c��IVCenKR x��Rf��%�O����=�'ž۪	 Ӗ�����N��BO`���4�ݛ����	�Q�ƈ�@ÖW�ч�7�֥]Y�(�N���!XZHaDxt�y%���k��;��;�O�W_�G���?�"�ua�����oz�F+�E��Iww�p{0���8���U�x-�����ج[z�7����� ߉����`�2e.�M��yqV�޾%�Q3�z��'�ps��} �gaF�y5!Rf�f�Z9�fR�&���M'�)u��r�t��Az�N��cp$a�+s�p�V���q����x{�Kq2��B�ĳ���յC��-���[|�*@7R`M�W(����u�� �Uw��~W�5AG���DH�v��m��׆��tk�����Z�!e��=��*%�aA�涓a@����֣F;���@���
^F�n���
U�K�z�ۂϠ,����)�L�J��:jQ��P��)�r�,Uc��}�Jy��@g���kI�8���i[Ԙ�h�n��8�{0h�/�v��K@�����؁�𝆓Q$;���fQm$P�4����WB��g}pN��~������e ��>a!�������Vʣ�-,*��c�-���C	6�`>f�Y��b@��x�k�\!���F3���믆_��ڼq��Ou�%`�t�,��z� ̩��2]�yJ�����~=�S*�$����.�4*����c���HkЖ����`γ�����w����~��Q$a���"X9<��� � ��� ����U��W���w;�=�������P�����=-�{��/�(p�׵0��P�OE+k��c��>'i۰��ZIW"��;��I��������j� �s�A��W��&v)���Sw��Ÿ�:��t�~(� ��~gbD;G��o���O�O��Y�H�=Ÿ�k����-�KԔK�So�~�O9-Cs�E�|�Zr�e\��U������ๆ��H��0��_�=[�WE�@����\����'#�!��w|��l�����j*�T��|���ҁau�r�����(F-���6%�(����1̺��w+]1[���hk��h��@�S�'h�����wS�5����.��8�	���/DI�..�%f�Y����J��M���R�Y۪�F�+�2'jV�{����	�I�7���щ���H9��ĵv���N4̷����w���8�m���z%Q���z���g��M|bܾ�d �c/���D���Y�L�{[U���Z/��`�ۘjY៰�W���I�
�[��`���UY,B̽yF㕺�i '�gL�Kd8x�w'.;��/2G-�*;����P5�f���@�����uod.|׸����=���;l	qx��:t�!��.�I��N\=���-p��;�ҨC��|C�U+��H(�:�XfOͫ�%��Hڜ��?�����Ӳx��t�j�xTY[��%x���+}κaP�F�dth�hEh���_�����j��j�5�=B�V�~���q�3��o@!���?�Ҡ���Qra裏���hAu�b0U辯>3���c�O�������/�w�����+>���E�@�0�	�IW�N�n<J��BC!c������bN�{q�L �^�]F���;ON���9�d����n��eXFJM��x�_�*��u��(L�!�f��]2���,���ŕ�C��O����=u��FQ�5�}y�yh����1>��0h�"��h�O/�����oh�.�\�Uw�@��pE�w>���Ru	����1麟}JN$o(wt��m~���`�E<j��U���l�iC� ��.V���0��xu��.��Cͼ�P�ux&�,���*KMd���Y6 %�X��3�S��6�����^���	��g(ߚ��f�(D��7����(Nw��), ��B����$6�3�~�1�I�(£rA�\ޛ�I"��J��`��~�P�iE���*[�����D�٤��J�~�S�&v\���Rm�Fv幾�T����
�t牗~[����Ʉ�{���櫗�����٢:v�ٴ��\�m���P[���e{�ɻ��#]Yy�_pbfL|�o�޹�ݿuߒ�I>6W��>��6�J6���e&��vͣ0c�����cu˄�	�>�!��Az]�Z������&,}8ǫ 5�+���]{f�G4��p�֭~�/E�+0������Cڨ	�&=�+b�_����Ğr�~m�R���^M�Q�
��ًá�@��4��)�;`5	�\v�Ü���[4����*���.l{��Ɲ�i�($���AEw@�>R�e?�p39)��Ғ� �N�0�y�e���o����#��Q�!��MH$�	��Ӕ��*�Z�C�!�/Ԍ��z*{�Qձe�k�KxB��,��\*�����<S�|�f�^T�j����5@CP��Z�p���T�-<�O~\(Z��Y���,	B��u���c�;Y��WoEu��#X%�Ý㊻�����YE����t3�1*zC$[�~G=l�Vt��c�zZ�n�zW��Ǣ�i�ߖ��ڹ�*يtxQ#5�-�*,.�t_�����-L=�H�H5����/2w��oy��g����#ْ~��'�i�fS�5��-�l��i^�2�8�4	��1�֔W�.q��v�����H�S�r�����x��㽾*����}Ka��R�/ �f��`��N?&D��,v��(�d��¤�`�H �+�0zKh���(�J�b�񥧭Ce��v9�<W �y���3��|���N�>��T��H��Hk��n|	��/tH�$�@�؀6i �Nq����߿:Vs'��%�dt#������	�X���>&�R��oG���.��٩���H�޴�|���2|��(V:��|�@�^����T�b,�ȯ�h�qT�57m�x�&���sD������
���U�:����e���4F�-�
�����@�����W��F��M������K�)����bӠp~0��t/^Q`q�#���?)�q>oKYE����9��o6��RF\h�H`_Ps�Q2��)G��?˱@���m�7���j�2���56�����:��=%� `��c�օP��h6RA���k��X��
��=�K���[;���t�ή|x<�%���#ͽ){��}��	��D{�9P�֎q)
ۈ^̩z�j�ȸ,���>�aCu��6���Z~�ԓ�!�ӿ�"�|�|���ŵ�&�������bk�+}��W��H\�i�d*�Q;ӥu63��*�y��������B~8�a��eD�A[k��:�v��#c,)���iԸ������,�u��'ԍ�'\�6��%�78����~�%���X ���R՝ YtC+�.������VH��:��B�AM/xa^5u�TO�R���o�+�=�����Z��8lp
�C�&�<��,��@��l�H>nP�ӛ�hZ�8�帖�֤�'����flPh��e�1 ��EW�ȟ�m����hC)����R�)��E�5!R��C��çăb$%�9̉2OdN�@K{��}/9Ŕ_E�'��c��Fٮ+�����CAIoD�����Ԟ,����t����:�)嫢��r�k�Kcf���''Ҩ�y���.��w���+x�f��|E.� ����]�7�]B�Օ^ʹ��c}E��tI�;{|*�Ld�i�뾚�T��a�+�$Иl�ѓ��Ǉ0�/:�����q5���1��!hV�M�[����&O����g)�i.��.3����Vl��ƸXe�'��{�N�!��+�d���݃��<ȣ��c���~���r4�3��,����z!��.3v$���Y٩��,�YB�w�X�����$6+�X��+�:�$�;��R�������`�)�ㅒ�]i"��ЩjR/P�^hS�n�7����C��0�b��9�4"R\�k_w�Aʋ_<���V�'h����+8��Т�cmeG�]8�ڄh�C���_f���?q@��ȑ�>	y�'�_	�I\X��ґ4��Fi�vv��(HJ��i��f�tY��tB4��b�6���M��$�����TAư�b��J~E�%�����F�wԎ冫Ò���h �r�:�y=��R�)J
P|M	-��VT�pkw�"X��O��^$8��f���'B��-N����_#avuR3h���.bc�Y3�Ν�U<��@�=F�x1��"Bx*�����OT����
��w�US�P�2*�S>��>�5����o�;�Q~7�x�Z(�Ǭ�%q������
�,��F�ə�5��Tȩ�Y[�b�G+��f����/�V�iK�<�5@�� B���+�4�*�wr�[���-�� �?�j��eA��HS���7	P�⛊l�_p���`Ќ"�	�1���tqk�+�*�� �JM���g#&)�����v����;�%��=�a�i1y�xdu���rʷL&,g�&�\|ſ+'��>YF���8�x4
�A�R��u��̞!>֓��Zs�e��x�d���'�Oi1%c2P ��~�E�}e�*�9�s]��	]yk��o�������ˍ���ӊ��ە,����O,����B���Z�rN�x�ǴE�	w
�]��+靈��XBh��v��%�Ѽ��� e��n�@��;K@E9�
<�xo���zك����Ƴ%~���0i_���"�9�)Wå�i>��9J=�����z'wL��"&�g��9E:�L�炲�m�W�2~XO[Qӭ�c�s�~��r�x��+����VA�i�]s�TfOPn�)�����d�"�QO[��&�v4�B�w�M��T���X-x��hR9�-9��w��g�h'O�+��Xg.
����V���-<���3����F,�W��sT�r@��r`"��x]&����u�Z��ﵸ3�~���D�C gݪ�U+�:�GJ�f�����:5�#��
����Cz�ι���6�r�1@9^�`f�>�q�_�9�����v��?�g�o��HnR��~۠��k%����%ƶ�:t��EXw%q��a{ q<b�r�V$�&��jv@A5��ܙ	�z �3�[f{�&��_��	]�г#��yv*��ȃ��w���w!�6P5(�b�$zm�9%�0�3�_��,vh��2���m�zq�\bg�\mj�F_�5�r���#��N^�FVLs��/+���¹1�	��Kmqb�߽s��Ƕ`�9�gð�=������=�뻟N���b�G�n럏�Wr�)���RX�MK����nSj�ۅ�-����]�V=��S(��;���\|dL�s��m(?�ͪQKo��S�tB�-U�$�(�٧o��zR_��ux���5�����6#^��<�N�:�dw�	wQdL,����lu��6e>�yv<���՚@ج[i�oE�9�T�`�ѝr]K�)-�b+k봰b�H{��w8�氌~P^�W5��Jtj��u��#5::|�I���/�FYʤ�4S'�Ö�P�F�"�F6]sn0�Lw����Z�T\h�_]Fa�E���D\C��td�)��!����D7�Z��\M������DƼTq8�|����	Cw�d{UDXX#J^@l�^N���8�/���~5�6�\��P �qhp�;�-Bx�����<�Ͳ���#����.H�W�Kl��,3��[
}R�Ta����=&�~p{&���N�Z�S�i���!k�wl%����hGR�o��p�&�C��'zu��D��`�z�؞�ӯ��I���c@�.(��yD-�U�QO��>�BfwId��&6c�h?���\i��S��˕� �>���y��P�^�VN$�s&P-N��K����ŀ�G8��(��fb��)�_�޻^��X�0�;f��j�����y�2���k���J�\�Y�~	oZ�ߠnq�c�0�^<|~���j����u뮾�MP��Ɍ�6�Ga�!l4�/N2uh�gq�Q�1��ֱ=�`�����u�|�ib����l���Q�h^���9e�v@S��ᶩI�x�"sH�Wʺ�00H�=�,���g{�]�U�}�;}=?5��H{�.�v޵�q�K55�H�Y�\��H���<������S\X�����Jv�Q`KQ��e{H�����P�������"�&lWA��M垳 ���.��KNod�(a7���E���_f,j����d�q��H�Ǡ/e9��`K���e�̄����O��r�H^�z�N���|aB�E׫pV�v���=����M<�ꥳŕ�8�]�t�9Zo�u�-�ǘ�|�c_��.��-�nD�b�=v���+ȸ;�����{���_?�\�W��T,��f��y<�,������ ���J���W8�N	�ݦ)x�l�n��9��w��ƹ�E<4&ڜ)�.�)���xIi#+��+�{b2��a*+J�V��)Q4�W�	��j����uh��`Q#�+��J�J�p{m�����q�blO�ቩ�D��Ǧ����#=<��VS�>TN���Z� meAp'�O�G��E�w��Ӕ[̥S��` �o/mBW�r��Dz�������8蚓yΒʼ��9
���za:�[v	fi�~Ҋ�u|/�8���'���E3ջ��rbuz�#e	�.Iw��Zbw=d%���:�l�U#�(V9��a�H\�M~�y�)����|��a�^��O�����p.��t���dl�a_�kT����b�!:9�h�b\iq4B�r�tr���:�����f�8v�H�mR>�k鵕O1U��8g�f�l��),��������Ƅi�6풬����;�(͌�v���$͔z�1��橞��@}������"�[�;�j�(尯��.��4ǖ�l���v@nx���o�\�F��Z�Z1S�eN9Ɨ���9�/�q:>�t����G��DI��My�V(�q����>�³�Z}Y�D2�K8�~u�X�ɌX�8��),(�Hc�s�Q�%へPSl�a�A/T.�xS�С!��;|ըX��v��0o�6�qQR\C�/O���E�h���R�fzR��YA6QuWR�s�o��I�;��*E@`=-!h{m��_���ػ��#|��Ib�ي])EH�v�jV ���H�&Ȏ�(��.����%���@ 36ׁ��)���o���j{�J�M�V3��H<󯄀f��Y����E���Wv���y�A�uL���_i}��L,o~���=�oj�^h��긛����EhEѦG��V^� 賰!���ৰ����QՌ-�;.�Pc#6��X%�B�2܍���i�ݗ`{��������:-;��%?��\;���^[y�os,6F}�������`�D$���逴��|�J��#7'��z����H��4s�t�atTYpsILg�,J�ô�[�Z▁c�9�⢯�_��m��a�+ӆ_��Ac�%��v�87���Ҽ��D*-Xn�q>�wP�5�@���p8~�*�+���qN�T@8�C+@���>!�䏮�Tyf�.7����{q��y�j����1��./�?e��P��we���:�~��	A2T�D2rEJ���X8#�|��NL\*u,ADΉ1���>��*����?��,��-�K�	���gJo���5���߄ �r7鳙�s6*�ot�iJ�R�;�v�oJ��)p�Y�:&U�$�2]�Pb�y SV�W�Q����]�|ٯ���z�Ҥ�)>]R,��e`�	sm=�Ux�;I��\��+�F!Ѣ��2���.���������ɇ);�Y\��LB0sm���!���y�O]ښPnI9/l\jl���}���� Ͷ��]b?�4uq���v�:�bb?۪�� 7�␉��v����Dm��~�Y��q��9��֕�)RM֨����e����ԿB����.���g�O\g��\�G��H����R��9V��=��P�Ī`Ah���f]�(%L5�C�s�-�����x2�����ϻ���G������%���2�^��C�g���{���IV����a/p���dc�m����/w>[�z��9����8P�ً7�lb�P��<�	�~dwOt*�������3�Vy�.��dr���Q|:m����Bcwqr��D��"?\�"�:�>�i�o��k����%:S�g�`e!�!�p>�|gY+���27�!B��ET�Y;Y���a���	����;�X�jBW�s��e�6f�F�A-h}AJ�a��1R�A6x�����5�.�����k8AI��ա7'(Vr1Eͷ(�羯�r��*�6�Op��}�ߊ�#��@�C6�>��*���3j��-pl�ch�X^�����n\���L�������3D�1J-�[T�Ǣٗ��s�[HV�S��},.��I���#d��F�ƹj�\|�A��tIW�:u��q4wL�����9d�똻�LAe������6���4��K�&�R�|*�{SþL�B@�}�+i�D�dU��!���(�;��X� &�w�w@0`����Ƒ��J���
��z�aǫ�5�}�#%�X�I4��5��_���2n76�?÷ȧ2׸��#�C�Wr'_wt�zjߩ�X,�08 b�
�d��D��_�4@�����r�2�®yQKr9�����I|��ۡ��'0�3� ���Ij>T*[=��T�z�/q��
�K�WV�t�"'���&.F�����Я�U�6�FJژ	���e�B\h�������,��ӗ���Ӕ-J��ôw���YKP�*���*��4TE Ƒ�l���������K̦��ր��WƗ-z��'�&=iG)��� ������0�@��M�Ϟ�{]�؅���Df�'�x���{���UX�D�)�H�؆u<ו����i����a���t�>�0>,{��j��g�>d]��gy����>8?�B��D��tx���S6:~g�'>n,H
m��W{qBR�W�����V$&�T�����q?�8A��I$qxO����pt|�7�7����sϠ��h�_@[�6��otw���!��up�ׄ*uG����*�z��ob��y�򂚕(�F�;K�l_d@4��TJU``ޞ�{^�C=e|)��vZt�T~�h�%�f��<<�;��qf1��#`r��=�Z�K6h8/-�����L��ӈ��B�`H����Z��~T��6�8���醸?VY���s���c���:�9OaE����v~U>�J��`�S1���"B���j`�@�M�7���QB@ �Io�فfɂ"X�3Y\��JVeKJ2*ԈJX9� 1�e{�l��wcn�/蛛wS�>J�o�@!��v�ݿo�=�sQ��~Ci�h��B���2Wn*�c�+6��|�$桄>�t;hz9��b+j�R�"�&cO��#�[����M�!:�35%vS%��R�^h����ha���O��n�&O���
դ��Kr�侇��	)ar.��קio�&4�[d&d��B�Kf9O'�7�c؈�8y��{\#�	(<S���D�D�k!s,8��{�<���kf��9drM�1F�s?�-G.����J�T�|�C�u|�>ќ�KC�-;�3{t������I�I�2/����I��������H �h	'=��k�&��P-��;R���O85�����Ijh	��a!��EH����Ri,'ꡃB���DO8C֕[�p��W�ߧ�{}�RK�*U.�l[�l�iq�-����a�x ΏV����c�_;%y0��"�87˗��M���� ���}������
_��~ �כ��G��@�8�w��o�c��|2-�'��]r-?�+<6Q�)�h����.�;�w��PPQK))(=΍��G�%����dO@���?e&P��A�/B�k&0}x�H���۸t;@8���m��vhВ:C�Dck±>9�|4x*TN-E��Q����ݚ���U�R���	��>�����X��Hhf��WowJ�6 Biu9{��)L��nSG�Լ�tfԣ¨F���� ���@ r����iL�����x�` ���*u>��gF����A��X�7ј(w�4�4�xp����Y���s|-�5D��ʠW_�y����M��!NJ�5�Y&������qЏ�]鰔�kJ��3��`���G�V0f���{���ޱb%W�Q:�dL��q{5������D�G�a<E��8S�;ˀ�U�"�h��C��8Wc~VR�Ԯ�Rf�_4Hp	�.�(բR��S����Ӫ�KlɆ�@��},yo���}3��#W9E0�_�`X�R�/�l͏�K���$�'~s�9����Kվ�蹔��+���S�z��RʙG�v�ŰZ� Œ�u�緪ط�U��2f=X�r�ln�}$j����Ō ��`�&[�.Y����s��i�h�X���%eBЄ�5�1�`|3��a�o�֎����� �I�ި�2�������㠒&�@چi`����r&�����3'�K�~=�.��7�]�#]�'T�é��i���=���{�~��1�Ըg�ҡ'Ϫ�la4Ђk�$.�&����\�����\<E9�.C��߅L���&������xy�m�J�7U�3�G�^��f���YO��:,aD[��F�"JYء���`�sw,�Am����
�j�X��\u��5�'�1UHC�PI��w0d�����ztR|%�=1�P�ѷڐ��iz8���fHh�p��-�y�-�*>�㑴���6��ǡ_����2&����f���`�Zl�<�� �w�m���<bvR��^��g�黯[���ʘ1o��9�J�	�-M�`�[fs97x�\�\�4�\_��*�_`�:^ �UZUŵ�����l-9AԸ!�+sN��j���<���s��춾�s�w�4�_��`��2�<d���m{=B�3��r �0��Q�� �/E-֬�+3zZ=Kc8ʺ&��<��>{����Y�$.�,��/��R�:�g�Pu�!�_�O�/��KQ�U.���I��֮��pXr:>�󞷅!�Ȗ>/��=��n��K��.�F������4��5��4�k-
�@I?ǱD�J#/��]�9]h��b�7@��+1Ш���q����pD2�r`)H,4h��ܪ���;�<�mKvr������;��;�4�c;k�.��獔A�mW�yZi�i�[8�]W>����|�iY
d�K$^��%F�x��5YEi����8�4�36cy�O%�p.V[� Hʟ&�f�8uL��#��Y!�3�3�nf�"4��\p����MR���ʒ��\���,�^nU'�J}�2����?��,�x"_���02�	����Z�Ѐ4�,���UZ�l�?��1�Y�\�
�\|�3�J�i�S�c4� b�/:(�܀�t=
zl��[ݸ��l.*�����|)1gl�m��Q��!zwJ�|ݻ��%�+��~S7�4mP9�e�1�Q��;t�.3��F&vb��|w/����z��zh
����Ean��[r��)����~���ԅ�s| ����E�2�1��BHr@��1���.� �]:Z��,_���=�{��p��>��rFX��;S.�J���9�����i�B2+�r+J� h� ��(Yeڳ��]|�0�Q�;C��m��$8qn� g���k�<]���.gP����sq��0�i���h	�9���7�[^W�������z7�游�Q�R�W��t�&V�62�
�J)E��?}�
XQC��t�P�P���5����=aC�p�7l=�$q�5� ��M�zjGF��wvk�8Gܝ���,�w�Et�	������g�_����~c�e��M�4U��oD�.�#J�->�GݫȌ���o���ן�{����xP;�R�A<M�RN��"�J���Ķ�n�2(6`��1� ���M�S�9���e�2�g<�ap���^�~� <0�w �r&��
����!��8�Q�����ywR��p������u&�=���+�}p����*��e^��Y���  �.-�\jJ�h�|����+����F�;�I���e�c��%�� �;y�,��{L���1����)�b�Ykq���ק���u���ރ��Ke����;(�.��A�B�qZ�X�����i�^׭� Lc����&�����$�`�����Jg1�V�C-X�7g[�Cqx^	aA}Apx�{��idPbv��#G/��ǍUe��QޘW�	P�qӹ��˩^%H���*��M6�!���,���vrY[S���6j���!���]����E�>ݳ��=H�rx}��1M��i)�:�l|��ۉ����<���g����NbzigB�S^Z�3�2�vG8��V�XS�ی~��j��e�C�g^L���x��&ϲ�����$�2)��N�8��7�N� m���B��g���(����φJ�2�ٙc�6�s��d!0���x�[�7��F/��_kN	�r��	�����b|���a�T���1��ɯ�`��E��ʪ_r�X&nW��}�����\��7 ����߼n6;�KD�.j��U���:\�E�1KT䲤��#�;�+�RK��Rܧ�8H7I�c�A�F�J5���QM������5 �C\�E��uu�m>��3|��H��2w��6��1�x�J�@TX�*���`ٻH�!d~fs����hF�����H�^=x�5lv�4�r¾����{��1%�����-���n�"�UF�<�\O�|���ۅ;[T:�,��G�s>����uJ7 	�Бe�n����7�>�o( �r{oé���5y]�	8TAM,UW��*�����\s�N~Zj�р�Z�|����������Ъ��ʮx��84�.�H:K3����Q}m/��
l��׭W:-��RAiXH�=��w���X��!ʝ����9`7	8lO�G�u�.����̇��:@Gu�;(�M�pZZu���w����'a^C���E��lSj��ϡ|���'�'����5f�Z]9̀�_�B�Ƽ�������C�pK\�[c��nes�`E��0�ڸ�;���;����ˏ�X�ȶ���l��e�'5�0J�ׅ3w�3^�	�ܓ@�n�P�lMY�F��X#�L:�@��\���g����`'*��T���@w�B�Ǩ�Iٌ�{�2X"FS�3��w�	4�.�9qN��XQjm���y�����ǡO�A�T��Z�}���*����\��f��	�i���B�.�M�ʠ�v��Ը��ۦ��~زj�e���Z���vC�N�}d>tM�X��B@*Q�:��@�k���ǩfo^Ʒ���6Ӧ�W��r:L��1a�虰Km�zϝ�����w���%_��a���q!9VuM��� 6��j�kEyڲ��q�
�N�#�:h(Ӣ$���r[����n�!)��(�<�7j�EG$L���|]ga?)+��ԗ��J I����xG������Y=����n'jX�_�"���z"�#�Lg/�.Ew�E�Qu���(z�Op�k�{I�sI4���k�E�kn4�ǐ�z
�}�fF���� *%d�޹=�I_��[�v��g� ]���U��ކ�6o0��R�pkX� ��9��Cj(;I&8�����e'��������%hL�v ���P�8���O�����,$䗁x����r�Є����[^A�x���� ����;�:�YDnI�Im�c�Zp�g���)���Z�О���j�qւ\�;��t��_���W����@��_�y�GE�W�m������D5��@�r��G'S�m�~���>e�L�1�A�3��q��w&k��6��q��;U[�{_b���z����D�=W�j��0-Mc:�CPl��"�P�{�RELC���W
�rl�����F_�&D�:XB@���3@��FP�Tj���"R�q7�+Uy�k
�ƅ�+KDjC�z�h߷{)'|r�� �H7^�gkj"����&�4�0��Z�u�/�c�oF"n���R��m�Y-wj�}iT��5�
:�ޞ' Zm�;�E|/λ�l�!)l=I�w)B�{���8�,���5�iud��	J�u$S5%#q<��`{<ߎ�P�I�P(N���V4� ��3#*x�<b��H��KQ�
F�$7�~�w�$�Uj��TKe��V��c#T�N�}	<�u�T���E�ߎ*�ξ�Dhg�YW8�Q�T銼�а�7o{(��s�]{n��P��ۭ�Ģ�\��Ӡu�¾���5��r��d�D^Ȩ��y��ڣI]-2��˖P��f��^���q[=_1%D�f�ѯ:`��Q��ai[gf w��Tx�����#����)���$xq��t/�E.�}�w�vtz�����)�=�O�B=�ˤV�媉l?�CL܋�B=�[!�
��۸����D��W��ь@
YʘWF�ly�f�$�ݜ�ڜ#!���X�m�y�ݮn�fmb����l���7�L�b���[{�]���	�}h�����dw�.Ү�����,��N4,�1��u�p�]��U�UO��H��Xqޠ� �V#|�����#��uaL>��!��,��qX�:k���+�%i�}�3�l��Ԙb>\�C��t�ԧ�35�E���FJ�9��'��J��DFΗX�Vb<d�n�O� �W�IS_Ԕ�l�5s��`�r�$�f�v(� mJM	�/���:&����UԦ1\�}��y0�F�ʋ���DQ��kp�&�M,�E4��TQ�f�6��rd������Ai���jd�;yp���M�:x�-����W�c�X�z���͇���:;��I1�B�Ӧr��֙ǵ��$|�9�J}H�D-����XӘC�J��e�v��!S�	~��!�q�l�uE�Zp������\�h�r���֐�xl��x�L!m����� a�w��ImH��d�-ʹ9Ϫn�V��haŬ�I�_iď9քiff�_P �ތ�%k���
�$�	�pꠝ|�("j��P�\[	1O.GϮ%Y�����i��RbkH���v�m=���;���7R��r�{ƫ&I�m��r��!?�`]Ϭk�s���2B�ٕrpe�����eP���^[L%�]�x=��ޥ��u����}�'/K^)G�����ϻ�W,|���T��P�Үx$/X���Z*�]���Cw~�����`2�*c�'��pFh�%�^g��b+������9�2s�|?ܷ֌T1���yOZ�-�OІ �0�y;�K=9_U�YO�m�̀��248����Ng��M��ja�i����<+X�K5���tƑ�eymXO�)��ՎT�)��v���2�R4�d�:U~���3�w�b�N��7�pY��V�'�����⤴Nr�>���q�Dj}vF��_�&I���/���➎�۩�Gf����|�� T���ޏ��-%=љ"W)p&!4�6�z�{�>"�N7���t�2�x���@/\?�~x�"s+6E��)�_��Mf�M�h�mN�aX<�'�3'���.݋>b�����vȇ�����j�.��AXؠ-�9��HX�0��0�.���;b ����*�y�� �\iN�w-(�C���:�h�*��r�lUf9��/�7&��hf��DbYluuJ�#��]$Wc�!T���8�p��I�ТH�@'�z?��^.��AB �r!�e����9��t�E�>kl�	�m��"K9g�r���U���g����$6F�o��<�J�m֦��[��Pś��x���
8�,v�[g��%4=?a�9�Aq����v�J�h{s��#_��t;E\�����yE�8\f�\QF�9K1��L�:�*C��|J�*j!��	�h��X��W}�n����Q"��gC�L���J�sc'��|��V�ٟ��K�?��=MIo�V&9�T�; l��+ �4{lG���:K���ꭹOƋ���=��_"T�K�D��^H����X���e[�zŋv��0J���2�X�0��
V�*�e����2�&�iHhDOPvwӼV+� mNB=���L�3�v���T���2..e#�E2?�|"޼2��Y�ݱ`ֆk�����-2�j������ <#�B��7�9Y���(�HW���#N�^�p|iݞ��N0޹�b�*��L�R-��ʡ9��;��50���/ڍ�W,v	��ͫ�����8����+��nT�+ ��
��z������＿�5���aqvKު�G��X��7K��S�a�����4�Ȇ�"��|-�4�"͓�4fd�oz�SK�-O�e%���b�P�;u���pF��̀��Q0�d�ĔjN�
�NQJ7JRow�ֽyː�%���.U��O����:޶�n�]�<Y� �C�S0"����r�$8\{#���As|�W�м��I��Zi��m��e7�Y���mN�ų��݃�����ݑW�	�rn(��j��U�;��=���ݭM ��1�(���>~g�Y)ܘ��W+V��Ŏ>˖�ø-�D }������W��7$���n��ƏcC��Ixn�א���Qr� ���Ҋ@���D�$ګ�f���~v3R[M��\��?��w� '� mN:3�Y��*Ȩb�
y]c�n)����B-cA갇d}��?��u�C�n?֯�����Uia�J$�Į�kT�%�ŗ���UM<�#=fh�4O��~m��>�ٙ�G�OGa����� ^�����s�Rs���+ vhn)r�%KO(�۝&o4rH�b*RW}Խ�7T�G`�B����Ϭѕ��)Z�w&�ZE�������t�w�Lr�zc�C1�}X��wFߞT�� 怮$BZ4fk�J��R�����V��-Y��X��"��d��ںZ��=X��m=$���c�Q�>b.�<����5
vX6�~7B��<��a˔�/����<)��F O��].�d��\�Ge�c�E��s�b&E��;~�O�N�'Y�-�"es�H��Rӣ�y��o�o�"0%t�=u�Du�Hv�u`�ȿ�u0�h��#���sZF@�J�ٌ2��FB����b�=�m�O)`�M���F!"�v��W�P�c�XG�'��l�8_~����������4m���,qܪ���@ݾHv�h3����LX�}��)X�1I�����E�0�Fi<�$Ц��K6�n쉉�4;Qp�0��Χ\��j����D�l���U����,í�P~u��-G����M^�Jw�7� 8U�� ��
���p!�@���nE�S���μ�#ֵކ��GH�+kѥA�q�aG~��4K@�f>o��^�d�1d虌���D�{�ʗ"=�}��J=�%K�w!bl������6mX@&9=G\�ӡ;8<�sb%.�b�/�����d�3���8(�z��J�y�)��S��S���FA�>Ku<�gb����!���-ڈ�Z�y�(F
��3�Z�6��l*3�[1��)�y��P�S3H�DB��7X����b����j.�N����w�\�	津xK5���M�t�CXJq�S�Gi��8�y�����g�o�LK ��6��Z���޽����)���G�!}�T�2�Nm�<l���]6�e,<`�0v���r�p	s�1p�����1�6��1�uE��%g��	Mꩍ�ͫ�:B�u�&n�K+
����d�
g/�3�e� -ߥ±��L�t>������R��!Q�D�ϝ�V�Ly�s��A璥H�g n���v~�CѰ��D�]DVϵN��b�NA(x��F�<&*"S��|aaUl"5�2)��� t�
���t�Dɲ�C{�\ym��V�ߋ����U�D�*B{/�y\)k��n�����x�D��0�qϰ���h_�
�<�KA��Jfξ��`�P����?�ݝ٣���0�GX:N<��>z��r��>�k
Y�����͝0{�W�X8t��K�T���LXI�w�r5�E���b}�����Ɣ�n�GM������K�B�ݯ��/A�&�����,��WX@�kVU0KLk)RY)S��i@�G�ݞ�GcM�u�m�c"Q�7b���1�^�ƞ��3��Ml ���C@�^������:��s^��T�e9!Z�#��:.�{N���I�Z����x�3Ɔd0��bF��m߻BBJ/�lx�滢��W����.��� &���s����_�T8�ڇ�d�x�d���8(�&�6*r��L�S�m���#*:��0��nԜ�
�����>��W4����L��7�}U+�2L|�r۽�_�3kWͅ�o���l���`�i6 �p��-EN�o}-�N#Kt}��A���� 6����a�>Na?�T�쟢�۰���ުCZΞ�UgbB�'��2j�`�[�eXE�G����m�>�F&���&F�d3��z��1:�Ox��B���<[1i�����%�h!ܶ���E��Ӛڤ��r}u�oI{��y���u�05x)��!JcϘ�����C ���W���h�� �^���%(��F���egq��S���-/�ƚIEL4������VB���h���в�(.l_��z���	�<i˧o}<��,�u8����ue�w�[1ŝ�$����>���wER%`���㹠q�d��w�9=C�-�陠=�,�T�&���Alc;g��w K���#��l��n!��N�DgM�m��q�p��φ�㤗�)����0�O����p9\�]=�x��4?&pF�8-���X�_�0j뚄��A)~��J�ɐD#��,=g�6���6M_20mm�|�5�H{�~�̂�����ƏQaw?��~�W�����]$�*@9���5.^��[��Qn��Yh �\:y9����t(�@�-k��ј��ԍ�8���AFmR����>����t�H߭P��ҭ�V�e�uQ���`�@*U7�WPBl� �sGxXM}�)���2�f:���m��w�T�y{�0P[�9�f����,ؑ9��
52'N]���rwA��\��wl�����o�dZ,�3�jI;�+1D�����-ye��VdW7���������ݻ#=���S� e��I�S���x�y?)�}��E�u��M�i�IC��gxG�F����,�f!כsJ�Q�V���rf_υæ�S�.�>G�?�V��ि{<m��-�"�x�)��҅�)kLNc:�lJ7�h�o���S[U#�ŕs�hi�'9��V]]�T!���)�Q�*�M�2Oϟ�y,4`�^ūS�ǩ1{��o�r�T�������3 k�7�j���}jV;��U��Oi���0�vX2Y�6 R������-N,
�
�F_Mȴn^4,ְI�`Pt�j%.��~G��gW��w���
B��{�[�b�ͧ�mv�����~�$����$Ś柹��(v�$>�c��pjeZ^�V�]�a�����*�L$7@�z�N����u>�b�h���	ڬ�E��{��ԽH2P��P�q=�+PD���@w�~�Zٕ�Eך�w�bM�v�r�fC�w9�M`��>����R���&G��M"t-����x��P/l�I��2��!`��U.� z�|��fg�WX\�0���#w���r*Õ$R;|����䧆Ն�8Ba��U����lՋG$��%1�-2w���������B;�?�1&G}%��M%z���rr�Ե1*ׁ�	�'�s�@�P�K2��ݜh��!Â(�)��	1��c^[��I�>e�R����A��KO�u�/� �iE��<Xq��Fػ\���lw�q�X�u�^�p�LT9�R�Vw�Ї��Y�іc@�v"�jK�`�qbfd�|\��Jγ����܏�J�(��H���ov�M��(qB[����v�`?�?�&�OS5�(\	z��?��^��!"��L#��	���V=�(x�-���x/��U�i=���Hhg�?5���3�|�����6����0����3bw'�]d3�˼�}R��L8
ܫZW���\��h�`��:I�~���3�G�f�1����7ρv-��.����e�0��j�ȡZJ�h�KK��H�gvĝp�Ћ���D��<�ФD�B�ۈJ�[��`�ڿF��^�,��\]�T�'Z�}����~�LQ�C�f������_��ޑ#V�@��0�:i1h���YV�B��ܗ� ��<�Hs����)�a̼��D/T)חWE(�Z2	+�G�	C���ٳ�f:��j���sR��X@!�͖�F���Ы
�9\̹���}���_�;�%	�67�J����l�~q[E]���݌��/�E�eB�Z�������'����|�:�E�'����Fݝ��]���\��O�!D��6m��mn�T2�r�8P��(�o
+|�I-�tW��6,�$7\J����˵��� ��U�ՏA "lB��MR'"'�!Z�Ͼ\��@~��y2�$�Q�M���i����!�S8W�����Ѩ�
�a$#՝y|��R�V�Xq}l���D��"Ѩ��kʨ'�'#���;�~jr����N��D����G�����~(���e�eK\,쌁���1r� VUq��W"���hoD�P�+��K䤽|b���&��Ob@��)��?�����w�|S����o40���2Ńı��PBk���qᙎ˖���+���>Ճz�/)�����=H�T�<��7[V�@�u�"j<�o�RT�,a�{��� �����2=
xU����y��
��wO�Z�=��k�6�����	S������1�|Fq2 L����ޡ������8Q�9�����a���m�|`J�X/�P/���g���yF*e��Sb�8hiH��`y�7��f����Zn���]1����E�}��O��F���_B��&�6�yV���7�D���GF�G���-��"=9�[�sŀ��>����hC���x��Ő��Ue�����Ŧ~DW	N�3/o��̥�4J�n���:\�ق������{�	�An��m�����
�Ti�2�� S6�v-P�v"�F
�}#k��]tm��-���0�k���dp��_ɦ�t�˗�պJ�.`��qO�i��&�`^��/�'�T��jj��oR[⡁0a��*}U�\/)��F˶�=v8�cV�6�d��'�b�&�@$jm�M�G9Т�t��v����]��d�_���qi�{�;Cꀵ�± �	^D���W����'��ڃ��VGHg�HP�E�,NVߑ��P �ː�����Ĳ�f��0�UFB��mU���f��G��$B@]���H�	���9ѠM�##^H*)H2 �P)����G� �P��&�P]:�2ɱ4Z�P�d<���k�Jg�/>��SV@��� �Ց�X�hlG��m�m��	i��խ|�e�Z��2<��T�Q�G�q`�0J�/#���	v�x}��׆����&�X��ſIl �c�gQ�~*`�̸eIPjh��J���Yw�����G�E7e�2�-�m�u!p�?�}�N;ջ��px((�����*,��EZc4�0�f�/�)�V[���<�f����pnj��߀A��ɒ���yN�b�,�Wp[y$^�V9��%�|�1��=0ϝ[��*y���魶���{0�!��u��h�O�aIŴ�]I�Іv�{�3I�M��i��Ԫb}� !ݤЗ'3,Z�^¡;���?ϭ}���VѢ�����d���ο����w̹Q�kS����_��~��lbEd�bOAa]M�zV��>o]=p�	�Ȋ�H󴡅\�����ؓi8M�����T^.�[6l��U�x�Z~�anAiOt�>���K�,��Nlg2.����N�F�mP���o���r(��I!�sX�`d�a��H};]�}�k�?<Yį=�P{����"B�]">5����L�K�~g�0��w~D;�`��&�3�7' Z\�Ֆ,|����Q��M���1܀��8�"ЫB5λ���y��Ӡ���c5}�b��l�����b�u��LML�xrv�B2줾�����X�08g��̮bEC0�!�i��r�q�`w��#0���jb�-��sɹ��8ȏ!��@���ê}��(v��]�{2Г���7C�p3 8�
�M�]f�Շ�����Nck`h��Q�h�gDa'��N_�	�5$��3���#_������lV�1�N��#4� �a�	o�7�f"�N��mOnqA�^�x��� �ٍ5V�zBPh���A�2�7� l�MJ��4a�Q�z���r��P�������.X�5=��2t��N�<��	ܨ�e�Z�M����2�&�׾)=?��k�4E�P�ʊN�	��o�T!���:��x�M&:V2ג�3�92dڛft�8-��i��O[����k�h�w]�I�p�g��W+.���>�lLh����X����h����K�E��w���"\'��?�� �X"8l`.%�]5eѐ�AJ�Y�4B���K��־��<��i�f���
|��9:���m�%���=�^�Y6N�銂)����R�<R�F7�Z���_��:�FSf!��S�{��3l��@N*$&���]6��}�Y�zN[�9}1�[FA��]���3�
�JZ-uV�0��P�=��}�g���7��h=og�޴�O��y�
k/6bm$׭F����ܒ0n�r�������Ud�)���zD��� ~�Gg�{��]� A��<-|ˉ[�^�?rQv�/0�3�`�;��}@k����=
���,��%!]@[W��6�
�񌏜K���W_�.#8�����r��I�G}p����tS1�� ?�]�vy;�F�1�ch�4�Zz�u���b�;�	%��g��l��@R_�J���3��'&~�,�Qk���c�^ �67[a��g���G����+-˓�ߦ$v�q8嬽��%�b�]\�^j�X>,�����ӎۃ�@X�a;�PMZ��� F��޶ ����yKlU�מ�Ҁm��IߪT2���l�ڌm���Rg.l/��Z�Rߍ��a[��)G�XQP/��BZ��=�@��ih�3e�9q����f~����7^��8�^=�2��x���D�A����%ד�������`I�pa/ʳ��;>��焆C��9H� }v�Hy��O>�2����O�O����A�DB�%�f3��J�E N?��$#m�Eaͮ�yؑ-H��8�� ��2S(V�u�3gҲ_cM�5'#+�e[Q�e�&��u�v�}�d�kp��'��qA��t���EC���~G� �#7U���A]�����QN���u��Ѻ%>�=-q6C�[(�V>���LIy�:�QMV�S�G��J��$G�5�}b>�|�������l�Mf{�byu;�W�A�5:��I�8��tNEwm�.��OKn4p�#��g�^vF@�wIMǊִTr�v����jq�Qx����ٵ�ebfB�O�=�������h��z�"Ym�?���d�Sɬp����O���X�U�(��C.�>��ւS���?ŒG�������(�K�m��,��D��C��T��z���q&�@.&��M����[;��Dy[����.��3@d�y��'����US�6+����"�H���$/B�ax�IT�ݸ�^��B�y-3���A������Ӛxp�����:��7]��J����0�,���HCt�lJ>jK +D����p�W��|�%��?t�&��&�D9w���8��L�:>e��Hʩ� PYh��`�x4�Pq̨���\k�!{�e"O��D}UFQ�z�'a��*��lJ2a%�k��K��f�����چD�����J/}-�kD�u=tt�q���0�w9��Ӣ+놌#�K3���N{uCj8Ex�  ����CΝڒ-���x�]ۙ �a�B�0KS0����Pi�,�v:r����x_?irH
!�X'!�9�.١�Q�M~�Ҡ=�F��6�ٍ�7�P����y3�;b�g9�Zh�v���㺽���0I&(5g�/ �<v����y��rl�Xv�Z�0�%���s����|��-���m�L��Df��M���=g�~��ǲ��1��%���%� 
�Z�g�&~�����e$q�q��@6D�+�J�+��;��T��&8�
��S|�?�-�p�_�L����]�>�6���Qq:�Xy�[��>��\��,p�I�!�Uy��h�T�ҵ�m2�3�{<�7^^�v7KdS�{�#N<:	x;b��v����y���
w@F�0}��W!]��(;��_�0Mo3'���CQ�b�zԹC�4s�D���:�� x��OE�c�W���CИw�"�"\D[*��-3���������:��xχN���ڢ\/�1y��Cq���rߧf����EE?�%��Ҭ���]��	jʰ���s��8��_�)3w���#*t>�)/j*+�"��[[1{��|���
�ە��[�U<dcO�Hv��C��w6툍�hN�7�9�XX�o��c��~���S��X"}�b�<�� b�����~,��Q"҂���C���U���Ƞ��ѫw��.��D�K_+Vg/�kgƏ��zX�\;�������e\��"B�Q�t���T��e�*=r�Y�K�%��6�����ܮ�y<NV�$�Y���S1bϔՠXl�����0�2b��Y:���j�
�O�W:���D��B�� 5g��,���Y�6�ֆ���k�'B��RI�B��j�+���m�۾�bNª�D�&�C������3�#t�M�%�\�������K��v�3�T�����'�D,�r�*����8P���� �Tԃ�޶����^^n���b.:�G�h&Q��oIh[����c��B��SQz�̺����
k�9VL��\�4�x��ݗ�2�ت�?��p��3���cj�XA�ܧo|��+�"�?�r{�/9�G�	qt�����F�f�^�Q��d�0��o!��Q􌾑$�bw�6u��}���s�z�Ӷ'JK��ǥh��$]X�T������d����g����33'��z\�Djz�X��ݛm����/тu[�L[�Lf)��;IV������k:�@�OxK������U��x�8�T�9"�X=k�F����|E�#M}I�vM�}p$t���w�r�ުK,�2���4��g�܁r !�(��ϯ�����`c:�,V�!�:C�e,#5�dt���S>�@���O�r	턻J��M�`�,��_bz��iK�̥�*���ڞ�"���OF�ԫ_��z�8���-�O��i�y�U�[�����G�X��H9���J[��8�fM����"�b�%�gƥY:N- ���
J�_�6�������EZ���S�'��@�I'B��J�u`z�d>/�80n�s�V�F�O�x��=`s��t��-�kէ�¼���z����u7M� mfu �'��A�Tk:�b��������`ˆ˼]��FbU�E��=y��C�2��a�~1`3j'.���7��\��Ȁ]�4iėX����%O����HfE� ��[��u
��J#���F����~��L/�;���m�ɠ;�^\�Z+������pJ BL�}8��g������I:�h�|�%l0��;\n�]�;S��7&�(�q��8��-��b�e&�,��ݡm��x�W6��\�҃2�
:�3K�b��ԍ����F�{��&˧?��f7��6�J��!���H���WR��y͂��Ҧ�Al���u��v�Y�rY���l��a�J�ʰ�誚^��𠐖*�����q!�[�"C�~�X+�ae�;NjX(�x��e�!����O� ��;��|����_h�-�S-E_?q,�>x���k fm{��9��Ljk�+ވk�)V��m���x&���p���l*�r�<��t-����T:�����{{;�i*�S;aU�w��.����[���òj��+]�x�Ϥ̓q�X�Ơ�%"tiz�{����ju����ϟ!��r��/ێ���DC�#�����gz7��(5ZkB0���vP�h�A�L��s�TL����';��?�z����A�P@w����v�Ny#p���$�������nC�-�
d�'X\�M[�m�BOX|�H��� =�d!� @�����s�'�0'�X��׺?�Q�Z�\P���.���.���t�
A�0cV��b͘��p$sk`)��V����(�{�/����ڻ+��jr�޽&��� @�ZJ�e��٧��w�䅵��g� ��LF��B7Y�F�&�1(�_UK��߷�����%qs!@|���d�g%���pX(�����l�y"ѧ�i��
��IJ��)YO-;hИ/=M8x7��*{��8D�+���+�5k��n�.�T��X�7�m���Ο�$���Ӹ��:ߴ���{6�l��^�%~|1�}ӟu�	�kB��$��c��lv��g���H��C}+n#vl�RS0� 	{��F=Xѝ.f	�9��BԱq��V�����3�o6�����4,����޽�1�AO��� i�6�˳�'�t��nv�^��=l�+��%e"λQw_zfT�
,] ��oR��~�=�Y�{L��Ϲ�>|N�5s���U�>��R���@���b�	t�	�lgB�?g�n�8$���Y�I���c7~I��Va����߶s`K�{'�b�������_��$��$?�Wxl����GV�Q�\���ߋ\xz���:ВG]D�3{؎穪���U:�R������0P�f���9<�#���1
��N(�Uߩ�Z��f]il�[:��i�A��$�)�Z�Y����V�cһ7u瑨٘��Ɔ���E��(/E��rs2����cQ��ç��9ȓ�SE}/�=��>�ڣ�ϙ��O�_���m�'��T��5����1���CVm'�X�$�J��8n�3�������	+���_q�$�9�)�c����$6����<��Կ&�T� ���XB����@�fuq�����ջYEn�VQ�����!����'$MՈ�
����E9-twIv�E�ް54�~��H�V'��XMI�n0�O<��l|�SRfD����$��ˌ�Q�{��3���"�9eeG]L�H2ܭ�J8�TO�l,��
���s�I�� �X�Yжz������|�AD��!����2�oO�=UW��Eu(�fv��O���y��<Ӧ�V�V�s��ۧ��z*ެʛ[c�M��p��Uf)yq�����w�5�����9@|Ǵ!߻��tNR�x�iMY�<�Qu����J�C�ɸ)� �aoUJ���,�Qx�$����&�� ����ح1�Tt�zڜ��ߛU��ݔ�Z<LK�u$�ѱT`\v雫�1(���(� %k�,�{%Q����>���=D�����}}�Tݺ��䪵�r&wk���5����F,�h�j��@Ņ;��yPq��ݪ�V�������\M��AhE�[���$��B�/z9�1߭deβ��Ϋ���� r|���^��#nT`���\Z��#�+1����,���UG%�y*.�d�7&�0x*��cF��s`.c����#��xȕ�	�9�8q���o�����d�m5&��'1������py��(q��=���m�`����><����PIX����;=�#��+%��n�d��D�B0��'V��hA��ɛ�-���H����T��}&�i��!J���J�
�X�P?�:Y�5��*C���	�3I�3�V6�ۼp�Õ���+�Ȃ9������A�P�b��A5�U�p ��CΚ�;o��&�S�d��Ɏ�:���x��KO���2�V��$�&�z�?���f�6�@��e@E��!XvFr��Tϧ�{���fA��HH���b���Jt�D闎���E�F����)U�W��@�<�����ÿ��ՖCSN�#{�H�}��!�����Z��@14�4�_z?Ɵ���r��c��X]�W����v-.�C`����I�!)2�\�w<iF3x1���*�;Qh���2��Q�(������1E��8�6O�����$�Ś���#�FR�����Ev��m��	�buf�B�N����%F��~�&�����-s��e����t��Z�N�>��%����֫��ߙ���3�Y5�2�������8ɢ0��yۀ��'N�gפ�[���D�����O�B�<����FV�9�u�P��C�GG�mA�8r�D�0ڽ��{�y�}`3�7�طy��9��N�.m7����9��� Sc��f�uW�N2����G��#��)c{�.����=R'K|��3-��+���{T��H�}gm���q�(��ݫCd���p���iF���*���L�ߠ��R���H%��N�S��� Ȫ�%�N� ���=X<^�oӤo�昸��0rAP_^mjw���Aݙ�@���7�[[-�V������r{�O�*4Dj�DȱѪ�v���l� 0Q}x��4���&���͡�%�N��e�J�2���vp�;���pܾ���D)A$k���T.V�J���7�2PU��)�8�'Oh��NR��B
���4�p��0���\yo�F<jy|!@����b1�^�(�� 1t�T���X_��4l��|h���˚����Wh�U߃l"�*4���7�檘6 QJK��]R��|_���J�Έ]`�������̍,����&9�L��.C�,\[�|�l##�o����*���#�X��ϫ	��t��`��\��i����;�q4i���J��x�e\ˢW���C�`5F/o��D1���7s�EhPG�B��u�l�8�D�s�����V �H���L�<{��%J,�E�4����]5s�A���Q���Gd�+ҋ<5�������O��۩����%������C�S���A����4�\�!⌍���=��9rA����*x�B8�>�hK�'b�`Ka���ŀE�����[r���T��<��T�qD�Ι�_`�J)���|u��5;?M]Wu!�u�zgp���kĴ?��]�:�v1ud"U���&Q�=�A9��R�z�]Q��x�R#�|J�y��1ë��l�����a��%�Ydh�	����j�BB>Ud/~]Z,�O�_^F�8���u(�vla�.�j�8�l����5ͻ�3&�b�~l��l��.���~��Q�;���/M��cJ�4���泏p"skw�#c�ϥPå�E^m�	d_?�ɳ���y~@^d��(y�,H�������R�:c���g_�NJ�{��r��F�D��~�B��##}L�tLv����F[x�1�=B���I�HY�y���D���pTFok���o�iu�lP�)0o��K*?Ka��8l���c�p�ԚK��R9���#Ј��:�<�J��2�?�j���K��#�.9��,d��5��_��.�&�P��e�a\��qd!=C���B���cI+J�����b�����#{�6�`����@Y}U n�C/	ji�p��:E�^�]�����v'ؓ��
�z7f�֐P��w�l-�A�V��h��Y��R��2L�e�z{E`�{����)�d���x4�?j���1v6L}��T���F*م7�\�kH�bF��[�����
`�֔�c���f�0pZ���-�~z���(lm��ڒ팛G�JLF����*��/�z_;���φ�D��0g���6u)L��/��2��P�����_ g��p�r_m�h>�wj�E�։��}���;1�)sv�,W;�(	�A���Q-�<��Lq�ѫ^�Z�Հ
֭�g��*s(�/�= ;�܃�!�`��M�uo1~�h�|��=ȹ��9�P�c�xV���|jN�oO�򄱻>�1���P�"D=޹�"�>��_U����S�kr��=�u��
 %MΛɰ-ob[B�Z�b�U�R��I���FN���x���`�%Sy�~3^�~���Cx�8(@����N�)X9,5}R�s���b�-�%��x�����R�]��rkeG�H3��S����)QU7%�4��j�
�>׸ԗ�]K�)h�������cZQu�'4]�v֜]�dH��a�To�lp�c,{���Fe��.�x>CR�s
i3�jݿ����ظ�����N		��ϺTFUXK5����Δ�=���ݮ��&��_��	:9�TK�}��T�8����DS�5�\���oO�L*��n�3�QójE�^���Y]��;?B]�ɿP��IL�?��9T�S��Tͨ��x�g_�]���-���P������\Y��J��A.���6$�y��n��ᘟk�h�ry�B�9:1k�l�a	��i���D=��'�z�} �^���5����+��MW>|����p�:�B,i�E	�UG�k�S=�����!U��~��"Dk��8�w�K	�d��-���>�0�����(I��Ml�p��6؝0U���`�7�R��5����A]I�kJ'���Wc�ci6q����Ja��(���Ie1��0nI��z��|ֳ���Eh� �tRT8淪�A�|+!��/LI6�U)������ʦB�{��s<"��4�0�������qӜ֞��g�K�U�Op�QϺ�5�B�W��n��nOp�j�0G�} iR4{��}jwLxڸ�����1�\�f������:{���B��Ixi�+�jC��G~n�1�t�7ܞ�=����Z��qZƖ(�����e���z�����3r#;��lL�����l���w�|ݡ��tL��Ӊʯ��3�_���s���r+}Co�R�T�CrM���b��w1�"�+7��'��Z؁<Rf�q.@���%JR7�숁��\
�V��G�4��MO��r
��哝�'��E�Kph�k�E�70K�½d��eY���[��&P�c�Z�\#�����y�q@[=����@r�<����n��i�l��6����ˤ1>�O�i��f��~�Z#������_���ڑ+���Lؒ���]��0K�Q�0V�E�2W�~[�+"�C�Z����YY���7���
�?ƶ]b�pB�Z����5���3�9���/$�F6�cB��*�	��4Om�w�y��Z���Ӣ�X�Jb.�oP|��\�/h�������}v�*dCrؚ���qI�x��ԈA{	��_�-���0yk��i���dr����2���bn+�;E��ߡx��z��u�]��-0�Ny`7�(.1"�����Khm��S�Չ*�E��3��xk����=_
�vQR�����FMj2�Y��F�Dc��񑈻ɺ�U�H>��8�7�/4�G5�6�V��<��JvL���gKB4vya Ue|-�%Rg>���r@,�fv-��pB��k����c���MN��rT�`����Ͱ��[k��*�k�TRpp��q�X��J������[0�������Q�$��[��L�Spr6���=��*K�SLF|Xn�Bm���S��������j�E�E V���W��V�!���l!�gxI�__�_�]�7[��b��S��*���1�u±���p�H��y)�B�4Û�.|�̢p���q�8Y�[�CM���F�����OƷs�${����*����p|���1�\�~X���xI�|ݗ�� Q�S��	�(v��8����7Jz�ӗ}$�)��,�����[���2�zi�`{uf��1���'��I?p��k��?Fa�(D�1����?�9e�{�A�Y�r�L�bNU�SrڈX8��F㈀@��k���f.~,C�b�93byva�����ʯ���ƥ�r���ѡ�s,i?-ȼ�?Mˬ;"��n�E��Q+��n�泾����xj�#$nН=�������mz����AZ����D\�z�m�l��S`��a�D��
'|����W�� �4�������縉r��H,����I�Is�{��e$���;�/�������H?P>�� �]���ʨ�A�_��`` ρ^�չ�
�j���亼�����}�0�s�% �&*������O�
������ N��� ��x�G��R���%b]WN2BB�?�V�=��Y�]Cϱ��oJ�Jzo���4��!�x��쵬)�;V��Y�fw��y�c���Qj��j���8���3�Z�x�\WY�9�0��y���Jc@Ζ�A�-L���$X���յU�x}�Zy�w����!�����R���f��*����۝Rr<���H�!O2To	�ʬ��x\�/ش��/��K�-��2��e�'�q�R�� G�WAg���N�|���쎂L!��G����$��d�M�����;���b%�����}��b��/Dٽ�y�f$�y�M�@&�w���f~�yԣp���=fE;$f 0���*����걣����|,�B#�K+ʎ2NP���qڎm�er5�dӧ6���"�]R~�)�-P ��^K��qwf*���>��<��A6U�v1�9�a������A���ӸV���N�q�����#$�M�
')�~�t3M��0k�LN�U'E�%���G�Ѯp �H~�f��\'%	47�]lF�~�� ��xV�و�� 涘W�:Ǧ�~�^~_��8��?���~�#vw2a��*/��e��]||�0,�nԁ��R1b"�U�m-�Q�gIt�mcL��t��s��v�F�~��B�}�DR�#���#`=Ͷ�KB�n��|@j*
	j�$^��n�W��̡�������Ł~l���	�TYUGą*^܉{�5�T��8�m!i����N��U%>a3~!cVw����@����1�#�3
�C��r~;�pg?��y6ր^8��e�-�t��Ӫ�\��`�4��xVj Fz��܎��jc�W�eKǒ�G#��3{�r��롬�D��s\�-���WZ��]I�՗�����[ ?Y 8��v������
��g8@��R��/�X%OT8�����l}_�nͫ���|�wPNn�F7g���$��-���z�������ƍ��"��-!��f�>Y+�C�/���U���Kr�b[sÝ2�]�4��^^�q�Fl�I���]�~�]��������V��l姘�YT��#.:�]�6h����ris���f;]����]OZ]��w7�[�M����=��m�78�n,�h��@���ێ��io���2o'�%�̂EfIǤ�B����E�H!�/���L�ѐ�=���q�*�;�uZj�LD�F�%���2�Ԋ'^��"��ߟFXw\P��A:D}:�S�N�Pjs�5�e��k���/T	�w��1�/��f�-�`�yM��n;0��Z�����:�6Y��H�٩��d	������缎�'}aWP/C ��f-w��g(�K��O��L8�
ҡ��y�v�+1�2Gd b_�KJ���|�T���k眩��1'��H� KPo���h�,�E<�S����W��Վ�!�ɔ��E2
����&=#Y??���{L���SGE�n�0L1�8Yv��?la�o|��O�-~H/1J�.���R~C�ۉ�� ��V�E00��t��*�����~����~`p�Z�� 5�W���6�*����K/1C�I �����Q+�B-��bt�/��s�q�'�N��~��q_��l��z�"��V<�a�����ލG���?t1�[��(�9�o 4�"}o��=�xQ:}�����wܱq ����+��G��!��.���Ô�X��&�E���U�J��Rt�?�[�9�P���Q�F��Sy�ʡ��Ŏ�@&?�!9(�7�,t�d}B�.أ����s��d&��X{�����-���E �?Q�w!k����Rk���E�!E��|׎���^��u��t�� (��jv�02�_[t+ۿ��8P����JKV����z���Ǧ ����D���D�8Z�8S����f����J�����E<��M������A�ڃz�e�I0��Y����y����4��̧�R�RL[��95� ��cr�;��R��nx:����$/	�۷T_�/�B/��^?Q)+-z�s�c���v���W�   -S���gnO��'/:��J,��n"�jRH^�J��� ,�W�a�a������D\7ӂwdKN+TP�چ���~O%sfdP\�x+�[t3F普T8��ha|��� �\�{Î��o�o�S#រ����YM�)��ސ�Xj������}ë����Oi�a0��fsnVX���U��[)G�7�φ����z��E`g�L+S��ND]G����/���]�Q{�*�f�u��t)�"�pFT��$@��1����Jwhh���<ʈ�cVl��^�5pA@,�z#%{P7���$��V��2ߛ,�}#�w� �;ej�l< '{�k]����T�W�����������,,A�-$�df�)���DD�;�V���_�̅u�.�����W_��T#�,H��^��� ����I��@���K�Q�)馽tV���M��E��ً�b��>�#7������1�Ï9�7}6M�_��:��|��t؃ mT0�븓y��AW��qf"�nΗ@�"Yh��ZT���q��ۭ�˪�G�w�ѧ:�QH��S�5Wɽv��e��,t��7���p-&��^�07+a,D3%���ҡ����OF'��uZ�+�p��*�Q�yGp)��	�`�2+jM�?=|U��H7���i0q�ЇAW~4~�z�.jth�*�h�t�T�5Z����<T�F	`�h�egf\�L�(S�^�C�ݐ@{c���z ڂ�mޱ�^B��3V�ќ���� �*E�59w����������Gb֦��(������%~�<��{Nրkϫ�sm�����+�j�ŗk��NE`����	4��Ok�w
#��P=�p�.�+h�b���3��>�2�d���)B�����K�jq@k�J�Ń;�U��g"s���p�6$E�˓���� ��z���iy��'����4��r��1�W\����!��1:��s�^��$C>J��3 3����;�(qN�D0h(syf�ꗐ��T]�@t���h�u���`Y�Kd��6g�H D{��Y���G����aY�#�qDC�$Ư�GV\�����P#������)�8y� ��p��a��K�����a�ޣ3�q� �g����)� �if�����U��W��4�u�~�G��A*XR�:�\���}���2� <���S��kN��a��LCqkN}�#gE�}_m��<ʉy�%?�������2�>��۲T��d׼q������%[�[t<w4�ԂE�pb�nO�?L�M��
DMzs�7&\F�t�*�hCP�U�t�!���E���f�<�2��D3i�(�7�GW�����v%��`=��"6%4��~���B���ݕ�Oy���>6T�,��͚R>��˨��+;�A(̮KxZ�J�R�F�{}U-��6�N�"��y�X*$�<D�S]�W=8��Ex!ĤEs��']��ͼQ��JJ�O�LR#�մJϔ�=j��eD���5Y��1�K&�:��2�RG=푙�)ʌV�W�=!y!v��z��.�T!���F�֖L$ʹ�@j����fst�y~$5�MnIõl���~��_�9.^�us6��/�k���kəY���̂�	aN�L�B�K�=�g�.�¥����[d�H�B�;�����/��Q�0�]�}�k�Wy��� �ǃ��cRd_���(�����E��	W��	q��VQjil�:���@mh��z+_��Et��lαgˌ�`��0�Ɂ���J�#Q����@��^��ȼ�)����X�e?��\6�<��Yg$� /��X�8�&qМ\E�Pp����cla���PM�E� �۴��6�C
����dd*��_�pʺôSJ7��15*��	<S!�F4�|�d�q��{��BVHL�� �3Eo�/�L���;�@�W�O�.ܘo6�(i���wi@G��b���;	h޾�<�t�QG�����/����S,0$�s/��s ǩ����1��"�����=.= �;?���ы��ѫ�a���� �C��9
=3����=���+���-y�6�\VG��Eh�oM�"[ç��+���R�q�ˬ�|0q[�V�ԅP�Sܩ�4A��Z������Mu�\�X�?�d�����opF��.ҶJP]�.4��(��z.�h =�ǀ�}olslk�ì�(�Y���)ZS3��x��?�v�!�}������Y�DH�3I6t/�0B��l�ø
ײίHb|�pS+6�"�o>+x�v�6��؊����Ýb747���e��~�@�:1ֿtW�БK*"��$tЯ?������i�����:���Eo�B�Hb�`3�mQ�*�#�X��,fk�H��`�*�Qb;W�Q�y��� ��hMQ���lwF�R(pͳ�f���Ȉ3���@?߲ 2ղ"��so�i�2�S�*�ݸ�d@:�(�?k�b&�����2c)���]Y�R+��tK��`��a�I�<P]~w�qXK��j��`S�]�Y8����:���ISm&TRz{����@e��vU
�D��OhF�l����wwAǫ����\���<��S�m�}v�1Re����L����W'ϻ���y�.a�<���CYT���E�������\�����9�M���6�x��R7\%*(����uPy���E�tçzlO��=�挴�3e0�Ow��;�4��MY2�$�}[��+���q��O,�и�U�)����lT�lǫ�+P?γq[0��0��j�=������;j �֍俓��	M8���Iz+��he+��V�)�N���0�W����"��=��d����nn������.3,|�2��m�E��Yt��h����KLy�߉ެtʼ��l�|�o�~�}V'��m���]?���r�.���k�b~r(��a�O���>2bw,L�x�h4������;)I}�Ɍt���2 �",c]?p�?�d�O�(@|����N<J�^DE���	���3CY=��o��q�k1�?��&�-�;��2�vDDVqBwK%���Jb\�|�� c�K��^pL�!�8�*J�_`��Eԙi*��?4��RxIyB�
B#���zCp��f��7 B���ϔt)<�z��>;N�'�G�⍍����.?�U�v� ��ܪ�.�.-�e^�Y�beH�g����t���L�iO|^���T�nx+J*E�to]�@L=�����:j��/u���P�FT]��u����,�1᱇�X/�������;��J僕�),�w�Y��JDi�(j=�d�p��V�1����Å(�>�m��ԢL�	�@"X[k4����*ˎ�x� { ���^�y֡ݍ�L�Z?4��c��չ�r
nh��u��c5Z�-��[7-eW;ד �1�t�5���0 �8�=H��q��oP�vy�0���;��S��,&Bѵ��f����+*dVZh����ަ�gl�*��V���B�e͋�g�Akg��Y�z�ӄ�3�W�� �P@y7�9� f&/a<m5Q�������K1�v�bsK�-��O��35��L��s��ܜ�w�E~¦�Ja+�z'��䓑���C$���&g�0{�d�d�`n�i��E��`7G#�nxjx��6l����\W����ik�~��`7�Bg��2�UH�y�|�9�g ��v�st0�jb���B�,�o��&�}���y��U6R���	uh6�c��o6��5`5�,�^�c'ZD�}�bBqYC���U���xX�Z�Å↞�s�q���8j7��4��EPלR�5��L��
/�8h��!��'�mp�7nN��������Eɹ��0g�J45��}�`~]��q��n�Jv}4��/�T�����x��-�'�Xx�t�Y�ۢT��U�̹t�DD����	'c���n� ��=��_ά%�w�����?�G����_v؊�%�^�$��zH�IL�~{蕢F�;g�i�WGg׶ab�|r4�I1�q�;�ȨG���S�Y��29���O�Tn���T:�8�k�ZÛ^���O*�a��dF�k�9�o��:Ҿ��o�c��x��a�6���`�1X�i�M*�-��6��Ry���s�ds���G�����6F��<4�e��`ɞʟ"���,'��Pԕ�.���#<������Q]���f�$���O?Ο��]/r#\��b+������=�gtFYb������kvu�7Ց�� ���[Vn�r��63%�譍.�'�[��A����e�K;�����\_E:p�4�7���ϲ���+F�ַb�ְ�~��p�C`3� x���[���j�����M��zGr�N։V��e�t��L~Ï6ӎ��Wm$��َ&���{&�	�E��0��e&�s��E���\����4�$8�ǘq��A6�l4�&fpn�
�����O"��^J��i��h����F�l��
Hh�!��lM��m��U7��5�����1��p�{?@@�$�4�����Z<�Eq���~�f�|�Y ��=`ݙ?��gJ�EP���U_�Y8n� ��u 9zS�_W��\��qwλ��9�"�3J[O�亡"K�P�=��V'�M�?N��v�O&=C�9k�V6C�����K��&GM���"�f ��s?�tj�`:�Bg"ˊ�S����L#�ю��\`��/�Μ�MS:�W�?f�m�M�9�x�P�zz�+��Ԯ�@D�e�gxЅ6���}	q\1_�t묔���Sar�[yS�;�4����۞�S�%ιVl��;���-�!"�e��"�Դ` w��<K����&)W��+�|�Ps���l�M��8b-Y�W����"��>�׹�3��·���W�K�4�i�!�Xii���Z�Be�I�p'��fT���z�4�Z��@�k�P��aY;��,�ika�����%{�}�`��dJ��̀M�|
�Dn����p#1Ҵ�1��3i�L��6__�yS�S9�CPࢮ�-��;��QEP�<��~�P�[DI�;f�*txk7��=�d^%��z��A�L������V��>3�,�<���W�;�Y�w^��7����]p�c�c��`���n�b�9�$a�]G��bmB���\�(�a��T1�@f���Y�')����Z��1�v�Nk�ʳ��@�n_/�`N�iVy���0$�"��7�k�x$>B
�q���a@�1�.}�7r��#i�2�|�����YQ^�oTg�邓8e+���N�3h�+p��w��;Zn��Z���:���V��>x$��B�v�K�i5�(�e�S���H�.�F�#:c�p�7��r�[�f�d�L9� ��J°�8���㛘�n �8�;�=���gj���s�q�ZWv�p��A�;?�G�{u���5�ZS`F w%�#YQ`�:�x/��G�TVN�f�ԟ�B�#�LU��68߳��뀭�JV.��p!��_μ!�����f'w��ֿ�>�i��$hdn����t�j�?B-�_f�������\�c�X��G~4�m۵����6D=�Y�ݭh���g!��K�����)�%�=8.�E�4�̯1y�`�����7S�g̸,L�����~�b�8�V�B"���۩�Z�cYw��$Ak(?��6\x���˞���3t�E�ľM��Z5`�"y$�߻W�F�1�ua�9�
 gx�%����iٻ��Z�kAhu[g����D���r�SMɓ<�e��2��<�RW�d	B�_������$ʖ�I+�=0�1��a�V���Iǥ�؂�Q���Ո�&��+]�����SE�r�Aj��z#�#�m~H�����>Ԟ��LL��45�����`׏33��ny��;�},�_��ϖ����r�|��-/ګ���I% b�'�ov�u#]��I�᷏'�`><���=e+ӦYy켛������)��Jy�!�a22��L*��/! ���3bƩ���P�y^�ym�ˬL+^��4�a��$F�{d@�Jig�Tl�`l�(\�ks>�.�J@���k�8Y�R�tT�"�x�򬚫���_N��ZC���L�Xe�q���;���.C���o7,�m.��D'^ K�gXHi_�k\/!�6mڙ�汕в�%1G.Q"��GVm�]���'��U�݆� �ف�PƫUz��Z�pʘ�'��V0��5 �������aI6J�L��g��@���4�i�Tؕ�@װ��s=��z��~�;_�|$l��x(������m�q�uaɒ�>��Lp�;�����oQ�N������s��!�FVR�� m�o�����X0���E
�� Q����Yz�v�lbgO��,�thR�wK��&v����es�w�N7~i�x�]й�~$H����՞��U*�������#�ݻ2��.�Eߝٰ#�~�A)�p�^Fn��ʰ�e��Mx��PnN	�z������C���{�I�:�F�T ~_ȓ4�9jT�U�� �[I�O�X���j�dW���^�rH�*��K'���FE����i�wƓ[Nޅ5V�!t(���T�hA��Ԇ�A�/���b�X���>@��m�ݾ<�Kr@�a� �v��oȟ�FXW�\*œ��q��އ&4�9f�[�����3��a���F.�D����\D�XS���"��@a�&[�M� ��!p3"|b�U}�A�,-�>mi��,v�/QNȝ�%�y�O5�I�#`Aqج�[���ܫ8��^u]��(�a�xX���o���n�Ne�s�<�|�������#ԭ�Z)�=��ŝ%�C���e� ��2_Nς8(d�;������#���-�Fe�C�F¼�db�Z�sX�#=�ȉE�:��#N������2\n1]&"~����{Ԡ>-1=���i!m�+)/|��R(S�܅��A�tV����s� ��V	i�
��f�&I�-1-�V�$иp�C�<ʎO���ك�JK�hܶbܟ��c��v���EY��1�aVI��S�� ���A6c��7�iNtLg���<]l����}�����U4���Y�k�[p���I=��h+���!��Į������M۲����D }�� �p����j�"�h�������I\,x8�2j��~ٴ���5p
!c�ٍ�c�B�-	�b7 �q~���:���ѮA��lXN+�6QC���*㸜j��1^s�~���p�aB����8 ���V\�rD�z���:!����D�_Y��g����x�����x�i�e�@�����W��8��׼�ҩE_� 2�xKz��� ��N�_�kiF��`)� ��; ��xk��r4�H�-��$ǣ�vX�}��9��!���d`O�����6)M�E`�g��/�fZ��S҄?��u�}�;tM%=�8+��mUQq�&Af���n'n�l����_x�x��T�P j�CG�4܌�A}{��p�L_Cډ�Oˌ
����1U4I|��Y2~���`@'I�����,9:�%�E�IO�`��Ʃ���r��9ɞ�_�;�M�!�B�^��,�8�1� �­�������U���Ibs�Id��B�.�K����Dߴl�f���Q���.�A?Oh�ê�3�8�.
>��Ǐ��?��A"q���E���Ŵ�yj�o>!�T��n�fJm��&��.]w�'���kؓƍ�3����tIϷR���u^��5�5�}���t�N��P�j3�$k��{l-�ۘG_�8�j}��a��i"d��3q��G<���0ik��}Ød�%91�m�S53h�Ӭ�w��0�z���Q�R�ٵ��VU[�0�yL\�r�l�\P53���]���ʈV�<3�6��k�-�sr���>�Y�wlM�ǴR{b��_���Y���z�=�!εPcU�ț�5L�DX$L�[��'�e��s�"<-�9��4G��^�wT�Qc�BF&�I�m;wm}��e�/i�(G��F4���a��$�t���.H?(��ބ��}�����S�2`���`A���p/6+�-V��ih֝x:�n��TIr�*N�n�A��C�b����g���tO����ǟ�e|�a�8�������=3���\�A�+K�Rd۬Z'�+�7�����a�M����%�]jo�.#���.���������9֡S����>�x3lA�ؼu0�ޱ�p���E�ʧ�����S�MO���:�'o �A\1�1V�=��{��*��0YX�n�y����\���N�,Fx��[�Rs3��>V�Ve͵l����E��7�����Z��U�CfsO��]�vf�Âl�g\��oo��\�J��hw���PsF���h���~P&b@�Q� 6B2!�ڍ�5f��s�.\!�%��p{���o3/Q��`ߺ�y�	g�D�XN1t�շ�m�V��H]�}��_�@v��l���C��|.�U$~%$U�8A$��_�~NEC�� ��=;����p��6o������Q�@�"�1��t+�?������]�����8m�&��;t�xH��/(���n(��)��*X��8�dҘ��bxy"5��cjikA����)��̭��'xzr��L���=�?hPW�+�_���<�F*��vY���N.�V�ǌ���h� a�
|���3�!է`n�����k�ѵ鸳��ḧ́g	��-
mړሑX���[Hs(�+<���t�u}V�LՅ�qg���Ղu=r�g�1s.f�r�H�V.�T����#��;dK�h�o�3)-Y�!�����)�ٕx��3oH���~G�|�e]�l���5̆�<!h�9����&^૶g���.&��
�����-9 �i�}�
Bw�S��*E��Fw�℟sv�)�P=Z���;��}��$t�iz�D`�(B�w4�:qYO
f٥jw�P��8�K�a\��Y<N	>�m���Y|4F!)`��-���f&��l(���w"i�b۸�0?e{�|�O�{5���J�o�nο2�����,y�565	������Q�7�-���u0��L�$Π`Q����ɚ��$�D�Ƭ����B^����nT~V$�h�T3i׏��+�5~}�}�';�pbw.��{F�Ґ]F�X���t��#;2Π����n���)`cܞ�<(�r�|.�yWB�E�Y1�%+��]�;��m����_�]�cX�K[������Q���>YS1�#m���sQ���������>��W�3Go�8�"�K6K�	��
hs1]]�9Xr�h�K"��聑��qDN8�ҿOUd��XrbiY���٭طЁiHv�0�s���J�-Eo��������F1+�ب�3��+����1��a�����$!��^�'>��1 ģVS�%l5�ȣ�k�`��=����]/������qLĿf��qvV��N֟�����Bu��mh����@C/���,��Rx)�����1d�?̼�/6�d�)�����8��-{Gt��"���s���2����f�Ԑ1̢H$���$ʙ�T���!@̕Q��xG�`v��X@#`mP&�Lz�`Q��Ȃ�W�=��Zr,O�TGݚac(�(x=�.��=v��i��G��vj��8y8	�~�_�����++��������W"�� �?�a�.��]C v�5��%��'��$��A�i)�)
�@h�W�	�]cdf�Ay��f���!�(�)X�s�����]�y|9�T���&��8�����Mf[]V���l[Fg�@{[0�"�"�����)�'B�{��S ����Ԝ�?3k�
у/ɰ#����^
#؏?F���G̵�����zi:${H��դ�(��0QLC�6܋���b;��*Y��\6�lB_#��%�uI�i�!������%�VC4ϸ�lt��X��Տ�w��|�D��!5X�D��(>�J�^��'R_~�����(l Z΀�{�F	�a�r�&  ���?���D�أ�h=+05{+bA������]"�5���V�絾F���z���I����ˡ�ϰ	MZ���Q��z~��F�NSI
���L���V�(4y��K��t�!�7�(m��F��s�2�[�[�|��(�>�q;�s�Ǽ�7%�"�<�-�k�����&�!A�����[�N��Ņ� mBaCp%�{��9L���t�eD��z}�*��y	-�s���t���;8)t�aƳ�[�G~��ϱ�壨�z���`��ڄx`@z��h����%D�,�j��8n�
����b~^̏�a��Ǫ�C���^p<LeJ8�����U��<����$^b��.S�%}�Y"��
����L�*�'ՌH3��v�7�BS������������^�.��٨0�H�"շ�I�<��e/A~�AWL��bɶ��d���1��"g�%�D��QSo~$z��8�m�xP�	�p~��Xß�y��`��&�I���8�6`5�A��1�^� �q@�������������vd/������7���# ��P����]&U{��<bS?���8Q!���xP�Ѓ���w̴ϻo�Y[�t���﯏���ⳃ�-V��jlM��n$
c>�h�jcТ�u������3����$ʜxg�&��˃(9����ƊwʿP p�EԷG�g�_�5O�qm6$�~��~1��;b��aX:��VH�����/�y�*ܠ�q��Qq&�s�y�9�9I�(&��'�iv��������������?�(@c�{���j��}0I�;z��P��ʱ��	{Q�����彫�e�W����^�wJ{g�WA�=�G��٪����tb�𺵚�8Wv�2:13@��6;���5�U�+�ҟ�@1��b��y(Z`���nPH_	~��6��L�\rRɘT-�8�5%tx)xo�)�z�Ό��%=?J9kD=��a3L �lI��;���H�Ӗ�9J h���Gbr2U��{m����
��p�2�hG�z���F\��,���Z��r��e�p��<�?��y�m�����It,�b|�b��a�t\��?T����>F��;,3뗶�h�
$ɑ	S]�����؀�&@����@)x�&��<��fA�h6c��~Rެ��c���1*�]�.f�ɹ����ݛ�lE��qZE#��'���{�s�K�?w�&B����H������C�����Y�����$گ�\~knjL�yb�� �^"JSA��9g/i���b��v�Ɩ���	�t��@�&��B��_ ���~?��\9D*�ȳRI�5�>�E1z���;r����.ݶ?������bw����B��\ը�o#��Џ�}m\踊):˹�j���[�dkf��U��|��E��JCpi�ye����Cy�}�A)�Z|�t�S�<��ǖ��zm);�Uw!�֊�'��}�B5o�An��S.wIQ)d�F��w��(�"���`"7�O��#��W��r�7ռӚO`����*IA�����۝Y,"��p�L�+J@�5ګ��U�rI�I��g�`�qBc���'L���+�q_*٤i�9�R^�,*�Ci�XB�AvV����������?�-zjd�T�^V׊P�wk����%54�I53x�wb���3c!�"�Ao�����,f����F���kL�^mT�;����.wK��ǩ�@HR�N����õ�#""Š�蚧Sy*��}/��-�!�y>�c�#�X��C<I�-P>��^��
Z�@�#5Z�)�1����e2ϒC�3BL��w[�A㋉���G �4���"?�A�(d��YS!�b��5`ԐTԨ��O�����\?(c5���@�|#d���~;�W���M�z"EG-���}��!|L�N)�"�dT�͹M=5�BS���g���(��X_��oя]X5�m!�����k(ՠ�P�)�`rR&�ȭ&��#p�&K�0�v�}~7Q����sû�D��x7wIhH|�q�s��F�X�v��:�	��ƝwE���\��0�-*�U�z�����՝E4<��"{ܠoh��ф��*���T��X�F���+T���@ ������)��Q�uJ�������7¶��ou��6�a/��xi�=D�_�D ����|��e}O~2�hd��n7~��4�G�궣D��Tm�ތ7���7��J����rJ�(��-���X���ji�?�+<PB7{/�Z�I�`!�I0p�E���k\�y�x��	M��In2SZV=����2��>��� *,;�w:R`S+��X���RFO��hK�̒_���W������~��z^@���j�l����-������f�rE%Q��ї7�f�W�az���VUdY���Ƕ0�n)V�Y SS0�u�XU�
��_�����?��M$;h�:S����)*�cy̔�nj���Nr�2�C�,1	��A)E��^|*���gu�1����if��+�!�C >�&���Y�&��o�Į�<���kR�eBr�tԜ�E~��|1�C&�|�kQ���L�T��q�s�Z���%�����m��[�mR6F�N�L<����L�(�M����������ܹ�f�a����t�/�<���,9 2�A��@�Q�7��떽��ZyK(K�'J�4��-R�߲�.԰�*A)�?��E��W��!W-{7��L�*�.��9|�NJ��|�+����w)�X�۩r � v��Ł�LV�gj5�1��#�������D��[�;�Y�EvL
�^y��Bg
Ĵ�a�ϵ��&s�t:���9X�F8$߅Q� s�p=��y���M^����D�Y �!����Q�/�M���^����+�i3�閽xU܃:(a�b�*;��Ū"�%cSǫ��+���V��:���s4j�ԑC`_��M��`[��:�sX�����v(t�ʐo�_����a�j�t�]-����[T=�5�������2���
EI�I����N�:\�>���>-��xa���ۗ��p��v�dz!�,kE�ڨܭ�h�4�2}���B:����X�#ߟ�Q뱂���j�^{������AbÍ�
��6��N�rY�,�X�u0�G�m7�{U)σ�@��!Dp�&j_����s�P/�@�餱��F��x�l� �:��\$Cx?JъD��j2lQ]��ͦHs���	��d��&�@�<������Q[�kjޑ�#�%#�}�i7H�}��bJFh����,�zr^���t�>��n��'�4��T
9绍��o>*e+�Xm_+��}��:�D%)���-t�(�PȒ�8�bE��l��Ku��[-�.OĎ݊ui&�$��6@1Ȥ�b[{��
2�U;�J���%��e��Y2���|�Q�R�h=����B��2Z����cR�oU.����eVf_��׼A����c�Z�5R�Yt�\���j�R��Z�.�n�X�8�˘���@�����Q�h����2?ө��p�����+�^������W��A*����5_߸�L�\"M��X�ԃ_X������T ڄJ��f��
u����3fq�ϟ.�M��qk���{���Ԃ{\K����H�R���zvJ�W�w"6Ρ|webU�F{�$*t��0�g�5����+g������v�\+��Z̙��*[I�C�b_XZbχ�#�M������E�kW��̑[�A�3���,3>���M>u�|wt��b�xp+B*�dk�nX"�����B!����@j�D�~͛��� ʎ
g=�9�XV�
`:Z��ɻ�K-әM?�L�L�@�j?���8�����`+h�z�1����&ӎ[_2��?ؾ����{�,��$��}ߥ�E�X�Ƒϴ7z��7�C�F|y��Cצs���O�&�U��LT��_�lM���R��c�=	W�e9byε]=����ߘ��n�]�)�`&����H\Q�C���
�NB�b�2�Q]������C�]A�!W;�����ф�g����r>[�~�MT����Uڦ�trW�(���2�B���⽝V��LD���W�&�b���⫤������A�Q�ֵ!%h�7��C�r^rF.7�j�#�Ba�9�?;�N�>!�eT���N������O%q����1q��Sh�K��#���f�Hy�T�#��>2��9� 0r$-�� ]�5�1pլ��˝��3*��,��l����1���"_�E�ض3�꿽`C����T/�qdsz�஥�b\�O�~���
=^M�������)-x������6��@zd�S��q�RM��#���5%,�ї��;�!fȢ�6Dc��	���8�� �]�9y�` �X�T�:&/�Y6���� �,К��jet�v��Ha˒��E/��6t���X��hZ�q�3��ƦޜI{�>����MTI.p"�T: �Gh툷�� �F�5�uɽ��s��źm�
/uE+O��E��=82V���ks����F�^'��}a<FT��?Oaz�h�v̆+x�fXS��#C���.+����H��/�B#z�V�WXZ5�u��u�
�7�a'�� ���f`^ln�u�i�5��}������u��I�aw�#��4�����ZM#�{��so&�X��������^���㌟u�y��|���M*.�UǋR�~'S�fڳ��!��]#pTWLm4��*LsϨ��M�ws���p��"sJ�٨Xi�D^����[�iT�w�V�+St���$��G��^�*��3�n�5���y��kRx�~Է� �y� A&��sf�-LLh!"�%@(8��֏<k<�����A3g6�T�f���%�����c8�R�v�d8 ��ě���<nΖN�0���H��Q�ԒI���t-�2�7Y�V
)�
O��M��¤'�>zM=�W�
����z�\��z��3+
�g���}��ȸd_: ���Ο��\�D5�]�D��a$r�h*A� E�Q��[)�}��b�w���-�ߎ8�
7W��[3dM�("
?��+/If���iw�I+~6��+������i��1�\1��<`��ꫀ��T�B���	H��}�6��V�X=���ךr�{���.��A��Qgu�~;����?�=d7v���*,�rm,V��Ҷ�#˧6��t ��ER쭟Ə���m�A��Y�f�mV$��Wg�k���@��=�6G(� �/�m��h�KFjv���/����~������VE��ɃTJѝ�Np�W"bf��w��y�}[A�+�=Tί��[����vt�� ��H=ikM%��ɺ��Q�1@��}�u0�ؐ_InhZ���
"KMsE�ۦkBMp�"�IÒ��LW��=#���������ɚ���	�:Fޣ�ஂ��7<k�?��2�;��dc���@HE7�{�}d�(����ȯ�>��Z��i���gT��i�hfYk�G�@�ch���p?��5�a��w�_�2'ѱ�R�����Bᗺ{'�դ{{�EX;���F�b�Uϳ��){T�C��9�D6G���[����j�[���ى۟T�-'oP�g�)��Q2��-�#�$�ΐ��>kq8�\�|��C@"M^
����k|�Ȑ�@�0�ՊO�i?�Tm���k*�9��E �Z^WW_���ǹ]��~@ ���Lx;r�A��6���Y�:c>��r�����,^-ч��eL{���a^ֱ,���M���7�D�f	7�G��==^�p��<R�wM'�$�6�A����V�uߍڔ�����.�Ӵ��F�g��M^E'�o�ޚ���P�����W)<_�w_o�f@�>�vFq�$Oe���F�ר���aó�����S�"����6�Z��w�x�`���y�x��=�C)F+�EwK�xV���l�/�>T��� 捈҂Wv���8�������v�!�E3���Y�3	Y���鄿=x�+&p�ͪ�l�#�2j����'���9���[��_��ZZzsO����t8�n�3����5���H:�����ri�r����!�`�A�i����E��d�<&��#=�/T��u�L��[����S��W���9$?_���N��-�`*o�r�q��<�xC��C\��1{:۷kYt��`L�����YTV���k.QrQIY�,]����M]
��|�O���hG�����o��k*;Wr'�7�Q_ʻv�,���!��^�b�P	&'M?^z5���2f�t�2�ɦ ﴷ]�-g$q��6^�}C��T���B#�wMOⶹ�oJ(���N�$-Q��Z#�Á�q�ψ\�	��J˞6.Ze��5�E��~c�n�#��c��� �
�S�5:a*��lQ��_��o��!��"��"�*�pi_M��q� ��~Ƣ�E�<�4�*�i��o6��Y���po5bZ�S�޴�ItJ�)��\.��A�d$�SXsaŰN)_��E~S�QP�#��`�����
8���G�%T��\��~ϧ�7=Y�3Z�����!*�evk����d7R`RИ\
�T��)p�zf6�A?\��YCjE��s�RwYa�34��WU�yL.����ZІ�'�҃�+y}Σ�6'	���s~�@�ۖ|[��{y'E�-X.�[N�����V>�çp))�M�;1�C!OmBƼzR<Y����F��+��hRҜ�{6��nTI@sH���0�u 9�TM�(��
kK�^ӻ��7�)ld%���$]H����<.*�*���[ �0����VRF���$��ս�32_�2��6��@��J�Eh�|���|Rp�G4��ȹR��C�TC�S� +M�� �S�y���4��]aɇ]�r/��Z:��WF���p}a�+�/���c�C#n��ٽ�*A�7��bɳ-6i�Q�`�h�7CR�>?�����Zt��Ŀ�<�Pv�����%���p:��h3����~eG_�%)C�5�	˖�E�e��^�а5�gm3��i�t�m�%vɰ�[�kC� �d�R_4I�f㤒�"��FET��~!�ߖ��/�5��$�B�x}hV����^	�K	�R��/" HٸZle�P�8��7M~��Z
���ͣq$�7����Q
�|^��Z?Ey�	 ���ڋ4�%�`��m�Օ�L�Y�ȊN��_��!z3
FѾY��R�Zj&t�*�U�Zoh�2�EM^�^���!7�r픔[�0	�4����E�g�=����E���}�m�7a2��ŨsR�J8��|{�}*~k��{�UXi_��
�)�����4�MRf@��8����)��_�e��]��֔F��;�0�e����}jē1�h�(��eޑ�Ð�hd�]7���Y��a�*x?[f~�/(#>����~㟽��ZT!���p� ��C�V��D�'���u+�o4r�uV���2�vy���X\�Yۊ��{�q�lH�!�$�a0X3h�)�uRy:A�!���|^�s�8'���	����wM#V�s��uV���M��Z�rO�F9@׉����(�Ԟ���w�k5%,tmkY��t ��m}����n���GG$��
٤1I�z@���y$f�3�=�]̉yNwm�ٓ�j����psPy��z�n7��#�,%Px���F��dw�͌Oݐ
�%��̔WE��.�B��eap��&�K?�B�:�l�_g?'!M��#�!���Y�}Ƥ�-��]�bi���T!�f_e�y\ ���9�jҚ��bf�Bb@���z����Ѽ�?:E���bR��
SfI�V�i	�sM/D�֏����hWŌ|w��>힘���,N6OZ�f�W���y�K����ޣi�f��n����f-�k��9X���X���eA����1����ע7SS�����v�a�ޤl�~L��~T�&��a��*M77S,
�����Ƣ��L�P��@f|�e��;I�i1��y%��0R�N;��5�)����$d��o�/J��V���׎��=\O-�_��[F Mh�8���Y�P�F���i�(�{�#z٥����/ �<�� ��
u?�i��%;$s��6����m3|��NB��I�_�����#h�x���nI�p�����z����RA��
M;5/*�h`�+�)H2�����8����B� M��r�N�H
o
������-4��?޴��}��1��$mLH��*���ɖ�b�eu%�}��!��t�	W�tݎ滓-�`4$�f��Y��`��*pX?K�[�O�`�����"C��=��ɴ.�f���S.�?ݫ�0�պe�+�RN�Ne�N[�2�����n��A^&�>�TB6{C-�u��~�4����7���h8y�'�/�)��Y[�V�۴i�Խ��e����T��Ovw�d ��
���Mۭ����ܿej� ^aK�s�!������|�����������K|�zl� �**^(ǀ=���&�h�	�G4�.#:0@'�xMiY<���L��~3a�>mMa�JC�xs�Hǈ���2�3��YgFķ�I(�(!g�V�`ߠ�����<�߯L�(E�!K�ʃ� � Lh �F�T���<��6��9��~���X�;+�(� .���$;7�v�S�/V�Ǽ�O~�뽲��P�1s���9 kǣ��\�	�ƟLab��Iߕ��Iq��6~�`�C0e��f�v�@�r�x�o�1��Uk�6QQ��,b<)��,4`�Ᏻ�vɲ��������Ћ�$Z\A&g���1X5����"���Ui��z*,:$���n��H~p�9�P��\�B���T���_^�Ol�a��	�x0Y��E���Xܰ �@<su�Y\�|�,�n���#tA�|� kIT�irqt�
�����������
���P!�|�˧Q�^�:Q�٢j���VDu*�
��#"@�� N���D�J���s(��^�^��^Uf,C�n;-�P�0Sp	�B�<���t:�|�/��u-�n�%��'���.m��_ȿK׭���7���/*ʔyb�z���>���<\�
*��ŽT<�*��"
:���(\�7K�%{���Z n�&ɺ�üVn��2̈MHZ'�ﱭ��k����k�\l�@B̊�SZ%����^��k��w�1�hKb��[�qp��Hn�9�S΅Љ>�4�e�1B����ү�1X(����A��̷�J�!=�zNr1���/�W��a_g���l˒��Sm�sE�v$�b��T����dA1�/78/�6/��&�j��6�K�qU�����ѕ�p�wD��$*���Q����ɛ����Dr�Y����)M�ӑ�H�=w��T�S��73i ��{��8��U��ރQ��QO�~�Mur��݇p�����Dn�9�����������\���w�*���K�wK����[��f%	�ޢ/�<2�S�qÇ1���~פY�8v�Iח��練l�O�\��[0�&mn�FC!C�0 ��w�PE-ٱ��$���_co�ž4���/Pj�M� g�ݝ�Z��MM/�{B|7	���ڸ��&��77�@��n���NΜ\%�e��o�$:�>�ȫ��}����-2���!c�I��X�I�^�����w5���7�rTsi��.��S�v�5�wg�ލaEE��I,�z"���y=�����@P�>����+G���v�7d�n��.*�������`|nEh���и*5��ӓ|̈������ ח�����c#v0#2U[�u�w�bZ�ĝe��m%��в�r�5�z��)��=B�c	�7�kq�lP|ˢ%�]F��ʟa"P焋����ֻ�Ãf�!��3��ٸ�ah��Tt{�S�i���N@����᪰(Ώˣ�ȓ������l��0C���W�mܐ�_�����oLq�;�b�[ݜ����2'l.M�}l}�(Z��������Rՠjzb/ �2&�iA[���ۃ�����!�TP	.�>��g�9Kѧ~��Fb�D�=Z��"&�9kghU��w�A=�KQ���P0�uj������
�����q9�Ť�z����(�?G�#��:F&i�9����Z�aZ�*ZՔ�<�r`���8	+3�Ղ|��UnhKH�C�n�q'��kN���O`d�b/��7��^�^g�A^I.�xG���W�l�k�J_a�b�␊/#`����a�Q�?�#��ޜr�� ��z/�GB�ƪ2YR�'XvA�<�i6?8R��g�xz�ҩ-:��JBkm�*��M�G���*�1�|�<�u4	� ћ<����<֌Eɐ�C��S9֧������cc�T��Sa)2�$�o \U��N���|�j�e�'�����B���eȏ,)��pJ�������X�� �ú�G|��j+@^��e�����	�.2�:�� $�B`u�*ୡ�퟉=�c�,�uNW�5M��I�
+�Tݔ핇����Gj�͆���v�;�±K-���뽯�GKu�~�ns7ZL��m��P]�8�����*���
A�Ԏb~����Y�Byٚ�f͙��T�y6�7���������m������FW��^���Q4��@���W�Q~)"D����fÕ�� p�$M��`}��x,����+�v��� �s7��b-����?�������V��ⳝ����
��;��G��WlR拲;M���
3�=~��]Z���\e�w~5o��|?>�)ȑ�l��>�s�f �+B!�y�G��[E��t��*�_��e^���wA��t@��c�U<�;�]�h��<a@���(�#=���*|��m���V�v`�=���^�bN��v�s�?p{��Q�2�j7�4[����gа�E����2(;%&`ս!��1)?lθ.���<"G�ꉂQ�'�j��f�A"̐Unr/x�l�l�����y���-jh�ɕ����0H,R89�a�s�Lik�?q�5�[�=��`���h���%h	��Aj�������9�$���"�<�qf�'���
��С��j��K�\Eo��Aa;1xI�����9y�|���1���tK?��}$��>��LX�L��*z��0��`$Q�J�kv;0쪙�ۡVN�}�|�L�	�������d�J'V�P���M��³}���)=��Uu'�U������7^�l��#����Pp��[���\$q���׀���O��,��z��Z��U�D6xf���BZ���gK�.�*_#�ۋ�*h�	�D\�Ԏ�J���-�������GaĬv� 8������c�6�<75b�῅9���i'x���3����$+K<��v����cpV<��x�ܣ�|��ѓ��ʁo�/MtA��A�^�D��
�Ahӄ����H�nR�݈�;�e2���烎
�=~w�ł�O ��{A-?�J]����ǅ��:Yę❫%(�t��QV�ڃ��m��(�fH�"4�}�;JKJY����_���ܐ�ı���4����a\ɇn���)���7?=y'e���e\n�<��_])#N_#�������$���Ǡ�v��(�G�
�Eӛ�u�}ڭ�c1)��>ᢛ<<�����"�|9^ը����q� �Kr�S�k���T�$Z�3�~.N�=J yk>ݥ�G����E'�5wu�C
![]#{Jq9B�,�Iq��'C��Qkr:���J;8��soT#	mh�����$����ɉY	��A+|;%���e��f�<�DD.I�&���O.q��m>�����ڊ�3��"C3AmN����Ŭ�֔ѾM�cd�D���GJ;�j��Z��΂�a�nꩥ�ߦpY�9�������f:4²�-6��xU��u`(��d��g G| a��ẞ�7�c�#�$`+,�*���>����B�U�zB�����n��
��w��N����!M�P��S��y2|�H��g�G1Va�Q`]����A�8���
0�(�@�[G�Jjْ���u�z��M�����Z�i�k���6����*+,���Vɹ���ӴQ�B,��i?�Mb�Q2k���`!�Ķ�)�	~nVsw�ܗ��d	#ߖ+j5�?��x�C��}L2�&��n۪��|��*ysG)�]���Ҋ�IΛAy2��T�A��� ����&��|��'%3���}�"	R�8}��"	�J�Tn"D '�#F�B ��V�IH��u��H�C�ڹ�1U����\��& ��g����al�4�4|�����tH��O���-��͵�NU��)uP4��h'1�N9	څ����(3��G�A�a��0�`��c �Z1�e��-�����w�:oR:J�]Ӕ. B������6���E���S5
=>��E�w��V)ЭAn�>�&�&SN���mls3��<s����=���AسV|�N��"��G���P��E]�`�M�`�0�}�a��?d(�E��5��Ř�#��� ��Yx�{���|L�k5|m(-;�\�]��gB�ö����Ҟ���mq<����\-�2e����v�Uۤ�O�v$	���%w����4$RR*���M�<�����dA��\���1Ŵ�ԩ�������j�}%Ђ��H�#cjj)@������sQ��mgke�G%^>M������n��
���5�ϓv�Y=J֕����ٴ���sr��#��G8�����z/ng�H���4ɴ���dL:���Usyr\�;A���ę�Zc"�����$ȧ �x|����
�ɜ�cF��s�\oyl�R��j���KKy��fC�6ܐV���c+3(�e1�7	�r�f#?���Tq�X�B�6�aA[�<x�Yj4Y��D��Si}�����#�6��jiǹ�}�0K�(�bc��Y��Ά�
�����7zU�W1y�U۽��ꚟ�3nQ醯`q��SZ&i�5Zs�b�o��K6���Ça����݆��n���c=U�0��A��N���)�`��󎻱�<�`�H�K>g������kA�\�l/�;nҢ�~�' I��93�E�L.�[��6+�B��Z5V�(�xT]��pmK��w��v����Z˦o��5S�/�=�����$D�}_�L2Ja�~N��J��U�/���P;3ۘg�54t��>z����Gz�1}{��/z�s_��p��,{O �Ԑ�$	��[��I��$̃�3�lE]M:K��[<�B�脅��2�}f�^r������10E�8��+NE��/*�w�C�px�Zp\
VM�m�S��;��	���,Sf��*�F�R �t	.�����VsX.�6f�� |���;4�B}JԄ�n�y�1c=Tl����>��L�%e��0Ӏ��c��!)���������T�I���."����3+VS{Ã�q�
�i78�:��6�ʧpa��V�7I�Rvq��e�s�S)A�"��B��L�I<��@�d(V��O;E��������L��n���P����9�78I%["���o@��(�+Q���=}?9�ͳ��P�2@�v��Vm�^N��z׾�X�s܌t���)�SΛ�!��� M<��Jj����e��z-;�"����w�Q04��s�h�~���Y� ��-���c~�@�W2Ple�h�M�����롾�9R�a�����V?kA�"���`p+=�&��Yl�m��u��R@	a�D�3�&��-J�cQoϸ�N;IL���!;h�%��ޝV�(�@�N[���z�mD�u�)Jl�#n^�`�s��A7��\�������A3�
�����Qb�2��g��l���
xm�Z Ɗ��F���i��>��ݒBC�!����AFP�������D����M)g������1�J���f�&i-�,^ ڔ7	U����@�C�.:ilUt$I���l>�gs��U�mv�݈C�V��ߜ�d��_@���l�b�uLP@��±wjg�=�%�J!!	n!��B-�����J\`�d����:2*��yk�Iʘ����GM"[��g4�ðI�9S#�\�{�3f~��n�v�̡�x���Db�%�JMg�)j���I�Eb�P�ɘ�V<���m�v^��CQ�q˵��5z���9�f�D�Se�|оs�s \8tR!*I������ ��R.%G�!�O�ԷRm�n��R �b���6�ɶ;�ky��;"꾢� +aee����pk�kX���l�$��ͣ)�؍�Z=��.��]C-?S�ߧ}�!���ϛ�E���Z,��6�\��Pz�C���h"F�7?k��<0SZ�֙U#��_�w��J��n�wm�p�Vö�0eJBc�=��s���K�s�sw�F'���(-0��y�!-X����#�&÷�.4{����#>nŪ0v�HM�n%����4I���.D<���H�E���YQ���G+n�&�%�Qˈ!��v5]�kIY= �h9����\���ϑ�A^#�ӡq�Nڗ���4�*D!Q��{���s��!2OO��Ǆ!�!����>�Ӂ���֚Ǽ�Io��CIX�&ꆆi렽z>�#�d{��doZ��V]U8�%n$�7�h�P#�Ql}�zp�A�c��;���ے�-H��➻�ЊY����Uǭ�L��>�S`��O|,�*k�L�V�����������m�;MU�5�AGٖ9lS�� ���U�jFX:46v*_c���} |�� �s��k����ol�8Q���w���g����cE��K����~3V�F�)�R�C�X����.������B"���=n:�wsZy��7R���f!J�u�x�J��;�C�D�x+��*�9o�:�XK���l��`)���B� Z��E�>{���quD�^4�O;��¨b2S?�ʾ'ߛ��a/�̍��Y���"'��\m�5��=��'?z�hk���&Kx�
�ZEwnqi��T���S���≔�*�<?h��l��L�Io�g�����r?��i��޲�7�����ˑ��-�nx���*>1Ia�a�H =>I�a�կ�i&O�K|~\;�Y�X�nO�CTi��i��b7���`�Q������x�p
_	�7��>��Yks�|(j�K�T ��AG#�N�7a0s'�̝�mba74izo�S�[�d$.*vw�ua?�D������q%ݬ3!�< =�IrkkI����8r��9iy�}
�zP(�M�AdW�V�v=�����܏�� ��g���4��5y)2:	�����vV��%�&N=�d{���,�I�o�iK�G��OjZ~g��[x��E>�"8��;��*�q.�x<'ZU��X��	' `}J������'��1Lb���n�SOj���|p��#��-3F�gEQ�Xd��+�-�t���[�,c�6�+�;��؆�j�1��"0�����)�I-�]��6Ci��hO��,���{�S����{߈�/b��gO�z����[�[�$YЛB�3�yL&ߥ�ҭ�A�6 �4b w�gL֒������2d���	����ϊ���={�@�R3Eo�$��=�!��rc �P�Ck�&��ٷD�_r#NRj`��.W���*��I-�%���"p�?	�+*9�3���`������4a�k_2�HՕG�rT�~ai���y�`�z�~�pS��K�S۰<S��֯P&G�Åt����~�s}NG�tͬ���� �B�h�$������(��C�����^7���X�8����kEI�6z��" Х8��BU���W*�(F�n�|G�18�pA�f�����R�� v���a��F���̔ݱ�Pf`����Ρ�-�I]gj���6r?E��`�G]��i��ء�5�T*�^�*F�#_�.�0`L3!og��yP8例�B��iD]C�M�{A�Hf��u��v��y�r&�n
��q;�>�5F(sWL�Y��w�
	�K��"�(�T��ܘ7,e�V��$�$A���#dޝdss8��*�֗E����?X�9��x��TQ�9P3}�`�6��o�]s{�v5}H�}�QJS�;�H�}�u��	�1e����+�"Ho��7X ��"yP��^������Ob�MŔȿ�
���]��C��2 '�����q	l oÜf��;o��瀠�ݮ�w����&�`���k26�6~�I;��Ө,���	-��|�^f%�Q`��n�[4�ug]g�6�n�I���,�]d���N5�V�d�U(���<&Z����*�N)���h�7�i?�j�8��U��}���c99��rb���X��"�*�S�k�?���C��U �	(�h�DmD�#|�ԩ���Z��E,<��$�)Ж�G����8�]�=�=و�g'	�#��ym��:A��)�S�?!��Hɂ���(*e��V�Ǔ	d�EL:��D�ԕK4�#j� ]q�V�B;>��Q.�c�'�p(��S���ڼAR�?�P����&��֣��۩ش��.h��z�9�h��2�"���� ���xƛ�Ć���jX��bb`B0h�"�����K���#�!�&���������y6��Ku�Q8��X����\�Ȣ��:�ڔ1�b���{�=��sܖf�M�n"��BK\�0n7S��;��¹:������p�6	z:����b��Q��	�2ݚt��!��v���@&��l�-x�jc.,�%��"���	%�tK�W�t
�"�B&�:�5N��ʵ±~߉U�Q�-qY2}�#I��5����yۏ��I{Е�\��&:�
���Ra���xlt�����G���d#�����fc��2\p�Z6wkIw����k��<W�~O2��B������,%Y;��%�S�݅G\n���sG*vE����Аζ6�[�d,7�Y�ӄ�k�yu|��F�>�5���"���h�Z�P�=k? �)�q�����`��L�̖��W��b2X��<{�e��)Y�:��j���P.)��6���3��:����N�ܘD��g�a��A��j��yy��Њ��\�%��
�HC�63�K����mc���n���Y����UpЊt/w�/��$�0���X�/�����������Q�y߯d�?���뜼7���k��Dg���� 1��y��!�Ψ��Z[�}3��@���z:��@$��_f�\�����	O�-�F�qr�X�(!N�N`f�M�[��f�5��=�s,��-�=ǎd��	���,bb[���L���.)�!�Xۣc,�w����0����J�!��F�p#�F/�ا��yʉ��%��H�#xi�IQ TzO�a-J�F�st4�}���'���(՚|�,�&M�X��ȼ.�64�eI2Ooc�G�u�Z="���j0^�!v��:O3�����}�L�;mUJ��
4/��
)�:Y��:��jݓi,D��I�b��M��v��lS�h���v7�\��b3����*����fb�j��]N������t�wSK �UR����RH �Q:����z�^�h��)�8F�TBy��^Gڄr�
$& ��(�h����B�4�A�B�M)��:k���E7�AX�D��a�����7��`q����z~�#y{�\GH"�b�ܭ?�������:*�n�D�H��O2�C%1���c�,{(�|����r�@��n͂�M{��D2�)X�����B������?0�Bu�\�_Y1�I�PV|1�B�Iw\� ȗL���S �^��ɵI9�����xU����ׄ��V�Vo[���y�Bp7�SD��`����9��ݔV6 {5��9�M�!ے��Y�%��D*�9��i���gD*���q�e����z���)�5�ݭx`��a��Uחv��\����Kv#��|��筐xj��$�$_��n���<�����|���y�Acz��B�7� /����!-����<�ᰳ�X��Ă�4��oӣ�Z-�$�4{�:���P�AM�{_s+pi����Fum4��;��f�D����#�������"_Qݜ��q�?¤��<eeZG_��'[b��� y0���yfO�V-�R+�W?adgϯ���(-��W��V�����T��7�[r�O
_f������Ř�w���a�dA��J%;<��T/�w�F�G*�"	1�WL�Hߣf�ʙ�O6�:�&�r �r&��n�_�\x���;�;���u�b4L�	��:D�T�
�蛷���	���"���R0���h"j����%+�v.�,pK*�j�H���CMU�HzDO>|⩜N<OiYq�ʫ�a���ZI�G�<")�hh*��k��Ҥ��T��q~�7,�5�ܐ��ْ��	pa�
�$�_8f�\�F�����>h��Қ��n'��0Up#VSd���B�9�c�<��lF=�A���f�;7	�zݖ��޳ϵp��{����\��ŏ�y��!�9W7M��ߘ�fL$�B�ӽ�oe�^���1���L�ҭ����0[���,wT�M'�� ��;��l]s��H}�2���L���#�=dg�ڃ��=��I$;���ۼgG(�'\Y����޴�%Y{�m�H�k59*�Z�@�(�]5�1%���-��n}�kE���ǒ�8D�z�㟇d�ɴ�u�h\m�|YE���wy�� ��f}�k����b���g��E����S2���A�N*G�����D��Bj�Y=��j�����&�?������6��A�=�2�_Z�!O0�$����b0]�J�s�>���n��Ѽ�\��A��!ԏ��';H�Iq���&�81pe�Rn�ͮzՂ>�T����ְ�hJ�<��/a@�f#�Q�f?����~�2�fڕ�JlƯ��Im�0��m8TGe�������O^`arxZ=����U��tu�����U�'�� 1c?�jS"ӭ���ZN�i�5����!��zs{.N���<Uz�rEh��p�_B�E�t�I��/��'f�8�'LV"S�������he}�(H��Pr���cJ�����!*t��{�g;\L[�5�7dJ��)�� �Mn���3���r+�u���DH~ �N�� ����In_�QF��-U������Q�rLC`�<����oQ$���7a�G7U��Iٽ\^��~>����Ұ�<IY���l���l$�cZ	�KE�`��e�I抝���M��r��~���BX�.iUe�αbC�sZ�Ha���3B�(e�0
���w#:��ߔ_<�Sj��&0$��,�=}c����Z����Jr�
O���^-��
}�\�䞙�υ2�c��*�璬�>�jJ2*sl��l�WR�x��؋!�R(��r�-���[�0�.�=8C�fA��l�</�w�[F�}9��R�+y&>�ҏ����|s���'��{M�;��Fہ.�2l6����i~n���9т�O����r@���d����נ,���/�he!"�H-��U"���Bؖ������c,��L���	��`�͓0� ��K��J`����ǧ�]l�n�\���d�c;��c)���1��Y%8Z%��\=`���([�"���,��{E��%HT�6�� �>�A�tA�T��1� �D�����1��m��ZҰ����m�D�X�	��9|��`��A��k�m��XLy���ȁ��ʏۉ��*�w���`���i{SY��S��G+m�>8~��U�N�6-��)%�4'��
P�~8�X����!���v=�Ԉ��7L�����b9��v�)|���'Cr����_���NP[�C��v~x+�B`2s�hM'���7C�U/��@��1X]�����0aT/gw�D[�-g\{E1يw����Bmg��m����6��_Q¢LG��J��%��V7-W�0\
uz�yii�2���k&�!{�'N���n�|��I�菝�2�ɾ��}���y��ZSG�9�S���վ���<pw^��YR��a��Mxs㩭����_��̵L�H]���	�z[ɷ�D&�n�/}j�a�-�W�w^z���5q4��ઊ�[�k-�g�����)DA˥u��>C��>3�ʝ����v�-�>�h*g/JZ�Eݯ����*�z$��q@�;	�<����h_P�<\�A��瀷�3u��1XA��>���U�Q�m̙���o�&"�PJ��fM%�TH�w�K+ק����Ry!���Ȗ�p�չ�~��Ǭ� ���<�Z��k\����iL���`K������_��d���j�����w�F/=�~"6	�M�Չ�!3� n.���NWPÌ��)'��<)��I/Z�������@�OR1��Ttx��`��I���g�a�z�!L	:���[4���l6Rk�§˕��v{,q w&W`?Q�V�2����_��ۦ���F�5^�iW�,qfA��N_@&/o��&H�=�xc ����#QX,9��|�@��j���n��:�a!��@���~hv���i��ڒ���]���#_ST��Y�w��5�������V��f�De{(#��ʦ�Mgyl!���P�ӥ��ub���&��:�yU�����"�+WRڎ���h�'���(�FU^�L� +g����p����0�����LD�Z-!������w�f�t��F/�}_|S#�?k*-��x�#�o#�Е�	r�f��,R�Y�'XU�ر� 쬟TPK�*�t�k��Or���,�]����#��q�3$ՋO�	�	bd�S��̕����|�=hѤ�>���uuߘo�$q(Kn�RF�)�x�>���̿+�裒f�֎#z����?��;�d��W�k�����a��52��-����tt�� �c�a6�M��Yp��n�8Q���c�_{Xy����z��{b����-x���2gl�
;��]+@ػ��\1��¦t�W3Ծ��b��7��B�.+�G2;�eI�&�s�
�Xz�]Ŵ��J�_)�g��ҝ��0��	0��WW��:��_��K�ڡ�ż��}$�������4d�N�d�5���,W8������$�r��e
@�����]EZ�S�Y�p F�5.E)7D
a/T��p��·�a�<�{��Ҡ����/kĐ�ó�A 
J�Wg�F(s �y�xw�{�r͹8��0AƲ�,��܊�s����M���y�H�g픷�nH��R^������1I�bl._w����Pdz���
��f�f��r l'Pj�,��=��1+�J��>a���rR��XVj⟊�#�m�O�΄��YX�:�̂�U��e���O�gW+���a�K�Ev;}8�Y�(��`H6���2!fF�bO�gA!kT����צ7����~?f�3ɴ�=h X�-}�@�jeR�y�)�>
̈��hÆ#&(C �I����&H��} �I�n;�����_���9*���Y����\��Į�:&�o�!��#�K��u|	^�H3m���>%(nw��Q�@,E�s ơ������T����P�'z��NNF�p�+�1X��&ǌB�:5}�/��ɼʸ�4�[%�=c`������( �sB�.�Dq[,�����Hp���v.����}BE�^���S��:�~b�G�Q��-�����nX����vW���>t�x�iX|��,w��i\
ХvPJ��W��9��M�l[�h^^р�^���pI ���ۺEl���u7�H�Ϥ�A��!%ĬF@�~���6��_<$I@Ⳅ�&BN���K�㻞�L.�9z�Y�c����WL �:��`��%3*�l��<7����Ç.DT �q�&X(��mo��ש��'�E�Cp<���D5��Gl���j�	Z�8Qg�)0³n2���x�M��!�O|��Q�F
x���y7t77�8c/W����=q����]���x�=
Sr�ڭ��i*��-�@-���x�7�'ጋ����ߔ���,��*_�.�*Dj �����"�� P�sN�n%�Js�k��8K�'��9��)��0�p_Av�������K��Z9�_�������%�
V�мvn�{Puxd�[;����Hxǚ��⹗Ŕ��k7�\��4T� �����x�o��q�%�+��iM��8����������	N��|�0/-�� /� F(&
Jj�5`��oqZ�d��Q6��lt���5E��v'f'l�	�s��z��S1�v�� ��C�'>H�ο:��~dPI�7Q�;d�C8��~�H�8�V"aW�W�ux�fX�?��A�m݋X`�bb�2��8�:�]�bW����"��}�(2�<��^,��Q���,>طs��W�Yn���A��C狷���̼!���ZC�Bk�E5��$��Ú;p*�0<4���eOH�d�
]�ٍ^�W�@�@���ܲ�WJ{��`1���D��X2���A�ߵ�;Q��:�RU�J�soH߿�ӭC���ae��fa���/�"^�7\��9�R"WklZ��h,�6>D�1�7�tƫT�EԨ��/�'d���k&��.�>-�	!G�ߡ{��x�較�1���=u28�NR���'�5���V�A�@.c��^��A���u<��%�6M��3�
��Ӝ�W-�_�=�W��`( f�F�7��xc���h��I.~Y�V<��C�3V����sp���J�%`��]�2:�%��!as�Խ`B�ATu>����N������_ā��OAI�ԃ��Z ��+"�A��Qu���UT�l�g�?��-�;�r���g���K�Ӑ��D��=�5�udq��Q��Z���G�2��:�"	���뤎f�e�Ӎ�x�Ʉ�r��x2����"p��t��v#�ie�#Eu>��=(�?1k��K L����R��۳��H ��P+���2b)6�%1��-��-lbr��]ZI�85t��ɧ>}⿋p��Ә�G�?*�y8ۄ�7��jL)�,��Z�^�]E<��Z����Hhݳ�#I��ȡ�h�_=9��!���3�if�inS� ��q���#mm6ʛmm��P���rX�����X�*٧�`�u�,����<��d�������҈j��"��H��%����A�Ԯ
M���>� ��!q���%�Ԗ�,�9{	�=�T9 2�k������Avv�u�:�>q���Fd��(���zH:���l����q�:#�Xh����Xo�F9�}�;�+D�ƙ�^{��勷����~�m��A�-->�ëRde���A@Y���eT��ʽqZK����[����ǝ��mT�|����:�k��mZ�f���Y+���63�J����?;�S���� �eD�a]z ���E��?�M7Pez�����K��.���Y�WOg9�Y��}��t=�^�=���h#0̥V/T(�u�O��ŊZQ�.�2��iY��/�s�斳з%EH�{c�˔�E�����"��)��֜GF�F�eBuSv�2{EͲo8��@뤉Q秬H! rY�����X�9�1��a9���l��,	[�cr�u�e���n�v�C[��\���Ѐ���K�ޑ  *)sp�������
��ˬ<4;2	���u5�G�7�j5�!rbY�S��ɒP�ݭ$���4L���<kB��$�̚��TD	�����Aʈ��f�0�������4Y�$���I<�6ʱ_��g��D�2�7�Z8)l�?x�[3����r��? N�ʠiR���� 0j�d�Sf����1�s���`پ�dk��!.&U����5�����ҁ�x��#|����Y��L�{�)��w�Ub�}��QҒ��_֔]=s��Ӂ�q;6�Ƣ��FW#��DG4��~�Y�`pd0*�o�Y�{�ۙ���k��}����|���(�Y\�,y�����b�I�2�3���g�~�V�� ����U9��	aA��;���wЭ��
j^�r�gi�U ��4��0h�I�|ZR��b�.ލ�"1��CPK�l���ƄK��M"�����*sk��''�%[��H 
��MX^2������e�Z�ʣg��P�ܻ���M=6�:ܐS�`�@=�/L�Q��X�r� 7B�'�rf �
�p^�J2V1�D�ݑ�;�Q�����~e�2�v�VMb���s:/'���5��}����F���JSJ0���ڗ�ILL-��|��l�����{h��J<>]�V�e�v�������ށ�% ��2þ�n����bF};1��ˢh�y��8;�lʦ��1\�>%���G �D��bn4E7��hX�N`QΆm��P���^�-Y��U$������M*�A�x*���e\DF��ËIw�c.�)�#�;*6b&*�c$��
�!�(.x���X���,��ߐ"+�о4B�tK��c�$�fڮ��ڀ4����=�-n��F�~��u:=�P~Q�])�xPrW ���&L��$j���k�
�"?���ׇ+%`8�Z��Z}c���ҍa�������)�.�ʜ[`��!���'ef�����p؏���V���|��f�D�>�Z���|��w��Xi>-�����.N��I."����u����D%~��0rxD��*W
C�ݺ�-N�"�C\����٨'�9���i�d���Io����桇+��nZQ��}
h�,<	k6�u��Vg����������(s�-�ʽ�UcBD��N����y�x�~.|_ԨsN�Qk����)�'Rs�]Z��"
P>8�7�IeEc- �Kє�;�vF�=Ŋ�RR�D�u�I�BU�e��3��[ =7ukw%��@�RiC�!�h��z�B�i� B	cl�n2
Όx�?b�N��v�t��pcB�����3b�?0�+���bc�-�c)�Ǖp ��%��w��ñ*�QJ�	y��*,,�M�_��;�f��V�����0߷���y�y�D�u�"�C.L��`�>j����Y\�yx���}����w��4�e�U'蠨4�P�4r�w���I�e5X^�T�2��?�ec���~��7��̥���U�����G��T���8E�f6M=� �44M"7�0Bp �B!�8�yo��(-�R�&ߑ�b9sO�����'���R������p.�N��j���3�?����qab��¨�;�C��t��x������)��$e�;%ш���cy�m̭��g<b����['���� �1J�?<ݩQ�#���h��&͢�.���f��$m\�3+� ���p<����FtS�m���WV��/ܿX���56D>z�&g�%
�>�)��8*h��#��q󴈊X�	q�HX+����Mg�B�p��G/����t7�H���I����!���ϋG>�[��磊�۵�N����!��	������Cc��n Ts��NV(���t�ds�L�w�+zU��~C<�4�[+S�G�>QY@զ� ��(f� ����ƋJ�^�ϼ�d�~���C�Ի�O�
ƅP�����?�I��@��H�� NOʍ<���;���&Wx���!4��ȊT,ٓ�<]Ub>Ԏ�����T��̟�0�Y4��`�w��"�.�� �Uz=�K{��0")�DRV����K	�0���_�&�ˤqDzʲl�Q(�����_ɀ`.x��VU��zTϩ9��y/�[S��L��p� ��ޫ�Or�-L���#t|��3^)qQ c�oQν���2箜2���zf��Ebð:9�(���rX���NVL�Q=F�g X �1�&�i�<�Իмb���V~=^�E�5��;�����S!n�����S�7�Gy�x�UZO�f�BW���5>�5/���1#����ܵY�%~�( *)y�:��P�*��,hd�H�.W�����l�z'uCl��Ṇ�_>A�M((1&Bל����n���46{�+f�r}��\�0omݪ��_a(��\﬉v��@�#�qA)2��ws�%�3I3�[kx��%�x>�!�@��cP�r����)�k�� ���H���Xf���,��X�*���k>��R�yFL E�mWlM5c*�]M���}���S�q&�
�P�fu���R��g�~	�alS���C�]�;Ǣ�o>~͜[rX�,u���,H��pN�	��
+zQC�ji�M��f.4��X��y"W��O]m`?DH_ӓ��.+�0C�����g}��p�y#�Q����<�Yt�*���"������
�v<N�c��vv�{m�8{�+����([D� �����&G&����kzg���Lw��{u�sNƃ�V��^NZ�lAh+�\d&���"�1|���Y��_ѿ��A�d�%oDԉ��R�)��6�N��/g�*�ɭ�X�?X� m�؃Ojk$tJ��6K���/�O�4�zz��1JB�t+悏:��X���y�g7�m�1Qmg����.�۹,q���4�X�r���Jm�c���S��8e�Ӱ���E�?�ٯ匦���a��������W��o�i�q�f��0�4/����㗡i6a�|BU�囘r�/k�>�++�GR͡���>*%�ˡ�`z��,�.��b����� �Ck�9C7-��c�[��~��t�iT��j��Y�׮�9�ڼ��V�툞�zm�|
�n�G���9��gJ��������V컒�m�����ar�ƙ3��zF�oʈB���vs ΐ@l��q��]0�G+H���-��[�]��
��H�-T볱=����#�2��_
[|uD*�d�ӓ� js�k ��b-�t���1ؘ������)��j�7E(��&��,�غR���;Z�ÍN9L��1�L'��������ym���?�/�x�]m�8�8�B����{@��!��/*����ڑ~��=q:a�8k����;��MzF������&�V�H��\�'=��a<�mU(1n�#p�^M�ӪM"����X���Vh"�يX�ȁ3F7�s��'�֦\�Z�F?���A�
>Ki91691�?���&�`�In�#��Rs��^�\M�����D���
x�㮭�?$�4� ��G��W��������S�C�^��<�
�`t���6Θ6e�6~~ �����h��IO��3(
���a�b����{O&)Y���d �;��4�{:��V`a�i�hT�-t��Md�q�X͛��v�����k��ݖ�Jw��ۜ� �q�v��U�H<�ka�,�$g��+��49����jn?[�(Gƞu���Z�-�pE��lC.W�fS�m���l �Ƌ��c/Ԉ�)��*6�)YY�Z�ke�&���s���6ٗ�<�p��3��l�z��.x��)����Ei<8����3p+Y��4�^Y�UH�T���Z�5;�R��������`�ro0�#��:s�,-����@7�)ڴ�>����L�{R�)��cQ)�����M$$���2�X��}��
<Y��>Gn�+sD�0b��	�_[��r���3N��7���
���|����΄�R��6,��d☺����]qcd/=��O�h�]܉�z�	UG��eT�-��A>��7���&�L���&�o0�����0c7�@.:�XmH���`ba�*x���ue��*�2�Ż���DO̖�����Ȍ>Y"��g�l�}��?[�klW۸Xv�.�[�?zo�	�:�v	/.���GN�� dz�)�Xȕ2�ć!p��D�-��WYcCG^NA�R�� )�z�6�:v� -�
9��,W�����
�,��`�e O��
�%XJ��}n#<����Q�,�`�*��m��w�y&h��0a8g�r-�P\7dD�ٌ{Җ��v)����4j����zk��E(����zb�q�v	a?q�JE���ܜHY2{����۱Z�x�8I�ow��aD)GT���w��z�}�C�������Ⱦ��T* FBl
I���!��. ��L�|bvwn5%��nX��C6F$,�d��y�v���injo��G��Q����.�.c�H�s�@�;���7oꎷEn��~�4�CT��C���;�JՒ��P:�=�ꅏ���P���˴tO���S�x���o�n钻t%Z����І�/��[��M��3�!�~\̄�kY�~�����m�b��a�3H9|<� �_cG���D`K�t�-�p�&�Dɸ�l8l�o[���h۸�d�R������A�v�-�q�%:�ӣ`���&Ȑ����*��	�+N�c�q��5�e����?�6��yi3�ofJ3��4b�_��{�s�U�^l`�+~�<!
���d�~k��f0����[�4��=u}(�p�t�J`��R�	��>~�.��N��>m��\�����:� "m