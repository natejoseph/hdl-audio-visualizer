��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\�ǩ�_����;�	��g���`�SF�Z�6v����(E�ݻ��<���� �1��4Ee4>
*9�g�Y�� ��3�I���mw`��ڸc~;V�!<���F|�Q�o�;�1�Ϝ��'۰�8n^aU��q�� K�y��l��㱫ry�B��x�!v�h�;��&!%�x�b&����_��P�,����A_2�	\W墺&�+�Z�t&q�T����!��a4|_	']^"�d�ys�d��[�k����ڦfwG�Pւ�$��%tCc�� VSq��g�����c�� k��y>�D|�#/�L+E%�*x���������B��H̼ú���Q
HO[����z������`��K�O8˖���3�ش6��Y��6>_�e�U$�0Im�4������!NM���\QSx]��~�>W�ݙ��.{驙m���ꋂ��\�LBh?u��A�8:�9ZƯPL���;٣%���m=�l�c�[֬�c�8gu�2pW��F�4ĳ̉���=r?�m���7?��I�D/�U��J���n�����LjAI��Ϳ���+W�&���ǩP�%�2�ҧ<6�T! L�^"mY��u+wbX�RT�7� �s�� -�"A�}��S�+g��Xl}�/�-W�<2창I𾂌&f�bx �!O�"���&/�L~O��֡e1v7�V��z�~G�|~�&".t�^Wψ�p׼8���ୌ )\]��ʏ�v��R�`Di�<�G�FsS Ylm�F�>�}9�{ ��-�Ȋq	��͘�uOuAr�DQ�cͺ��͓���h|�߻'f�נd��w��~a�=s-1��?P��L=�Y��h���F�1QZ
�<Y��6 ����)	!�v~4����m�\ȢL����ȵ&�~�W��j"��<�n��C  7���B/��ᦐ&�C�*d�VgQ_�Wk?+7T�2=KCx&�s�,�T�p�s�u�}�.Pӡ�ߩ[�zkr�o��C7��o�(���a@W^��@�	������Ud��G�#�^G���̆J�GHE|t��L42�`����w�@�m�'ȃ92�vFJeD�`�3�)�W3�ɰ�H�r��|,17M�E+����y:=k�Y&�D�	��`�0���	1�2��!����.*�p�0$�
5��M�l�b �\�s���QS��so,PJ�/H��<�K���}��)�A��*�x��+�ڋ�=���:��m*���Y�P����j�71�ТTm��+�:Vۀ�p�]S ��p����z��:�J�:�ޒZm�ҝ�~O��`��������!�_�[�}M�gC��a�f�Z���{#��`a��*��tI��m�א$�p�'b�Y�%V�+�h=�u
���"�´	�z}7A��obNk��O�^.6�sq=}�M�-�>r/
��K�31�!@��^u�(�k�w���2����fu"6i���� �_�S@�������q�i������i�F���q�lS,�}^��$��k�;/Oj4p̫ʁ30�I�O�k���K�)
t����O��Q�sǕY�ɕh��ʲ�Q��4��_��\�C��ht��4�K����B���ZM�ۜ|�|�����uQZ�T������զ��������Y&yK�k��X!)h�6�R��5ᤗѐ�K�����3x�����k�َ��b���4���M�r ��Xĝ�E�u��d��v���X���܏/WU#}��A�u��]Vo�i9Pk�`��O��ӵ����>%	��S�����}�x�Q��[$�-Q1k�8�捈��cT�}vV�u@јk�<)�2����:h�*�Y��n-��t��5�߁�u:JN�ƶ2�f�N��=!�ʵg�b Y!�-y1#)�Z��ŬW������w�ot�}���]�H��2�cHny�uU�ٓA�ڪ����}�L_\���VJ>�d4����h"C���
<)�M'M�oqRn2.��JUo` <�#�H�Y��G�Ѫ a�^�&!�I}z�g�:.?�[E���:ƍ�Y:��7��R6,�ʨ^O�M%��W&��(d�����h�����0�� �ߋb�L��~2~B �L+�X����ί���L6׀��p���$�ge�8�[�˯'% s�T��ؕ-J��'��$�R��2H�!��o��M�{	{��f�'���~pj�����	�v:HQ��q�7;7�}�*���&�dy��w�p�Z(����U��}W�
&)�DV@�s<6�������GԚ�X�<�k�<l��`
����Z�.RqU0�,�Goq�S�V�wvy7e��`��@>,�@��{�DdH��@��xf�m����)�o�z�)r�@����9�R^�&T�+���*�㍜���"������ipMl��L�>�.���6=�;��� ���w,0�&3��xu�>�k�T���~����s����֒�0V= Z�	64��j�4��M�t̀�$��.s�l��U�Dp�볬�O���_n�٬���P���#1/-ߏ�-Ҥ�X�+���7�
W��Z#<Iy?#����!�9I����;�������㍝Fo <�n�B����ny����|9	�������㖾ʮjz�MZ��S�ֿ7�xp	�������+����+h�Ug�D�һLJ�0OO��Y���s�t�َ彂��&I��6N:�,�1e�0L䢾��+G��$�8��?�U�MY���z�P앏<������2��Gb�>�D� A�
��FuS�;8+~�H\tc!�H��_�6�QL'�����߮k?Ѥ�[����&"B�XpwQ=W��s o�Ș�X�M6��_���f���8��p�垮hp0��O�ڹ}���:L���~��y�qE�� �Un������.0~8�p�����w���S�!0U<�r���B况���5�D�bm�~�.��ڭ�솕M!X-��󬣻�	�D%�e����;w��¾K'�Y4�#�chq��^��mVC����:�ݭp:�	ő�T�þ��Ķ]�G�K�X/ � ����r\*/"[e�]������z��ډWR�h�s ?4 O�Rmx�Z��&��A�bE�R�!�����äI�I�.���F�)Z��P�Y)�_�X�`
�s�}Iz+i�Q3s���>K�ٲ���y�p��}�0���-�Tz�-����4}[�V��H�OU�4��f��.���r^�x�K�W�;���>?Jv����� ;^��U�U}X���x�ј6�V�b8H%��>*�0ʒ�Q;��T��+I�����:x���x#��Q��vͯ��ٰ�~�ƛ����Ek�˛��6O.�v˨����!n���>�b{+d���ཌ-"��q���T�	�aBi}cA1Ah��Q���|ԬSo$J�Hw����D���!L�ul�ō�Cס�I�QЃ\4�
�:2D>�Bӕ�9����)��Õ ����h���U')K�ׯ�~R�ib�A3a\\^qo���̥��s|��+O1�Id�eWg��S'-Mtht�0��Ls���(o��U%6��֏��7��zM��4P�#�	S\��Q�i��E��L��g5M�&1�cx��&�n���)S���?p_5���;7B��wf�Ŗ ��V)��O�O�T0R)�E{qm�Re�Y�Oq4�:�~�k6~U,0���kh(�H�d��+ydtfc)�=є&�f�r�5�L���YHݴ~�P��?��i��W��`����zG�04ؖ�T͙b*G�7�tgzY��=I�G�*P�)X��	�Y,�/��jFqKZ X(kX���B�>��f���{�}C���x�-oH�;!�8�)��`QLZW=��t(��O�\��#�� ��_r%�IB��y9>���
b��GzJ�k)��8OM�@,1��}�F��r��}�v9Q�B�!2�I2F _�T$��=2�V$��Gx�l��� �
�S�A���_�J��Hip�f9����m�*
�o�+R��ܰ�J��##p�(�(Zvan�����_�FDQ��&�-����u,U!ȸ<�?���?����)�,��@�'������7)��_�Q,r�/ӌ�?YT�_�N`�A��S�Hw�p�0�sr��4b���@�f,�ʭ�
"��93�`�/�������0�7�C˫�O DE��Cɶ��i�ۧV/�D�/��u.����z�[?��o��n2ƹ�_���*��b�[��t�ɪ�Dw8LB^����ڠ��}�7>�$�����j扴�r>m���w���� ���R"�/s�������tH`��'r�ɲa�ǧ�%C˪���Z%͉�\���V�F�.����R��HZ���L�Y����/�"�fTl�a�e3��±U��@�:$���[�`o1�>�P5d>���/>
���VZ�x��	�x"��I���Wxu��^�燍���a�D�� _��i�a�e�c�p:��3c�G�R��2�BѪ��R��w���g��)�ه
$��\�KH ŮtjB[pL�'&y��J4�/	�`Z�7��H��[�/B)�q��6(�a�=hS��*Rҏn��7,l����eC�_��CK;>�k��}�esQU�U��֏�cA���2������o2�2'A�I690�fm�4���-!I�7��T�*w"Cv�(��0��c�4-��������h��,��FP�{{���Ee��Yhh�+/Zɫ���k������8�t���f��P:���,%�
�F����9�a�XFU�%M�N�77�~stl�W���/r�8����P�eM��~�2J��y�_*kP �߶�9�;���hm���J'��:_m��xe&��߬��v$��]�P?�F�@r�:Bf^[������H��A'eq��@��8�A�`���+���#Ҽ�[��rL�Bq��2z�Bi�7l����A�ܶ�!�-Q��+��~u��1�,���m5gBg]r#�T����<Cks`�"ݧS�����e�r*��R��7э	�k��\���-s���G�#��F��o�QN�lo;}���1�m�1l�\�-Y�y��M�*"�pѕ$�Z�1��4UbC]�����R�7'����k
զ��V��.�
�F�~�I�\��es�=s��O)_1Q��z���.[�t��Z��C78Ke��U޵7��}��h��]pY-/�߾ M�w,�98�V�ղ��Y�/�'3���_���E6��� ������:�,�����h��:E>b��^4�+\�с�e�ƪ%n�^��Kj[K�����u�}����ZC�����ټ$���7���<���R4�f7����H����n@+*g������J��e}�-��ۼ�9fs.�Y}>%I�0	]�\$R��vNN'��l[z��םM�X+��p}r���{i�p/�z��c������}E�_7K�^��J>�b�L�H6�7E����`ZAj���?�>y��ΐm�*@rc_F�����^,OR7���[�G�m=�S��Z!S0���%F@�ߺؕ���@=���cί�.�f�QnS�iX�����]fWi9�� ���Y��O��[�����̘��d�Ob�N�z��iU�a���HL.˫�:Hje�ӗ(\<������YCw�T� �a)��XU��4�e�V8>X�G�voz����=u�vqϝ�VJ�yԑVx���5����1��N�B�!3�����A��oT��ҿDLH�8y���=`j���W,yN��!�Ά�h� �q~�/T��|)�;����u{���?YkRz�g�[��>����I>�-[�Giȅ������{T�Y� *��*�%fx�<oO������ءf��i�u�U!��8l,e����"�e�àZBM��%��Wn�"ie3��&Vm#y�-o��b�/p�rï�kÐ���F�JH÷��M(Y�}���O%l�-�Ƚ5�z��}*�U9 �o�B��X;�OfW�n�'4�OM,޺l�$1��8�)B��t*�o,8��?��I�e��v�bW�g�8�����V�S`ى �񝌔��o���|��8|��E0[���)�Z78�ް��A�P.�ܚ��8O�1�$���q�aHZLn�@��@��k�!�O΋*�BGx�K4W.1���Kuq�#R?������ I�jq��~�e��	���׻N�U�����Qi���9�~߇�1���+�r�^"��br^oi����5��甆Z�����z�.���D��hK,޹�y��e<���ї�g gS�;U�t����⎈�]�"��8&�����h�H�3ֵD9�^W�OJ;����Wϋ����e�;��̏iA��@B�,M�Ю��L>�֑�d/| �q3����'��z�8����C��8:q-��4�� 2�;�)c� ����ܘ��s�+lm-�Bv�g��e9&.��}�Jp�����h�ܭQx����C�	�d��0�	|�5��c4�W7�I��[�S� Cs��վ ����N���P��-�Z;u��kd��6����|�x6i����~�o}�'��Lt���@,k�<�}v�n�@c���WI�<������<�*pS�4%�v�*�X�E���W!��*o�[�m<D��̓�t�X)P�+]X/7Y��x�Co0�&����ȭm���6�g�l����^� ��NdL�৲���)�H;D2޺�;Bjo�:S�B�&���0LS�BWF�ب�Arf�ǝ]�[���\¸��[^��g�����;��]�A��C��l=���l�"@���Q��2�9��R���;Ҧ����iE}�{��顃�o�v�k/Oa꾄�=�k���$�m�=�G`1܅tK1�4m�aHw�����.��AX�\̓��X.g\$gn0��VR�u)���0�����08~Z�N�3/���/�yXcd��Vj��͂�_6��߽if�cI���7�3�+\��F��]�<�W3cՄ��>j6���mGn�q�L�\'�w/����(b~꽎vSoW��3%2xry�k�a��r����N�7�@�'q��o4����0;���Χ������h���|��۴4�Ѡ 0ih�Q.��yA���.$�d�Y����o�Q�O�C�����6�_��U�P�@$5JI��I�X?���2P%p��|팳R#�H���l{ޜ��t�|/�v�c�w�HS)Z�w.K��p�dS�r�ϝ���c	�`�0�`>E��~�X�Փ�?�5N�Qf��ryi��,��Ẁ�v*+IK���ޡ�-�:S���?qz��$�R������ǋ�}N���=�6sP��Ax���0���7�8e�u���I�Н��G��q�`zE�C��)1��U�3K�.���s�_��t��Ӽ{8~���,k2�|3��3l�&J-x>v��ؑ���o@�x�o�vU�����ݿ��uJO�6�_;�|9>� 5�"'T�!�6R�M''�'�����`��	�f9�_���ܶ���+��ZG��	�IA� ��l�v�V�!��W��N�F�Ӹ��v�����Ĥ]l�^�@����&v��aj[l�I�]���]���ƶ�X����M���� �h*<w�)��~� �ޡb���b��>�q+�N�6�i�+�h�n�X�g~��.�&I3EW���QG@�Ms~�e׃����jҰ��̆�c����Bp�Qg�U�t!������ūX���א�mdĬ���b	QO:m|{���Q�
�]���5����|��j�(U� �S&�� ���$�Fo�W�.C�j������~ͨڴLX*�,��!u2�H���ω�-yS�@�ѭ�09s/��DA:׭+Ŷ´�olB���W�,q>���Sm�e=�R�ۋ| ��("����-YKikLV,A�oY������xr��O�!�%L�r�bC��۾o�B��Q�m�WݚƢG5.
բ����q��N�{x�M�Knz�e0#pc�bа�JH�i�%�|��Ԟ�O��,3�[��ۉ�,�XsL�Ol�x���
���cU��$�m�dݿ7t�7 �XÞ��@�|-�_��'&�1�f��bOR�/X�1�^�~��������;��ĳ�@����}2�fL��q��`G����5x͎)kmk�AJr*�*�O�RƓg�(Z&���Z뽰��)�]S��&Ibhls��1Q�W���I�H�,�W?o�ۨ0=MaL;k4�̣�����K��H�l7Tkv��/��j�;�xv���������l�5���>|����z�l��2?(�6g��Qp�"�H���`�����)��؆w&:�b����x\��|P!
�̈́�v#�Ҹz��48�pz�MA���tr��z8!�B2@Q%�M��7jP�>�)�/�Z��T�y_����;�E�'�La���S�x|oS�A~�_ؙ	H��z�H���{��z�u�ׇ(M;���J���Lc���}�&�5D��nv;���j�{�����`t�U���|/�}J8h��)�o���a���R���o���X� 1�����Bɪj�l��	�L�\���6�qԥ�ٴ�u���.&kkM�_�x/H�z��x� E��fo���<���2���н��ET����IV�w0O6�����}���������txb�d��q��]�*�kH� �ffH�i)�]Z���<bJ�dg"����=`G%y���w\�T��P����}�*e�Ҹ�b#�5��>��V��-Z�3��y�r�@����h`@<|3ds^ۋ�:h��Ts�ޥP���e&S��L�k�o�F?���x�e�]�6��<S_Q!���Q�#�Iѣ� ��yS��\I@�^}b2F4�k��(��7bq�e=l��#_J�w�g���9b��Z��֥� (�$^��S�Y�h�s�h�<�*&�SW�X�g�ӾQ��)�����I����� �Ô�;ɞf
�آ�>�/d7�	e3K�Jrg�b\��p݊�_��#N�Ŝ
�1-z�T�o�aT�XY���[߄�qE�Jz��������˼+��U�!�ѧ���<	���L�|�4^
��84�����:����N{��/׭{ ������
����V�~�R�RI�>�����r��xbv2�B.��6�>����t��Czh(Ys��F?��m����a�pw�P��n�9�@؜DѬG��H\+ç�)�L�VӰ�O���]c��e�/��i�ɉ����X���v«�����ZNY�7�5���yɸ��/�qb(�Ŗ�8j��-mD�wZ4g �RN��)�x
�Vp�z���4BFwpL�B(�]B��C��Y��^�+�\@���N�Ao%��R�<Rk�R>� H������8�r����p��H��.\D�>9��M?v{/p���x
�jk���T���P`�G+��u������i��&�~[��Я�n�r�S��Z��w�&I����i�EQ������-��e� 2=C�R�f���)ZMD�"X����7Ō�g4t��q��)�nx@w/�_4*UM���o�/�"�������dO�"1����`/dk��Ҙ�x��gc�ނ����W���%ǽLړ{�o�wa��Ă��fT����
,�@�]������3���8��>��&�~�x��k;<��.��|u�y��]�����2��B�&<�=j�"�:���}�����]������06��\�с����S��؇�%�2�j�05-X'Q��1۝p���u@�!�'��vp/Q�XR�)�<�FU̔H�� ��\��m�y�v$�ܭ!��h{O�,U:m#�?��>`m�	��92��`N1��J���EPT���5\�;+J��J�.iDː������W�v�`6�,D>�lO�����K����������7�I���Qp�ؼ���p:��%��H(�;�ֳs��{�7�;h��r��5����|(��������	\mJ���`��´8��:u�8֯�&v����
�ɀN$���$�����2�r�����^8�6�-%�c�W۩�����-Մ�Xdee�RUs,�P(PC�pW�~ɒ�������}f)�Y��t��Τ}��Z9L�$�iHw����x��4UhI���җ�`
�5o�2�/�ʬ|-$�ĳ�������Or:-a�̙|�;$�H���P�|���Ӻ{D�D�1�
���dP��\b��yi�������'��j�@G��uAt3��]y2?J4^fj�GɦFA�/#<Bj^��uOqA�g$�D%
�!�G��mә �9��D�k	����Oy.x�`����8ǀ�hi��Y�c��r8G�_$�q9�k���u�?4K��k'��Q٢)��-QM��Xg�G��������ϸ%g&�E��%�~��C��	pU
����Al�@����geZ�]�r��C�s�/F���;ͣ���)�8bl�ɽFݽ�`�"F����pzw��j�`e!&֗v�W$�ⶸC�IT�8��sø"�d�E�oD�wR��eL��{r
�+��F߾�6;���[�z,r�BQ�%֗*��B7
!M1�U��2��Kϥ�A��e�я}����N3"݇��5*5b.�d�j[#��A��^�H!�}B��"l:���>U2�/q�헎dl�9��.�����q6�����TPj��׷Hċ�Q6�pX`M\�R>,y�_d���,NU�
�h�&�T%E#,n� ͸
�j�x��O�-)�	� S�`kd�[� R����A7�	c��%��9�ۄ�.e�k(�N��t�Ð#ξ���,�a�PuE��H⾹bY�a�ċ�T!�N�M��%�vѳ+j��%�.�>�M�L��ׯl�\��\�I�p^�Έ��|T�U�"���CY3�z����gS䷫�Ք�m����uh����8��m���Ί������L2�~QK4I��?�π��f|��9��r�I�����Yu;*=N��t����fA�9!�p5O�y��>�w,/;q䌪�E,��ߛ:f�����ڪv�i�H��X`�ѷ�R]h�EE���E�W'�8�\)`Yo\t\_�&�ʳ5����nj��i�O������z`yL9E��S��`!a.^�\�(��m��S\mQ�jO��
�oB�ahy�S�x���{
���K \x�V��]��C}59f�%*�
V�iwLp��<���M��^h����ϓ��.L�e8���3��+C.�'�Y}�k9)���A����\[aD��0�q�#2?����1F ����|f���v"�5��K�
��w��c���c��s��c���x'>z���z��DZ$��0�x�|�XUЩ��n��	pX?�BQ����b2>�~�3�j�Ѱ�0.0�$�aؿC�oD�U]U�2�	��B�HG�-m�h�c�+�9�z|�N�Z��8�^MC�$������ٸ�N�֡��,���G��}d^�m��L�,�ܧ7T��R�@}?�%� �$=m�a�(�EL]%)7�ҡZM�S»	#�ХpX٠,G���0\MC��W�n��)b_���T�B��)���a��"�5LKy*ٻɚ�Y��yn�'�k
���&�����&�_��@�׀����Hlb��\��6l|��ݳytz���q�^I�6��x�N�w=t{�";�7�0�P����l�b�/���o-�X̽.G7�����;��+�A�z�9��>�>j'>� p�Ҕx)��ﲚ+k�w��]<s��sO�d�q�ea������hT�A�y��\���I���vRT��x��떝1	5v�Ί��|��2�ǠZ'��5&�RbL^)%���3M<�����}׹15���*��;�#	J/Ǎ�

x�n�t�!nc�K��y�(�S�Z����=�I]ڄ�
�B�c�OO�<^�u)g���eH���7ڍ�aP��mqM�2\�s�K"�a#���c``�2x�bv�Z��{}�5��d3�����T�� ƀ��VRϮv=�V���;�Ce�薬 ���>cZ��t]�3ɔ�ꥑ����M�w6h�
ý��:���8��\��q�-��hi�vc���S^���n��,����?�+��n�4�l�2>r;3�R"\")~|����T^eʜ�C�ۦp��!����e0'��Ko�Jp���Β?�����[ܽ�V���(X��lu�3����T��6�����u�j���V2V%t~�G,��M��E%����\��n��í�Wxu�<�y5�� �����ͮ�*OЖ�NR�QC��eg���u,��5R�*��Kt��7[�/��{��?f�o<����[�Ax6 ��~��g���-�8j*��Gt@Vp�~�[R��k�����P������o����r�����7K@�`����9�fɸ�>�Hc�1/$�a�,B���(��:��t��<gRJ����T��]N�{��P�Xʩ- ���.[�x�,0�ɑ?�^j�'�����G{�w@���MDU�a���P����K{�G�!p�3��(�J���Zc��� ��܌t���]�s�ۊU'pKQ'�������@��v3#�T��T�Ÿ#c�i~ �]��r�5�o8��,�D��Pf(k{?Zy�ˏ�c��7�)�mU%G���[Zϯ�,:���n69�O�e��ht�btu�jآ��Ǣ���d$J���������B��a�C���c�ɂ�a�����ĵ�,'���<�7���Y|=L%�bgo� D�	�<��bY��7�fr� d����ڮ>�H4eq��=- �2���Y�!vm��o��B�7�6�۲"W2�/=D�H}[�r��h<�)��R�'�|G�����c1��dND=�i$$��5�D�4Eq���^Y���6��
ڰ�����]���ގ'	-J�7� �Y�u��;4�����35����x���v��SO����#v�_�>'AS{*�F�vg`��t�[��xW	My�e�yǴ�t�d�����Q�m�p�4b�}2:�rE=@,_����K���N���P���Uې$�3:���$��v��(�Ѳ�}욆?Z�*q���ja��������r�o07dYi��$�4Q���Әw*�y`��[8�K��0L�Y����XP��Ļ�V?ގtZ�]��홯��t#�G�W)�1��33J%I[@��m�jsCI�S�!��|[��+\z�6��x^�=�������5D���]�o06��pOhW�6��zV��:����Ö�&V���kv���41�$,D�t�9J���{M��Q=�Z<�d�s~��}��~������舃!X&\��G�]�� ���m1����j��lγ�
������t;�c���OX���ɭq���[��XW#��)����\��HM�{`$m���e�N�h�C�	�0�fSG���_d9L��n�uW ���F����֔���D:�OÞ6} �]���	�j���psl�ꂐ�(��xHeYQ��v=W�����R�@�㱻����4�D����/�C�f�[B��U�`Z��C7��b~���ȧ�4�� ��	vÅ�}��1F��ѳu忀t����dG�� A�S/?��G�J*M(��EJ�= �"B�M?*�p�P�p���z��d���!> yfE%�V҇��+i�~{^ڹo�-Ņ>(��p��RomNh���C��X(��^m$|/���a�/Z޵�=7�t`�#uR��9�ۀ�E)L��2��v<M��\��_:HK��P�y�}�����O�}��r�ت�l�u+@w����H8g�Y�yM6�2z`,���\��뵇�,�]��X���V�vbC>�Y��5���XG�����$�Nr|V����ֵSŁ/Xn�j���wW&�g�N��ꠔQy�^PÝ��4e��5�������&p+�������a*��%�J���;b�e��O��!��	�հ�G�?;�JփW�-�����@w(i*B�����0^F�e!��A.ʈa��3>:�QG��?�Ѧ���%�5VC��w��Z��ь�0�!�yY�(xO�� v[���QWd1\��V̂R�˻�/^�a����#�?��(5#��pBr��O�H��\n]{����,X\]r\K��z{�����{�y���*m����t�t�p&�y���#"D���^�!oL&�|�K�c`���k�� ��*m���I�W��d����Oy����)��lk(Z��?���Ѱd�o�ǫ:�E�Ơ�XCu�(�_\���)-vĬ5V�W�*$��P�E���=-?Le������W��S���bL=�l���r���ۆ�?:�sCT�}�8�z|s��B�����a�Fgn�<g�5)��:�*��Г�A���tf��C/�Z�.�K>���U~�d%��J�]m���b��5�TӒ}�-�E�Љꫧ��?Τ�틏"�,��Ġ��y�o�<��cDa��[X�sJ��Cs����W���b���=�АL�!(�����!�a�`.�9n���U�?��~�O+��v��Q�YnHvb?K�c�H����R����%M��#�]�h��̏���"˃TE\�r��<���6~�4���kR���Z���KU!O��P���zV������TFʉ�bʽ�,�cv-AـG�����V�%?m��cO���n@ۧ� �����,/�J�\����d����	�+�9�H���u>�B�ɘ�vm3��)���V{`��2�p�aQx%Cc���S��I�t����S��J�r|q��d�f�(�ņu���~5��<��[yxX�c�XnA��&�=�5Dǐ�E��!���zG���#i�H@hQf�-�d�۩ͥ�3b�IM��6b�㺹��������ԈSV��lH�.;~;���d$haj5^��Gf���?)�Ӫ��ͦςh�?�8���â�g2�s���,,8+�* ����L�~����2CQ�\F�Y��.�u�Y��a+;S�����& �h(��lΝz-u$��3>*<���M�(�[C<yw�C�� �B�{��.�	I�61օ>B�����t��U�Ɨ���r��+>9rB��)vO�>��Wj��Z�n�)k�no3����'�f$���Ձ@H���"�u�@�R�EɆG��"���A�؉ez�n�z�<�����>��^��'�%n61vL�l�ɕTU��4�Er�4�/5�ud��9�$sK��Q�	�3GO8g5��-r�Q��Mi������v�
!q�\���/�3�;~2�Kc֌O͆q8:1G1hI�:�Iz����l`��D�R//��vM2�8dGg��։�߹P��l��'.a<��R�o���a%g�!s�?��6jaGƤ����"��DC܃��^w��+c��LP|;�K�n�*˅2.u���V,�G���?a-LSB2e�$ߏ��wU?hp�nL��q��իH��Ľ���I�O��xPKL�z��Ȃ�|�ݕ����F�x��I':����`�����<i$9B?!v�;JS;��#cF��(�-!m*��q�t~��������{��X���������"���q�
�B2Wa�>@���)�\��eN w֔��/"����{f�ؑ{=��>��v���1ӳ�!2������*�'S�W���~�]�:�Z�M��ԕF�·����ky�+�6܎������f���\�j��P����nsy�3��+��������X(������b6յb�vf��Z��F~� �J����aA��[3����8�f���ڎ�v�m'"5ݜ�9q��\w!�q��.��	啠y��j�B]���$:_�,�ǚo����[�|���8��V�
�j��>̪��/!�w����A-�ɿ�g���?dGI
�.糨�9��.�k��y�B�Y��;�o�d��O�Z���X�]˦��9�{Z��#���J�(ɣ]3��6�}U�6P[�8:2E+Z��1˚�,�,��VZ\�i$-�$Ѝ�=�Tײ}��
��:��6�E��_��c��IU�<�B�[�øV��qe��}s:����>O�p�Kd��&E�t�>M�O�<GBNZ��M,J*�Gx�ǮO�e$Z1�W^�Nc�x��*:�I^\�0��
uѺ���eN��R"�!���gy�HbE��=M�b��l�1��p�oM��+����h��->��^�M�/m�^k4L���C>�	fC&�8&�R�h�z8�'el�{3�A��D������r�Lj�{e�~. 2}�`V3�0N9J�-v��Q߯_G������y�N�A�c�:F\cb:��c&c�����V�3t�>��m��� "��"y��l�q�C6�;T��I�y|O3�c�F��Y���w��O�H�}���hꈓ{q��0�]I�^���cø�"��*$1�?�:�Ka I�ÐN�0���a#ũ�IJ�$��$N�v�Ăb[�ǡtl�Q�^0`7��+u�I{y?�����e� /��G�W���l��\B�	����pί,Y}�m���:��䏻��z��cq��l����&����b��&\�q�ܣ5����C�ܖd�d#�.�H_��s4 ��W�U�.P:4jk���k��y^�ݳRt�+�𜋕d��@y��`cT%x#�GU��QX��2�8�=w4D���Fz�nG��#��;쇇A���ZF�ܴ\�~����<������)����:�7��)4&J�ȅ5*�u�0IZ�#rI��D�:,�Y/��ħ;���E�0l��vRB�p�/�A*b~�4ruf�:
�U� =$�G��M�q��{$L.�2rl�AwhY6dr�f��co��J�q̞�ԲOn��MO�KP��W$:�n!�V�j}�r��f�d1J�V]��p0/���J#|���G��p�zڤZEg��t,�FJ a�������5�n��L�4	^Po��ˑ���H?���%'E_�P����l��D#]�`�Տ����9ρ���3�g~�:���g_�[c��K��*���ح;D_�)���N;�ұ�u��a��h�&q�ή��*x :�*5�-����Ƿ��W9�$.�,�K��d�N�=��J��e���r/XY#u��8U��ʢ�a5:)el�9�z��	I������$v�S�����,yT�v���%Ʒd�6�Y���Q�A�?����K�;��Rm8`q�ƖU��*��,��fD���u��6ZI/���Ñ��秃G�>n9?.��".�2�� ��1}{&o�e�&������M��r��Sj�'���5"�)e�`9��t�ㄅl���դ o�tu䘀�eQ?.�a���%G�k)E��p��{ �����X��$ċ��T\K����Y	�M2�iz��#�~��"��X7g���@���Q�w�����^ܨr�6��vZ�s�'0���ŷ0�j��r�9a���GeS��/�È#뻋{�,�{�x�RJ�%��S�e�Ñ���,=J�b=>0�+-.�]l�H�ߝk�k��"@1���g�6��M��j7�u�2k�m���@�M��d1� lK��	��i>�1���	s�ݝ
���O��`6� ��(Ė���l�p����w(�����סz��+����>T�v��4��E����Ne�r��合ѩ�وOO�P�ʸ�OSD߀I��o�R��UZ�dޑ�S���1.��)�����qW��/>w�Q��IƔ��T�kR���Ӝ���d�G�TVL%��38._����� ����Q�U�@��k����k�i�c��d�[{��ׁ����q�R��>*��[&w[#?h��`cv�1&�	�C�j:�z��~�ù��n�7xre�\��k���**-�"�d�mZ��uu��E��aŃ7�Jc�ʹ@Y�p��r�]6N3>��񜎚�J���zw��f�p�BE6�
�e]ɻ $ W� \4�9.�%�H�J�(�ɾ��Z�e�������7@9q��j+��˃���g��8h��t���O���j.��ۋE��j��|�4_���X���njy���!���o*1���Q�d���֟��t���;� �u\�]08���:M_I�!���5��2���~�-� �D�Z��~v�G<j�;�/�ƝPD	��hy�ϓ����Ԥ_� �����k�T��0��N�ţ �fi�W8��.w�mmϑ1\�:�	�B��ɨH�m�ٹ_��s�oqX�$�O3=�X�'���!�*^�AV�h�D��zH�!z:�	���Z�q1	��ϗ���t`���jȰ0#h�a�ș� �1�����'�މ�n�l�eQ|���Ϋ�ъ	��Ik����f3����!��u�u��!���v|�,��F	�r���\�J�	�JI$�+דm�;��GS�V�}�6C�>�Ӗ@��
��+��fc�w`:��,Vi-��!��|���D;Z��\'���5�W�F�$��AB�E��2|���s�;��[���M�>��T�,׳��a0��.�}P.B��|ۊ&n�7��2OE�F mh�Xh$�?�-�U�7�)O������(�jZ����g4R��{<0Ž�Zb��@o8,�.�X���6.�!�4��<zZ�==@q� 3���.P��r=xzA�Z[�0E�
\`̒MFq��" /��zi�J[���܊��B!P��򱄻ܥD��`Fk{�܏g�K�at�\ ʕ��{V!,o+��dD��K
����[ݒ�-�tpđ> �p.խ2�Xx{�֔����2j�֓�����̷�ZW����bޅ�F^�I�
^�ޏ��T2Mw��l��)ix���߯�1��?"l���������i��X������l�s �c ���J���l��I�j�5�SR���DյmDCu2�Jq}{>��.��O�/�a��3��׍��Ů̖K���:�p��U�FW�q4�~�I��Ƴ�����99��u�3X��O$�(����q�ƃ ̻��8�� ZFg�s:\���` ;�*o<i�̓kB��;�*����B)z�Lv�a��Oɼ=Y0������F����g�xÁ�:�J��i��x���W	�I���% P�}PZ��\)��3��}+�'2���e#�k�������l%�0ʯ�дe<��"e@�2�!+�tt��V��B'	Q�Kyf\o�;eX�;�5�u��N5�����/�L��j������T$���1����Jb{<���2�_-��?{c����>tR3�X87���k�ҰpVLH*�c�A��A�#�;S�>�<v
�0̄�i��jș�o��K�x�B*<����Y2��{g!��*�p�v��ܜm$<p�-�7<M,tq3��'����f�nN���*��^ \�U~?�i���%��(���~�r��Rd`e�.�T���Ʃ����WKA�"/֕2$��&ͶZ��Upw���A7KXҼ�3��ҙw��������s�B�KI�p���P�����P��@˗G�י�}��1&2�jߥ�jÈ�U�C3��/���8^ ���3\�R"���R����ZM�5��P/������Wk4ҏ�%�Z0� ^�]y#��;07$��f����!ž3zTbHw}Mﲅ*�磐*y�c� �@;+~��=���&9����E�һ��L�KV���Q��3�gSӾ�4��Q��ā~9�\4�h�SCzWޘ1y�h�>"�aR�Ϳ.���?�wZOa��4`9��1��_0fY�Z�k�u�����#�3QB��b�RT`$�m"҆���gOʩ
c�0.�.��j��+w��h:��m� �3����Q�үgF��aF�c��N����*"9?.�]�P`�Ղ��T,۾������&;��i]���Mp��xib%�
�(x����	�]M��Sn�����S�%�JnqZ�G�~�[e#�S��;gB<	^��z������_��!GC!�OSp�VN�0��⡚��9ї��Bl��pѪ0gFI�+<��S�K�N��e^vG�8
o{��3>Q9 �bq�f���ng����]�w�t������ ��1�d��.�c����䮓������>X�� {�2�`B'2��s:$X��
�@������!���S@���`�Y�3[ ��U�oD�~Ů��UԜ|�����H��@	QK����)�����8�	Яh��|����Kv$�G�ѓ|�訏���>wb�l�5��^��7g�hQIϔ��EРE�7o7�8�����)k��\�58���#Q���S�!5�h�>����E�j;횖�m!���#��I��_1l1��A;���H�kJp�PP�T�(JE�׻����.��P������)�v�9=G��i��"���v��<��<~5��]�e0�J^�2���^�J�_�tY��v��UA2hsa6����B�=f�v϶��Y)�cLJ�u�,,e4=3,�S�>�.Ws�I�5̬Ұ�}ʱ+5�}1�O�E���%�1_�6ĳ����B�Fb,��Z6��O̫�Jh��:4��(M�$�8̂��!�$��P.�H!�r�݋��%����V��C�޵`�r��?o�G�ʥI��2:�y�d��x��V�SM>l�Cx�a@ ��c$+�ȑ�$11�Xq�l�A>�"{C�B`B�&%���+-Ƒ�D9L�����T�1��4��~�o|��)VF�6i���-I�.3]��g�C=��,�o k3�8_<��3����D�`V�It�2�Ԕ��|5�i��3�x�F4}�� �ҿ>A�Vk�AFu���R6���#����L\��֐ <XŪ�r< jϡ�Q�a���;��'l�e's	(��M�5[��qo��Gs�[�j� ӊ�[p�26�/ɝ%�M
ނ"}�ګaM�j��!vb<��8aA���	����)� ��$���7�*a�&�e�|�I����;l᦯�J�Y.R��C\�4S�`��{�O�*(Z\��gH�i�^�`�hYT~O���P}!'Į�Q��\�r���L��(�����]�(U7�v����(�݂���C�=߼.����zMs,��x��%PFaܳ/wJ�|圽4�j�J��y06s���Yv�����>9<Ӣ6����c}��YH�@ۖ�,�oW0��[Xf~-sS���Eb2�O�gr���KX���;\�A�g��}�Z=�s&R��r��Z�D�zEo�V�m����̅V��Į/u�;�ϟ���&-S6	.$+�6)ɋ}��on�!��U���^���O��� ����6a��"G	���!)��UX`���3|�}w}l5�'���x�^ha�G�]Au:֍�g���J;���	���NN{�,�o{�L��݇@-
z��$n�v��sg���y�9��H��F����ʒ{��_ġ�� R������G�'�2�m�K6nȍK�w�r����s��Qe76!��>��{�Bt�>���T�3�3"�f	�O�R����Y��/M,�Ba�$�卟M�����A�'�C���C������,�V���}ᢚ%(�F}�{���C-�
�?ǝ�a�ʹ���P��vm^faa,�b�'`)G�M���K^ux��\���l��:&rK҉�O�K���W8V���M;p�a�ssW��B��H����]W���Fj���.�dd�浴v,��N�qnj��[\&"!�ҭ��[	F-��gl�[����
�'��Ltl8�6s$���v�Y��e  �(�lD��Ʋ���*F�d�5X�78�Df�����4f
��=1��4BH\Ādr����n2�� ��c2_\��P��sf�	����@yYk���s:���jc�M���^��W떚�
:.%�|�)G�&��&$��:��Jc�5?٠D�D�9%���R��uC�&��$��y��&-Zw���-z��c�$���OȻ՚R�3_u�!����✙���,��]T���}^.�@]�'<�+=���t:�EY�]p��ٗ`=�r��׎܇�n�$Օ D$;G��\r��ǵv��}���!�*O�lx3��C��&�x_=��, ��;4A��J7-��:?ô䮻��ӏ�#Z����]�t%�4Py݄DT!����92���\����bJ���� ����݈��Z˼g�(�,��T{U1!!�]�Лr�9�'�����B���2���)*�E|�p:��蔆�M>`/$t1����<|�\�#K�	R�!��e�������v.�톶i��OCع���^�C_?��n�S,z8�X:��Q�F��q���QBTiX\~��a��̻DJ�lŬ"Պ�����8�d���JR���K��A����"R
���D�ߍ�:9�e2�Z�A��zM�)M�w�Ȋ�]~nŁ!V�q�L�;���"�A����6J�\�F��wj@�M���l���^M\�o�^�TI�5�}�U~O���b���:���4��� G������h��6�&4��h�L����3������l.�D�b���j�/���4kۡ�P�.B�m�>u�C<��
CNw|z�Df�/�g�N��flxI�������A$��"6��U�Q55jI�Ӎ�Mi�Ic��B7њU;G&�6����0u����֦�s��n3�~��F{�1�O/�Kb���n��3@Ufy?��p�n:�a���N��B���a"xH����(ҍS���K?���x~��y��ك�S��= ���+PxN�!q�OpH�$�rN ��hB(b�<S^�#����N�
�ܤ���ٷC%Qؔ�MR�����)5q����a�⛄���ȥ/�ڨL�/U�5:�+>
�A��v��s�8�Fi����}}�[��Ҵ#8o�y�>��7z�th��w5� ���c�?�Mq�ʼ�;�?�C�{0�`t��'E�m���-?}I�V]�1d�П�{3�wk��ihNЭ������«D��x.��'r��69:��6�)l���o:��_rS)�C��;f]���A�j�AA�x`
�C���ȹx&]���XH��nS�^:�=���U ��]���K��(�����L���0B��J�~��`4䘐�D��|UOa�����vu��B"�,�!��Թ���D]�6E�����汼&�}!��6"�����[��0h4�$N�^���w8���#��#0c�f'��[z���7����1��hH��xV�X-zMM-��)T��㘡R��$�s�R�}�gdO'6�TN���K� r��QG�@9��k�K( �8�"�k�9�7	�p��i�Չ�~ܕ���`H=+�ۡ�?�������yB����F�Xtk4[�'}��O��!-M&��Q,uW<���{TcW.�[�?
�j0P	�C@���O׺�Gu}3%;����HFM|dC�$��F����w[�Wb�iO�p��A�7���MK�l�˪����J�ĝzr�J]m�0u4�(��`�ҍǠ4�-���1-Q ���>�7!�����������ΗYǎh���ԹFF��b�f+^��y?I��֣��s�(��~�b�~���`QB��?�p*������"z�}�)��~XG�B�����u����֬7�BhϞb[�!��AЅ��f��V�i�'�����S4ؠ�+�zV(���y-���]@ɂ�uߋ]����j��}�I�7T���#h���77c��Q|�O�o���`"�b��<��U;�b�5N�����>�H�ʭ�+r:� }��|�4��Z(��^��u�m����DE��	]��Q ��6_By��K��T�42h�nD�=���;%��F��� ����[��������Nլ�w�{�@I_@*E9W�<�J��z?���ܔ�H�< f�.�#Lz�2��s�ݑ�	�n!�f{�xM��P��n{Hm�jh[�1dm6�p�`c6�
e��}�<� 㓷�	��:\��bN��~|�'e+���j�D�$5	KH����H͈ ��*՘�s���#s���V���m���t�G�8��Z����y.U�O�8�n�6?N'(�by�H0��m��$�)v�Cn���z@��['�R��-��E۵� �+��j�mKh|�=B���7��oЯ^G�y�E�e����㻖�ؗ��d�ڻ>��g�M��˻K�K��Z	Y�~��I� r�AU�V��z!�Y�e��������dL����W��B�m�k�ǘ0��UB6=5���Wkԋ5�o�;Gw�E8��	�K�--j|b4v��Suy��!�Z�ZfO��}��q�r�DT��Љ'��y	����*KѮ�vB�Y�lN�����s��@c�6������w8��-`0>1�tP�c��v�i��0�N�����l,`���ִ�
�#�Mp�h�1����g�/�_�؝�wh)fN�g��������,�-�*?�h�� )�r�|�SP	2���w�5 @ڝ��q�͜���a��?����kL�׳�1}���
i1��~������|��V�B�c<��M�U�O`�[�N���gʮ�^]�� n) 
��`5�Z�Vr�u��e;�lm���֌�t��(�m�&��9ygN`����ّ!E~�J�1.��J��`"2��5��kk�mu�z�d]��u�ǖ�,Á����h|*����2�C5.��/=Q��KC��d�&Z8���K�����o� �_� W��G�nk2���pQ,��C��KK�6�"��=������Z�\w�(8�B�r�d�h ���sd���ʤA{+�-@o<��k��ړ
�,EM����x�����Y1 W���[/؋�{pk��<E�8��g��w�&�?J�"�د[�wfx����� �՝��������}��
��HN�D�q�9j�ʣ"�)X&J��5O~�S����P8@�g�e��\�N���iKEkV�F�;��N+���TЮ���Zi�Y�TQ���x���N^�(0���@�r14������%��eq9�Y�*����oq:��\�N
C��0�-j��c�)��̗�_wܖ��nV2�]j]n6�xy8�ˢ�NűA�u|� zY:�叙<ʩ��ПN�`6^������BL��'��v1�l��#�YD(��<U5 ���d[�ĕS�#Q���x�O�m�!��,�#R}��c}��������yޛc�뗧�&MT48F!5J�i@P�^Î�P�fKk�Z�	0~���H�5�>xw�f�g;3�W���䌍������:f�rS�'Tl���ƜZ$Df�����Y��)%_E��_L@�B{֢n��A{�ٙt�f�6��R]5�)Ll_����ӹq,��U2(��A�o�i�z�x|��l$���V��̰���5��_�?��:�V�_ۛn�m@^�~)��>x��AZ�YX���.a�a >�`���gNM�X��Rp�9��G�ָ���84�͒�8����@��m�	��m�2Ǉ�n�)��]Ξ��霹�2b�:�K��ޏOⰰ�CY&�Ťgd��27�]��I<�M�\b��hlwε���l �|�Z���1$K����Ӫ��Ny����$����)8gDD!+��i4�NL�M��r�j�����<Q��lc�ė����im�f-c����`r_�h��$-�ƹE�F)�*���� ��E�`.��m�C|ԛ�����:0X��FTD� �<,}l�/�^[�X;q�|Ǒ%z�L��K��(�
SNM7�����PA^�7���]{�ӝ��XR�A��Rm�sWU�������wgdr���k�&E���;W>s��?�xqg"���q��\+9�o�D���2Q+�g�&bW�4�N� �@�BU���FJ瘚>E?̋����iN�m`����ڦg�מ�g��φ�ܬp|�X����t��tO�L��D>���*:Vq�0���*�'�P���������6&LV��xb5_�sEQ1}�%g2���n=�N{�Ð �� �;�~̄ȠHS/6 2��^�ҀO4�}Ch=�!��%�?������^�`pU(�8�t��3~t�h��)��ܳ菤)����r�l�����ݒ�7Qgv٢4t����
�R�&�I��-N�?�J��;���>��6 ���Y��_5=�(_[S�h��$�8�2�놙@}�o���z�ŧdbQ�`�������I ���i��z����/��a��(p̍��ۊU�c%�XaVu�vx{���ȋ<x�����s�>��U��LYIL �}�}��
��W/�f�dD�w��澰H�����4�, �A��ߔɄF�����.�xJ�">0<$��y�=�(z���ȇw\ar��3]E@+`���7&�����)1�]a�rf�X6�pN��5�\~*i�3��~+3��wB`����$Trm�yHp�bƩ��0�<#�Lf�aoRL����)+��C����\3���Q�)�uݠ�����iFq�uW� ����x�VJD=����g??K�9��u�9�Q�J!�&o;|�v+�WȽ��M�`�'�1��+�Ncᜳ{{O�D�s�D�3Ρ�]��S-��g&��=.�wG	v�n+I5�?7#�/���o��D?Y�N�*��g���>���N8�ZS~�L���;��gg�O9���e�l��h��A�q���������R��������pP7��}}m1a�E��xV�։��F�ۃ�eF�bbr���@l$� �Tgl橢�}��1�S O�;X�-5R���������q��é��k�5������{V�ZQPeP)�����ʣ��v]�S�%x����R��E�ER�XS���9/�{�8z'l��-��=���_���X⟨6Z~��ҷ�(�ϸ��dC0ew4-��䠸��Mf�[.S(P���<r���}�~.%�����d���Yg��|P���h@dl�o#�]:���,�ڑs\���O6[��}�9!��L�g������4����X7K����Q������ty��ŏYk�����4�#��4Ge�C������[ZjCi����p�k���(�$�'�F��E�SHj�v�B8��
�)@���((�4����\��NEn�%Yp�:+�Φ��Y���^t#�����1sZ�#`?���ϣ���V�5��T(`�I�!�*1V��v6�u����[�����/sBl����A{�h���2�e�R`:����a�0�<'��*9Ω��v#������el0�5� .�� �U=�O��r�X>���3�����apk���>~�N�j7��,�^��k�Z E������B��]���E?�[S:�5�N!8�mQή������LAj�z���mY�P3{�[0Hc ��O*�A�ud1��݌�qT��m����U��y+�X��į�6�/���G��V����<�А�b��򗨄{��W���֙�Z��	���~C8�d��80���>���^z|���y)$�m-]�zE��~�a3]��QvcǍn����ߍM�N�u	C���������@=��|�a�T�_�6��SX�j�_�N�Vo"���@Y<���>� 69 ^���e{�l��q<_s�w������ҹ/IG�V2K������VV�n�U��3R���aU'��%���N��[q���r�Nq�KR!MӤ����t��d���sq�����3�	3�������������s��|*��6'E�<�4;�a���A��)�Y7V{ '�'R�J̶��K��д!�٤O�h<~|{JO)�D�؛k`F�?~�	�@��z}"D|A4\�Fx��Ӊ�D��|��L�;GN_}oj檿�u_V�í�]��$�$������1��ЦlPhs&� @�&�Yy�\yo�ưȨ�)0�����9/�����D�˛H��K��떪�~ Z� ��%�a{�% E�W��T<��u\�f7��FqU��np��K����7���������O����r�T��0ԑ@d �%(�U��M�JU��J/|�mD���5=;۫�y ���i9I�mhW��M��-
�v3�ʉ?�;Hu �PR�b�sE�oD�s�s?�ďӣ�?��j�4���_^��I�v^{�K�t�uߟ>�cHy��I�qb��<������?�=�A�!J�h�Ӏ}�2?��ϒ�9w�(�ѰCS������� ���������o���K\�����M��%����0M�F��BC�2J2��.���r�{�8W�(�K�`7��m�c2P��P�ժ}��+;�:�!����V�*�T��-���zq�"��ʠ)�m�YSy����=�;��C�_G���܉��_��;�-����DI�*�zm �����L߾oQ��`,������p��[Q �GA���ą���9-��L�[&����3#��;�G]v��#��&cW�����m�]���G�a3
7; r�h�(�d��ZuӉ5q-r� �e�sm��F3�h�����c!K0����{ f<�i�^=@�ށ��xXt��U=^�ed�iE���I����S�56����X&�w�&/6'���"+���ʌ(�s��B;�'Q^*4�mU���w^��sUO_�%j�����f���%vR 
�L.��k��X��o���_$}���� ϖ�Mn1it5�+�	Hg�`���~xՉo��Z�Y驢�g袲�S��=�VެHՑ�|'-s
���C�~�����D�;��vA_7�'�$�ݟDvK�f>7Ǘ'#��Y�n�K��.NzJ��E�욼_!��"��痱2�"����;%+ϊ���+��:�ݥ�H@��{P(J1cU"��~Lxw�d��sQ#����ͦ��H�R�/�7���0�P������R3����>�s�r ��~���8t�3$.����b�b9) �?�o�:"��bk.ne
�����U��AC�|�$c��D�Y�p*쩖K��{纁xzr�?W�q�`��$�9#�\��)��6[,���X|q��o��ڤ�6��=��0|#)�;g ��V 7�o�U�#=�l�vm�*ǩ���ç��?�S#UaB��fA��o��	8����r[�[p��V?��]ĺ��bUҶ��pܘ��8�ϧo����&�R���m�]i��®u�z��Wh���h�P�9�}�gw�^A�3�\|!ҥX_ȫ��Ws�0\�*	Վ�C���\�vk��O��IX���M�V��F���Gm:�ݐ�w>��\Y���^<�ƩӲ/��xܩ�������J[##uc�y�m׏�LCP<U�7�'g$���wt���X�+���hs	�nە�Kh�[�7p����1Ģ\"*��u�A�J=@��kij�� �=ʊ��>
�I���Ѽ�΃�3��~._�m���\-q�P�������g��/Ln�M�ܝ���#��U"���jc�G�Wu�iRj�;0A~ޛ-kF~i�/l�n>\���
�H�Ś*5�x\u��C;x���wհF�C"�7�6�Y�k�#�qg��Ν��i���,[�S7�C��8�i�uC�s���O͉�}bL��{�;R������h�@�w�J4)	ȹL6���ʯ�7�T�q���Y����Ъ�-�:�Yb:�at�����|GČ�V�_�(ӎñj��Y�^��uL�=J�d0�������Ϋ�ɂ�cA�U���JI�6�"��:��L� ��*��Y��T^2�M���v�7_,���A�a�'z2{��8���:�2�[p=��0R�#K�c]�`��?T8��6ɮޡ���֣.^\��(�v���&�`��4:,1��Dؖƍ�j	�1G�*�ư�7�q���!$��������3�i�	�L����fkE�i�q�U�.֡��Cv� 4	F��
�Զ��k 5�]�S�q�U���Fe����6���v���F��9�.l��ĨH��l�O����Qw�G��_CS:襙v���j�?�2y�ɸ̸�K.�t-Cê?� ��&�7K���p�OY�	TCXڗT��_�E�%��ѿ��Hu�o^�'�X�q��+���/� .��/ �#n40�O�:Y0`��S�9����Xj|�F�?�P�i�����=0>�.��*��%sI�J�g(:�"c�h��ug$1ɬ�Ym�j����*!����d�FGt������A����/N�:�e;
��zĎ*Icv�+��l���7V��$�xW��"��0%���c����+ r�kZ�y�L�|t�-X	��݃~��7]cY圹�ӧl.��0��������}:�9�x'P'�L�tx^|��*�>ɫ9��@�l���b�)ˠEF�� �y�g���܆�#�o~�~�ד�<��S��Ĥ"�1p��ؽ$W�[����']5\�p�T��"6�
5�0PJYѨ�3����$�$��g�p�
`�T����i'Ih�_w���Jt�'|�U�Ã�F�׉�msCg�2�;�b��2�[��L�P` d��v�?˵d�2Ҵ����9^NF�?{i�H*�_��|p�� �Z�xUs-j����ͷr�m��4���w�S��U��=No$pB����n����WGT�H؂�~�.��uX�"���+����(�@�,�D��oےX���>���� F�|�q;�C�;�2�p���v�Le�]�g��],���=!Q��R"�\��3�Ua�=�fg�=/�^W�p���oT N����nZ�0����{E���`����mX�f4[��IO�do���x����j?�m�7?ټ�R#���7��f?�Y�W"lѲֽH�|���_��0�4�E�|H�
���=��s����(��l\���Ű�؊��$�U�3��
JRx^��.�1��k��m',��2��jw�2}�A���#a�?oL���ˏ��:B#oUG���$W�Y�����х��v�C�Ś	��N	@��ca��xO����b--/U���Q��T?��k�Q �<ݗ��E��q��*#����������E8�[j �墭���V	�����`q�º�$��u@��N���w5�]<�x��DV�;�4d;��) -�6�k�V"�7�#����S���AqX�_^�7��s�U��Τ��E�Ӫ��.�? ՝Tۉl_,֯�X���<Da T%�&�����O�n�
8���d�%O�����åg���h#2�͏_�)�3d��� ݈�kٮ*�)0_�3��9�����;H���l����Y�!bB7�f�i.��`US���@�OB6�|�A�4�!tW�^��d ^+`�&��M磎��tK�J7I���]_�����-S�v�+z��D��7a���S�n�VL�+F4�o�X��[ty�A��j�,>K��[&�X�>�����,b���;���<�ˢ�KQ��{qJhˏ��yT<�}���ÏYZ�P��i��Cm�i0�����dMzR�ɰ
%2	&��P��!��� � ;~�������z�mV��?"����ɟ�6������_�0��yF�-�I�g+�~h�Q���D����nZ�lᛂ���!�4k���o�4�Z������Sx�v��*~g� Z((�
C�Z"������
 `�VS�= �`�kܷ��� ��o~�QK]���[^ !�,�`Z����F�;�v���^���v�����˾ضG=:�z2�.\�^V��t�$�@ �τxѲ���x_�["�������.�<��|}"lf� ����B�,B�F��ef}�a6�H�o�!>@#Z}�՝j���9� �&Z1�����T����YR9r e�/�jr�󁅼@�ã���S�d�d�?x�"�2����_Z��@L��:X�.����l��զ4��?�~��֢��8y��ܾ�J�����	�׏  �@Z>�n8�1@,i���g��1�]����߇��^�#G��U��F�=�,Q�nfc0�Lb��t(q��]�o�?��?
,�� �ᴹ��� �n.9[���R���#h����]�ū !�#CMp�b"rV?ͯP����=ކ�8��H�n�&g��oX��g�J���]T����� n	ؓ
�~�ݬs��$�a���4Ҿ<`Y�����sMu����Wʑ;�$�Va1�\]pi��\&l�W��;�!��`�V/5?��Po�|	*�����?6&5�C�n�b�䄎/s���!��1p5���q�LJ��a��pЏ���^\G�V�eET~&i�p��t�_���轷��h�N�];<�w�Ǎx*��"I�{.0���[��Z�2�|�L�l��X����4ԋ��K\��1���=�5����#�}���r��ǚM��Dd��ҶU���P���m���r�bYV���γ���,�������h�d��\������kҡ?��Y�͵�'v��)T��Xه٦��^��;�^ޟ��{����5�&n��>dÝ����	f�
�钷�D��*�}�;�*�6ʩ�a�e��+�����%���γd$�:
-�"`k/��D�h6�7�J8Ju=�عJqnL�%0����l[���lɀ�p7m0[�TB�c��R�As��.��n��5��y4�) ��6��2�H����H��j��,��21����dŨ2?m	~5�y�L�f����������|��v y���R����T����	��{��fyE� Kz\�y6B���dN�bu�)�Ak��It�)�F��yN��J%�l���r7SG<Ҹe��-aϣ~��8���&�P��ӗ�*v�I��F�g*���3#���%2���-����ơ8O/F�(�N�.����}��e��k]����ҭ�,Q�iR��FXݤ��(ơ\�XHZ"҃�M�5��lc�,�tr�dg��~PS��	��B\rb�&���T��;�^4F����Y�-W������FzEԯ ��*���2ļ-}Zjn��g;%t�5�v��m	�3e\gEa�����"gNv�-�]LS�̘�_��!A�����$���:G���~�tіf�����:��Suͺ��';�ޚJt}�N�_�t��Zޓ���+��Q���-�X�fD��T&Aҋ(�5M�I[g�"���es@t���lQ�u�ܫ�a��n�6'�6ج�;��fQ�� ����ޥ��$��]0�m4����8 guZڈ>w7	�<|�:0�g�����)  V��@6l�+�+�Q5Ryg"t/s:�-E$H�;zt^xR\����"�R+�8����'t�dIe�:�x).]i�t���{y���7�l	�"�[��m�z��K��|�!l�v��E'&M��y��������?a���ȇa#�����c��r��J~�]n��br��?� �����)D�*��ōYT`Ma������?.�{S��P�6�خk���f1�_rWި���x�o��3�S��e�� h��������)��L!z[����e�١e|��>�=�$9�Q�bȈ)��uC�����������Ҿ�\�cM)2V�����3ta%�<����A�����Cc���3zԧ����b��r�N�����3��-�S�H �8|kK�7�<ƙ��;���'�,^��u25�A� '��	Q�򉽿�_!�3cI��f�=�sOsl6Z��P�P���0��MG�3_P����l��Z3
{t�4&�S�2]QkE��i^w@�X�ʠ����2nZ��4�Ï��cy�2�I�*U��xXd�Zj8!$��_(��ے
�Ŀ�TjԌ��iD���/.8M�-�=�jV��������������,�c{+_��#�� ]Xa��h��������t(A��M4��N�&.�<��S"6���U�K���W;,� *�u��9�Ա<�*׫��U�[
]�x���w�~��D��{ڰIv=�u6ܥ�08d��_#�^[��6{A���P�.��7
x�5����x��$�U6S�x��T��
9��k�č��L��趼�'�ֳ ��A����+܋��������KD�g�t�R�b(6owIEm&B��ܶ�z��1�RN]1�6M�R_�0 oR�&����B�7 L�~��}��I2�5�xX�ٞ��ar�Q]4�5H�ӽ�(���*��l9��̲����5�w�8�d��$J��_b��t���n����J��;� z��2-Ln�>(2I� b�mg7�H�Z`�9�$�ؿ��L����0c�7��_��f�z��� hvg�p��ߺ]��q�6�Ҏpʎ6[\Zk���Ct�g����El([߮�sn�����+��o�ɼH�*���g'L����M�Jx���Z�U��r!�@���oj��4{�t�q̖i���oV�7Ov^n��������V�|Poc��+�6ȷ��32�Bϋ-�Sh����ST�|N͞)�h(��r:�	��W�=�����*�#&�3�o��V�8�c�B�<�j��2��)�",5�I؀��n����&��N+��u��o����Z�P�nS����D��2�?G�:\���d�ז=����?f�^͍)��Is���TQ��d�vφ$��u����@��[�pp,���c��ͅ-w�� X{N�� 3,������Iў�"?Z$Јz�!���D���a�ݸ=�!S���?�絃��L勺��DIp�hչ�>���䷕�buy���v��ޱ���	���1�u~��6���|��}���3��YN�ry�o�fb�Qբ�;3* �3B$?$I�ޫZ��L,�.�ڹ�BvfG��M�_i�!uh�q)�1��2e �^פ>&�Jn���c?6��.�ϼ��!u�Oh �a��B��J��b�<H�N���Ci8�ka����
󋠺�·�~�$t	%�	������N�6�#4�K�笧S�q� J�\�?��9��=8WX)��ٗXvt�eë~����f��_����E�!�R�� ��: S~<�dD&��
ƭ�	;�M��<���
~���]9XO�!ts�g��zxq>J�-�k�yJ�ٔ��1A:9�]���!'���`�(�����/���Ֆ�K�j�u�UZ=
�K�8ޘI&��g���n:�]�ϔZ�0}7� <M���o��;N���}x���
�>�����8k�ފj��AO�n�LDy0�� ̛dr�ӣUh_ CI;w;#{�:�ב�S�����iV�����䎰<�>����78.�}<��ui<����m�\u��W.����Ɲ	��K+��c'�F��½TN�"����b��?�c��p��'U�)TQ��^)�R7�'�)s�wѺN��\�h<4yO�ѭ�In�ҵ�P'�6;�O�x�% }5�x�3�{���^�!2�ޗۑ�k���a�{�>���U1CSZ=��8׊�:]�qβ����¤�u�|����^�[�_B!r�tNק#�$�� 0��Yz�\ї�Ų�������?�U.�lZ�V��4��d�R>���jv����5��,��p���Q!�J��':�����6G�~+*���'�;��wv��xp�)�8PYR<M�zmm��8���{��G_/���E
�ۂ���� ��f����ΈX���g�B!	������/�]����X,���������sf�>�S#�)jg)[ch�5eBo�^ ����Ψ��S�MFw�3�\��IUe#C��CTw䆵��J�ʲG(�gLW��",�;'���)�ג��n�A�`��s]��e�?�4�+iՏ�yFt��u�����2t���}'9y�
t�sз�
����[�m���<�w���;��O[�oG���+Sg�]��EM�Π- �@ �)�(m:
�sF�4�&?�)<	`Gj��>�x��f�2|b${�"h �N7�D2��㆒�Wd�7�#�c'����Y��vrO�oХ��=�0�o)w��~����%,�:���捶��B��:k��\6D��H�'�6�Bj�;r }����d aϔfo<�D1�t��Fj
˶{(}g�=�����;�H�-�F�h^���,�N�m�<+��޼�o����5��)��ԳV'�������u�k΃n�����`������)���V�c�*�3������eQ
�|yU*�;]�}���H�\<���0���X���;�%��p�hD�aQ�s�v���L���$�� �9���֡��v�(�7c��E�nSiǡ�I��I���өi�/fS:��"��A8+���h�k�u\�F3�9x<��7í�y�D��]�Z�ǀ����6ɸ��6���:f{n�)��P���`D_Z�F�)d涢��8V�Hv�i3�7/(Ȕ���^(��8=.#\��x{�Ap����<�5�`_�y��L�v�ߵe��KjeU�7C�$V�ޤ�rd����R�)JФ�'3����3v���:�s�i2�V�n�.T�+F>�=¤'�7.��:V5�1)~��8�Y��w]�j��:�ƾ��.���5ùK���ج�&ȃ��7�єƽ���fz1�1��#�M���ּ���?EaÕ���_| S^�2:���@g_��hJA4�?g�B�}���ݡ7�x��g^���(ӱ_gLc����>��\�)����/�I�=@Jw`N2+׺3�ȷ�QAZQ�]�Ăe���߅q���x:����"t���t������	Y�B�5D�%7��>!�|��B�X��_&6�˭	�l�Q��DĐ�y���א�.Q�bg�_��0 �8=�l�0`@{<��PY����o��,Bjf^�H�&�D��{�P{�� ]��)D�L�#����9I=h�^ť���`|>N�k��3.��2�cH~*�@b �����>/���k�:8�u�b���	@�&� -��p���� Ͷl��}j�9��.�U�ڵ�t�+� �Π�Jh�3��)7��H{3wRs��8X*�ܫ�2����By��>�-��}e0@��̏��5TE�҄�r��46��3�R����c�ʽRH�NK4T�漸�3�D+k{֓��%���wQ׊<���������D9�ݴ �,$΄��^�+�����Ɏ��=Lе�O�:g�m�|�@|�:
�;c��`�@y���2v��=� ��pV`����>�����JKP�=ֺ�!�<"5���~8�E�	<9^�0>\t��*`�P΋N7R�
êw��V���0[D�!GW���ܣ?=�J��t��:��
�ewۢ�m���n;�䴵�c�s��F#j��޿q�Z끲H?��#H�hD���x�(���#��'�y��������07k���x�i�Ū�o��45�5s���l����1s��g+�n:t:����|�Ɏ+��I���l7�W�=�ަ���pR����N c��k{G����:P+��݆*�N�tr�V������A�F(vN�͗d۴��x|�>�ZZ�h��[EP��(nbpl�P�|H�����|���B�k�M�r��Vx�zzT�Q��
�����;��!�ӿ����%�	\�_�,pv�2I9AҪ�e�_*ђ�`�%x`��
�%CM� ��^xH�x;T��X��$�.��0�����!!���:?�-0\ɭ�������@�� (��X�Os��m���xc�a����|d�e4��W��;j�-�T�sw)��^��Vyt��m��r-Js����S.������m�����|n��G!k���cઁn�ʧ-��8���j2l`�f3������F~1U���Eb"Q�3�7���te���r L/Ne��FN\�cSI��ϗ��s�>@ �>��8��&RY�F �Ӂa ����!��5/�9?�r���C�ÑݻR-���s��v٪(�s�����x����:��jW9M�^g���ol�HD�yzq�>eB��Y����;]��LV|�G��Ć642�~"��E�^�ڃ���9�X=>s*�%2�/���1�k�JT=yu=�V��t����ϾKj�t�2���4� ������ꐡ�L��ӝ^]��t�yXm1��T��1�I��n[Ć���!�5���,�%�T6�*J����>����4�����(�v��hTo�v�6�l]����B��T4����.q�gT�Z>�oJ/��ϙ5ys�)o$��tRv��~�+�(����)*�f�q�S��u��C�j�$�b4� 6���s�,NGҮ;������ ܬA?̯e� ˽<Q3��rBx���=�	�ܽ���N����X�3�=�#�@�P���u��]�zl�g�$@�� !Z1�>� I��qA�����Fjq���"�E�I��	E���� lW���8�z1g������=c*?���ЗE�ٕ1c���P��ϿnQ��W��O"�͡���?z�y��мs!�:ie�>T�S�1�Z�k�轡^�ljk�9[�s�igcf�c���@�� �?��o��7��7��5��q���q�lI��R�.�g��5�B�_Fv���㤑2�(���|iњ��90��@h eDv)��{H�c�N��[>�%:������y
(;���_��1F�Ո:�i�"�s״�����:�i��������y����P��A�V1k�ه\Z�l����F5����h�a����xb�i���1�R�s�ز#Y6��bw���J�Ɔɼ���{�FT��h����J'�Ƣ�f�/x����J����\��oP������r�F�6X}e�I�N��ƥ)���l�욕;�I[su�Ġf`߱U��0��F�#�?hj�(�lظ[�d�,���:�L���3���߀�v'&f3���M���N�\h��$�î�5�+�9�Y�1Q���=�w����g��+��ң����:��^�K�.�H�o���Ds,,��Xnn{��٨$���o&��xS�?���#��[������h�7I�
���N]T�,Êcf�>��yVX(wG�ʷ�0�sm/x?��}q�%����d�`�JX&��W���K̍��#/�����h`3n�0Zs,��T�;���wi��Z%Ն�`>���T��O0��5�e������ /V�w«B��5�
ݓm���,5U�4�5��6ɼ�cp�#�ѰMǺ�x���~/T3�닺��G8�9��K�H���{֠''Mn�+�L;Dˉ5�#l�8#t"�`h�a���Ҥ��K@�*��첤��%kr2����m�OQ������J
:N��!a�����Ͷ�pZ���\%�]y�E��F��{�]/��fï��v���q���~�jB�H9� ���a�r]�wi���:�H}i��N?Cg��`�+�Y�8�K��0����P(�ٕ<��gi$VH��\����D����	�s�;�o��j����&��9r��g�V�3C�&6+,�����2<<V.�J29�DiO� T�ew��L��4sQ&��mM��Y~��<���^�3����� ���g�$�j"�C�=8%J�M�����Cv�*i3k���Ji�/C[Z.�����&ĉ���6g	�2x׷��j]'*�m��$/��Ƶ#�����>��QJ)�<�n�������;���b�<��밃�q�;��atH!�^J'�U��ژEbŮc���#�O�c�쥤��eJ�G���p�#e���7Q �(zo�"���O�8��k�C��`�D&��Ҍ�5��Bc��'I�	"��J2���,$��߭�=^T��̩M.���a��C�*���	���s��ms*�	"�$i�C(&�!p��\=<�5�#���J�U��b����b��$SQ���U�����6�� �W��Y/��g�����,����̈�Z؍�]�؍=`B[��R������*BF �ҩ���{c����z�Ȗ���է�����^m�ސ?o�H<JǏI� Y�eX��>$�T�U�3�g�}�}� ��y�ܩ�A���Ru}5�~x��s���)U`����ח�Ү{q��Yo�d�V=Gi�I���De�"G�B3>�WT	Z�6
}����1�=����X)�j�Z���9���:�C;c�j��)q�O�G��S���B)]M#�E)k�Dtn�b(R��'�[��0���6���Kr�$��s�Z� �����Mc$u�Q�]95�	ś~4��)�b�Z�N��8�?1{6х���i@���Yt�.��E���US`IF҂��<�}��ǠI�Q�
t��?� �ٯ��4\ ����,����s]��i����
�7�`Z��Fj��C#͞L�m�q�=�VzQ�v���E%�4�?���L@I�PE�1#sk &o�4M�:�oQ��y�>
��s��O'u��B��պ�Ӿ� �DR��u��)t�kS?H]�/V�H�<ʵ���MN
	Ġ�b�ʆɡs0���?��8�o5W�O��WH� ��ҙ�.����7�Iۿ�D�?: ������ضq|d_���<�O'�e����[GV�����V��� u&��GG��ӫ,�8��T͒�3U���a����b2%d�(��#b'�W��ҭ����t�q��F�����R�F��E.\r��
��#��A�ۨ�^�f"����h;����aM��\���a���&��ိ#ez,Z�cy#�{5�&*D�|���_6@������/�<[���Ec`� �ځB%r��JA��������BA��䎀$���Aj,�U��[E��㦽8IX�ek]3T�t\��<��dZ�� �G)l�?�!�Df�^��NZ����X3e����Ь�a��4�ϼ�pS�T0���]����H�o�/�U�*�����ĝ� ^n޿W}����[��,q�O�v�����I�O��Tv�����f��	(ӫ��*c�>�k״�����/8��u����Xd�h�(�;G�(��ˬo���pf�2
�ܒ�2�|�)!8�^�3وW����}r�D��i=�jR�b�.��B��L�0�
��.6�Z�� �]톐:�po��5��5p�I�v^��6��New�Q��$A�W���ؗ�E�V���8�y�pq{��T��,Q �>���ށ��-`��]a��؟�^��o�I���|$�� �f�J�/k�Q�g~���'�$��~�,FF�,;�W��K 8?m� jr�Ϳ�lҺ��ee�4֏��.y��[�Dp>��U�VHZ���`S;�����>��X]�}��Ī,h����Dd0m3�ڧ���8O��VjI�N��y��5&�d�b%�y>�	t^\��<��j33t��\\�o���h��ptQ�v����g'cI�+�Gk�6c1D$��g�E�G�)�*��!�v����ˋĝY:���Nnݎ�׎�� S,���8���:�_vH�WA�w�`�$ǧu����nw����Z�L�O�}��bmm6ڔ;Ҙ�q��8������� �v};e�%k��d���nց�t�p���X�����~��5�	� �ކ�|�)��#w��1f
V�I��m"y"W�ucm��7�f���a�h&~%0��<87l��>\Xvq�#>;�I.�e+��W�@��yV؜FL�}��<�mgj�I*!�x$��qm�:f��[԰�ܞ�*%�$���u��?�^l��s=���r��}�-ye�وY���~�� 0��"�Χ�_�8�RTe&F9�qA��ݧo!����؁^�ҕ��F�@�b�ٔ�2cI����;��*����۵�\���i�����^j�hq;B�"�f���N��e�pص�q`�Υc��FJR΂b{?��o�j�F�̓�%�Y���7�oKɣ#vi���#%� �\^�Y;�a��+&��0�����8+g�8t�d��ۉ�pҦ)�M3��6�G��2��5�G�4oD����c��U��z,'��^���
�NԲ�l�Qx�X�A��L�i��8X
X����T��W2�����>���߄xu����R��#0}ȸ��þ���</a7}YھӐ�v�F�[��;9�-ݎc2j�y{�.�/����_��ͶTHɹ�APF���$��D �FB�}|����S>^�u���u��յvIsh%�u3��GY�B�C࿰̌�Ș�yH���M`�7���뽖�i_&3��6xa�����kSD����N���� y��S�Y��/ʻ���
� ~�56V�wܴ��"zэ�8C��5!&ZS��æm�Ȭ�����ތ(BZ�,WKao�6�ߌO�i��*����u��I��`S3M��Q���K��E��B��>��\���G��r�*͍3kf�\[:W?�� x������vҸ[|����Gi�*�-+���Od�ىiAezax�)}5��� B^�[֞`�	>�W眕i�SQ��@�ĺx��~%~�چ�����H��(���b�7����w�U�|��ї(1n��zU7�I(�:^�[��@��Z�C�ƝT�ҳ>�E��@ +H�C_�#���i�1u�ִ��~m`����ƒ;�K<ש�ucՃ����^_7�<a��E�(˺����v��Q�-՝��[[S�Q�J�����ԅR�MFier�&����qͱ���.k�+����p���q.�|�$�"�*�d1$$��J��߬_�j�QF[���yx�O��wL�a�<�\PV&p��d4�;u�V�#��kP�i��7��Kb�a��X�\4�y�!`��S)�w�P���x�޸i�!N(@����$�9��)8l�y�,ǵ�6�WG��}vۈ�Ţ֦Vl�<P5}֭ttڻ��E�5^�l���fb�$z�!�'��b�^#q���r���L��%�M���Na���P���-�����S���t��w{|�ࣧ���D�a�!���I�G��~�,�ˋR �ϑ���f��H�L����E]ܓ�k#��	,Kev�s�h�g�;�3~�p~��ԋ(���o�fr`���I�T������:�ZM\ѴHI��Q �3���.�=�tFp+�b�`죧'19$ū�Cg�Sz���1��Ll�>�8�c)@�\d]~�5�oCO��v7�@q �v��ngM���U����~�=Z��m�^��������43�n�w�Ai���$P8��B?Kq4��A=�Ҵ���6'�����b��M��X�oh��5��{����ײ�CZ:c�ƪ�f�}�¼�@���~]K��z������%�3K����<	Y�ҬGlٸ������`Ng,@�M|�g�ޛ�w���>����!Hʭ�&�p�N�H^g,�p;���旝���eR��Y2���j�qi���NW����U�u�$��Z?W�-��3K�<�f+a00���Vbh�ޏ���-�k����!r��=��,B)��]���b˗p�0���M`���}^r!S_8�p��{J7X�לٹ�QT����������QG��|�l?�bRt�����z8���q��7��\(9��������f.o�	�9?�}Nn�v>"Up�2Ϧ���H����U�(��.�6�oZ�6�k�^�Ȩx�طqN@��
f]�"�2 F����#{>��Ʉa,7w߶��4��Rt�vЪ��RT�Sҿ��Aԛ��o��NS��$�8< pպ�������{�s�O�P���t�>*��(�[C�6^�-A�J{��eId<�~��a��Wc��D�/����Cf���)�9�l��0�l�.rSP TD�^+�/���3u ����t0�vF�Ȇ�Bj)#�v�[�érX2���v��{P�D�
��Ƅ��(:�햣<�$�M�3� ·�u�ϖ��_�r��"�	� _XG���!�6/���v�UU?[.��!@Q�m�
H-�)��a���}]8��]m����V:�|i��+&?�I��.����_�#����Ꞃ'�"f��}30k��`J�p���U��N�%��6}��3J	���g��4��<f4~��s#6�mى��6�ާ��P���]�=����
��[�����0�h�ެ���Ѫ
]H�м�$�XF��_ЄC�)5���(��{����[���?g��x��+�O 6DGC��M����#ݸ��C�$��Za�K�{���T�،y�g�(}���5�9D���C�����N�-o�pޗ[�.2�㬞aQl\Y���ɵc
@��*�^/��GÜn�9@sk�{�ߣGsk}$�!9f�*���9v�aeo��|Ӌ"�Ӎ��,ԕ��[��4LN��5>#  ���������/e��>1�콰
;���O��!�27�M�C��њt	|v 