��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&��n?��1ů��> K�-� Dy����m�����|䰑fԵ�($�ݑ��u]Y�X ��x�%(A�Q ~6�f�Ь+��f*Ĭ2(3g�p�Z�s��ƒ��ho�u�6C��5��ʘuQD#� �]��:T+��n�M:`�5�2��ۺʣ+�֊�����<c�u�s6�S�$J�ꁕ�ڰ�'e�z��G(���E��m!J�Z���A�5�m��%��
����j�i��6C�DE�ɬ���=��ܸపr��%5o`.��SPLX���ݷ�]�F�2�nLj���ld�|2�im%lj��x<	�2� ���}B+q$�L��[i�ԩ6���(+������?μ ����}�����J�\�5͂P���å��\)GI��wٮ�)�W��G}���0� GA�{�K�}�C�$�f���7�8�+g��2I:CY����;��ԩ�}ND�#��������L���s�>W���iY�4�L�;+���~"�ܳ�q��D�R��/n[�9�N�4��9���E]��]��|����UJ`K�5,Kzi4�3�D��#�7��<p�Fx̯�����:��g�G��5�)�*͙7H4�Q��rVa<r<�G��&��G�6u÷i�O��(��*�quH���	t�a ��}�OC|�1��'�d9}a0V_�U��"�1�X���Ö����ϵE���Դ��5\VЊR�[)�B��}bww93�w1��ҝ�l<qd
{����mE/��g4���ѻ�/{)���{�f%��f����\V�]_�Y��C�M��+ 4��x�V�l���H�C�(/U�d$57e58m;1��F^7�3;���7�.p�M���X�Q�k*��qz��~Ys.#_⎭n�R�̞�X���ޛ#�/�ERFڀ� 1g%$�O��%��gy*��=��9%,��_��	Q2�5��A���X�f,�S[7@r}v�U8� �Y�eÈB�CG:o�%��ӊ ��P�ǯn�`�=Hу
���g��\��R	@`/T���n��?�O��~@�!����u� ���9����%q����Q9���(R�r9���r�_�t��N��buY9���,�u����?N�\!t�~�#j Bce<߬^'�����MКSD����h�����![�e'�!WEl�Ǻ�_W��� ��`�%.�u������Y9�W9ƶ9�Y�&�����6#�r������;Ƈٟ��������b���0�3������T/�Ҵc
|����y>�� ��A�����M�X�	򇩬)���Z�h�5������m�'*�d!10Wv��CȻ���]��GW�.����0GZ�$���=�n"5if��5B*�������c'2�O6�*>m��*�E�8)��޲�Sˍ(�QOZ�!7�C�(�`�Z%��%�R��綺VM�qؿ�v��`ɛQk;�g\��w!@���e:�2�����<�J���P���Y�l6��/c���T���+�V�!T������չ���f�M���k,��Q9��
�~����>p�Cs���^���� z2k����&�m�u��ox���,��L�����Teغy�$�9�O�M�������(����pͦ�Ĕ�3�x�@���D˹յ;y���=��r�7����83�]qB9&� �b��\B��ŗ�q�5Ķ�|1���� h�Օ���zCX�܁I P���q�l���K�9���h4���+�w�U�K�Rm��7K�ՐS��x4f����m�E�!��RE67N״O&	g$}�@�A�"�%����.~1���u[?��q3�$R�g��p��E,��ǱX>_u��R���3�ȼ�1+�{-*%J�>a�8���29���!WM��N��7��d�O����aO�-~���_s�U��_�Ff'�z!2�Z}��{`3�Aڠat��ه���{[�����@V'���!`�Mn���J2��o?����fjy�I>==σr��p�T}ԘT@)yIY�n*A�<DH�P�!\/7Rݗq������2~X7|2��	�SdnkԌ�0��m��ŷb<Ӽ-�q�0L{5[���ӛs�Ufj� $���m����)|��p;D
����
��}�71�X~ �@��,��d{��}�]{��1��&�/�}�-�?����[��!`�k*�Һ7g[A)ܩ
*�]�d�d�ߺ8��Ҙ�aXF'q�أ	,�!��26A�Z���C�rA9 �sIo�&qr7��Do]>�:��r�+On����YKǶ!>�:�구�!�-����/�`9`�����vɩ8��u�����>���e��<�֯��	I�D3�ja�f�Ҍ����\��t���C�T~qn��"$J�5���kD�����. F��L��Z(����I�~���?W���qu�����D�ԝ���M�� .O��Ӝ�g�y��M@��Fs�����4���=Yժg��)���KV�j��充o�D�<u�%i�pQN�[m9��s���:`Q��>��i�z��9ƃ�6��>��{y��{�F8�Ko �J&0A(�(��f�x�������.	붔+��AR���ZY�ƛ��#�N��-|�)�b�U6�T�|/�9�mYuM�Ϗ� 1�t��Q��沭B0h�OC�(�&n-����]�=��R�ꒄ���!L�`Ǚe���u  0������Z3$)W��!R����p+��{C��'�L�=B��P��jNn�$7��CHW�br���C+d�2���?���*�zo	
��˲�����4�B֘���"���.t��Hp�A:��n�+��bi]��I�������j��,��t�R*Ӽ.�_�R�
��<��2�o:x����3�6{n� .�!�O@��J����M��N�ꀕ���L�(?���'�N"��Ϣ����M��JO�{�u��E�(��FW�m��.�����T�*�|�C�������||ͤ{!]%P�b.؛��,͵�&�y�|^��(���(���L"mܖ�T;�yEWt_�������Фq� �R����ۏ_��G�w�auj*2ۋ�U:x�T�a�@�P��A����%�tH����\5�kP:�	n�5��h�ǣ�X����/���'��=�fsM��H*Z����&;�޹c�����R��.�ó�֮*�q��t>�&b�;tXz%�KR,�i�s��hX�8�ļ����&J�2sG4�r������A���c��Y��P��KR������<5����^���Q��>>�3j���0�I��l����ڽ!�T{��s�E�������IQKĀ�]/X�����{yCc7t5�
p,~͵�S�8�
��l߭���U����_��8�s��<����:X���;�M�=p��M[7I��3X�i�s�\2����Ӹ�0*pe���.��V�y&�+�c�)R�316��@�ъB�6��@�41"%;�]r�ݒ:� >B���2���hr?�0ߑE蛆P%�?	��9���� ��_@ŗ��8|��z\$�ωL�x�m�ϡeǐ+��b��L��_�����\r�4�A�w�N_�5:����[j��,Y�O���:=W������'�d!�2:$<��Rn,�,I�.�{�;��p,�Q�U�0ލ���y��Rr�o����8j��W�
�3�:��*:��h���hƙ
�ڨnP乼���Gv��r����a�!��ri�@�x�.��#�>���GT����+�=�S�݉t� Jٝ�S[��ڜ|X��H�::��`1��V�z���M���e5X0��rsB�?��%��d���A���OEx���/ �M�U�<e
�i(����8c��O/TH��	A�����6d��k�Yͮg����8G����dD��̈́���,��9�F۹�]��;�b�Q?�5wޭNA����#i?��{+�b�)�WL��J=EH����|���>q!�=�#`�,��q�,���?�=`�\;s����.������GȠ&E5,"a�Y_+=���E��{(7�mg��!3�+�����V|]��ـ����
�U���˗�fԒ��0���u��k�dn;�ɨ)�=���a-�M��P7���-IZ�y���Sbd�,�PVEW�փ���&����0�L��c�����Y�Y	|J��G�i×�c��1��fO?������03ESBq+����p2���H;M�4�5�<��[�S�y�6��,��>� =g��اB뙘�â=��,<��?$��f� ;�)�R&��%���;����z�6�q���MG�a�g�?���gS�	�Z����U9J�Ϸ]��P����Լ*�_ �B�'�_˼��f �,�m��Jc�M��V�%���Yĵ�X4@bKz$�,���j�����G��ӧF��]{�	(^����Q����|���
ɑSu{	N��)�zBW����r�R�I׾�����P.c��\�T��mư���I�R��oA$��ݷ�v�����q���e� ��:�˔d�O%��@��]̣��&�k��o`9��՜�����sp
ĥX��u��ͽK�[-	ߘ�b��z�gުtΖ��y$�MM�B�)Ɏg���~5V�$�q�Q�QX�D:�^���a����`T����wA^(y�&��́ld٧Y�Khw0qg7�*(�)B��[@t�k6��,f[;��N��E���"ǈ�8M�����+����bl�^	ц<DnHĆ�;���B�����tA�A�<�="N���2��H-�k�r�_�;��)ܟ���|�^j/�+����]6�l.��!���wx��3�g��zQ/��Ϋϡ��
�z�T�F�(^����;��v��˟V��)4���񿁄�'�ũP��AN�ÏW�b�F�"��8;]��.�#����ĥ�J��,N&�V�ʾ���]������U5�n��.�o3\��ۗȽ��,x��n�Y�Z�∄b��>��|�pALI"s!,�J+��6mmēe�kݬi�E���PD������Pя/��SSCM�ew����|��z,�,�	.�7�!��h���*��"���	��WlD�	�뙫y�طP���U��iX�T0��M��=k�N6���/���rc��O����[ܭ�?���7Ĝ�����10(0�/�F��Ӄe�ɖM��~0'�s��!�g�x�p�����S�2Tș�;�)	��~oM�0>y{X#˵L��kę->�3�U&��R�U`���rN�� �A�����T� lYV!���=q�D��ib�u0��Zz�>�C"�K�Y�{~5�G���Q|kN!�ɏ�3o�x�
K���'%��-����8��������6��9ܟ��T��M��1/�K�� Z�A�sxS��8eݪ��t5���$���%0����H.b��M�u�	$?�:�%�<_�R�Ӫu���^^#�é�S��T�P./&�"�{8���gN���u���;���\1g=���?��ftAz�wtB/����럙<Y���,]����mF�c�K�0�F|�jY/��N��G����U��0��C�T���л2#��\O$�rfQ�#"���Ve&�������~]"���>N�Ή=g��x�$�Go]��^�ܘ��ǶԆ�J�Dƴj�v+72�$�j�� p�f�Z���σ�]c�4{߸�G�*@�V�ks3�{�:E8V��&�ħq��L���!Q扈�jx�#Y{�z3#h�=Z��6�>��f��7�ӑ�	N��t�N��)���fK./b!�iȐ�nO�����а۪6�3�["W������.��a� $�]��oL��l�B��s��m�����d���E���@^j{V	ޭ�����bz˿F#�$>�!ԀY��јw<��z ����F�ڽ(��]p���^r����~�Jsr9P}{A0��Λ��X��B'�ȴ}rq��z��_X��G�5�����d�:��W�L�i�w������y�_��BE.X�AӦ$�,Pt�����G?��*3(ƅ�-5p|��׳:E�@��_�"� V
� C�f�"M�"g-���R�/���m@{
�oa�=��o��,u�a+����$A�,�o'���P���H��J��ɭ ��q��_V7!�3+u�pOk��	�M�˛���=���'����~|�KZ�����;(���ګ��` �e�����D��8��2%��f1������s	Td�J�^*o���_�4O���#�E5z��c���۩W	&�Vj՗�U=�!
6lMJ�Op۟�!�;��O�5�)Ĳ���ih����z{n����o���>��}�jm��f\����d �2ys�9��v/F7�]�u���T޾��~�]��(��JZI��b�?Q�	}�+�%�~�[���n��W������:ď�t����{��-g�~�?Νk:5����#P�U�VjSw�Y�O˿C2&�t_rЇh9�MI^�ψf�Q�'������}�v�Y*%+ ��*�KY��&�>V�^]?�XASt�>Ϙi�Ӡ<J�g�g�1����9����(	��m��=B��J�A�����Tn!�-{Z��O��g�a2�*<q?�.gD}G���9[�&TE5(Kq�P�H���@X�
���~-_��@��A� ���7^�y]v�h8s�d�鍧�����<��r�]�{�a��w�A���	1��l�3�|�*���.�˫j��&1eQg�Kш?2	Rʓ�ki.vFeM'c<�V�z�^�� 0-��m#�E��f�X�9�^ �Fm�M�]J�+���i�xmߤ�T����+�wp�T���)CJ�D�
���y��2}�`1�y����vW�A��2�z3quK���ㅇq"u���!�����C:����j����^{�cJ�m���N��/n��9��^�Q�m�?�)`<z��3���m�T�찪:�+�R���ڟN�I}�!���hZ]��.H��fH�A(��*O��,*�WG&��M��-<��VX>
��%��ƅ����PY����MlW�m��Z��5�<OC��JwD�c��]5�o\t	Lj[CG)�xۅ����.
l7���H��_�
��/̜LgB*��EW������!A{���C�D!�ۡI,rt���.2�쎟ń��4�
XkX�dQ��ZI��NA	��t~���yR�-_tD�ۂYےV����-�ߣ��s3��@ѡ��9����x� n	Ȍ0�i�o���½�u�
|�|M�	�"�$?�Nx��B��q���S�ܣF19n�HـT����9Z��`�m�uJ�:�HCmR�������6b��㘌H����5�Ɲ�+�#On��?�&�5WeP��SWAy^N���cnJ�Q��%� #���O�I�}�6T��O��"Y�6�&j�%����S&D�n��_sVR�{Q�����Q�5%�=���!�k��PO�@�6���ވ����<���ƅ�ֱ�!��b�(x�Il�
�[�����PA����(^U����S�{ϸF�l��祳=�����]7�w� �2�т�ztD�hp�,�=.j�mm�@�rjA���k˾ �����9��C'��@ޖn��C��Ϊ>&�&fn�*�5?Q~�i��9�@��7>�v?Bb��w������@:���?贴ʍ?"e�EՇ�fUE�QxW��vVA�_�
h��C!��=��'!Y��mz��=Y����i]�������l�[��TLѿ-����#09�d�݉��o�[yAB�9P-�yϑ�#��"��l,^!����!C?���}:��d�I�؟g*���t����W7<p��gK{R��#f�'j�T�����,��\�$� ~X����Q��,ӂ�#�����z�0���`e��~���r� �*W�'�0�+����d�("��Eڑx������F{M�3��"����S�T�7�����g��/ISj|��|�%�Λ`W��o-?��=u�YP9 �ע�L0[j��i�ۀ��9�*_.j`ǵP�Oڢ���o�9I7��w���ܕp�������?pٔ�������ga�[��_�/�8k��X�P�*"�լ�������c��qoC���;������8�1�"n;� ��b8����˜Gtl���4�b$�s��՚⎛a6*���|Sw�Ƥ���;�z��&@��B ��0j ���W5`��<�� �P������N��i����8�u�S\�Q`�������$�	D��uª���gM�0"�^`VV'��@�8���"(5�nׅa����0�}в��8jt��s����:�fIӬu�ǹ�{m�Ct������.�!��q���_�_D.V�"���9���A~�;L��;��򉱢q`VU��3�k���S G>���2.X�I�*�.s�B�,��� {<�,"E1��5S!L���[I(G�k*AOϱ�����L�t�k�j�g�5���伈io�T[�+R:��O�iT�N�H�(��S\^�~���[�O����f羨4�LL��rn��rg}��� ��w�J+�]���ķ��(��X7[�P���w�8�� �t][��*�1���]&e�~��ފ�Z�a�
(	?p*)���N1�܂|��v����À�U��	��+��5�K�}�$���Ñ铼IN�U��8@�S��M�[M�ܿ�*P`�Ď�;T\6�%��?��ƮB����IAc��(��^2uy�����g��
�''��Sg�sqY�ye�>v��:��1� ��5 )���(d0��'����a��Y	'i�`�nIڢűa��jP���F����p�^7�A��q_�7#+�L�Z�nR*�{wH��X��G�2p^JXWO7�9zU>�g���2��k3�F�c�!ߨ:h�kr|[n��1ZĉS��4\m�����)��d���9jiL�O���6���*ɮ��H��T�@>��,*�jl_��:���i�l��}_�?�j���o�����7����N����.4@�rqN����t����Q&��~ԣ�*8�d\H���6�O��L�. >���8\����||?�Yw���GT�-=�о�L�6�`��n�i/b�t&
�'dK�����]K)7&���l�_�����2���:��(p=������(�	?1��%�Y߶i�޹�+�Ⱥ�uo{^nF��"1>�2�!��Iˮ�8��=�YJ�x�r{E�:iZ<��I��Dx\4Ko�tK ��)�:�����-�7��ͷ��?Sa��t��:L��f1����y�f�4����q6ڤcg�������#���}=��I�r_���r��
%(�A�<�h	����x���J'U����?*5�c\��
�m�%0X�1�Mt�u\�������4�"_m��j�R�d7L�;�S�f{"7���� 4�ør/�5WE��l�m�<5�*�ן1 /n�bL���c���6��Za�Pz��X '+غ��M�|ΥK}�@:��iR�~Ȋ9�4��X�]���tqA������N�w��6hLݗ��	FW��0x�r���e�'f�-� �-@���/���~5XӸ3��Q���f-^�D3�]�Uhr?���.�i��.g�v2��]�ƭ`�־/x��i��֪�w0����H��9f���^��6�l������}_�wX8��8�kH3� �l�˸Kx�ZDz��U���Q)���o��u����q��oW��p�1�����nK����%�,n3���fX�Xx.���S ��nFd�������7��3 z�M������:ٖm��[f
��,�Rtdkd��D� �/�n���X��%��Q�v�3��}�����k����m����Vi��	Hj�L��>/��h�ܢGÄ����H�H0E��T�=�������$���E�Q�-ָd���!����C �;n��\4���x�y|QW�"9�+��^�O��|]�X�����|�$�XW@@XM3��%v���W��]�y�`�m���K\<�g=�%@#��i��A��7g���tlגE2C��̩��PLqT0�T^R�_pq44���z��l�SÉA�B������A�aF������o�v�tx7�ZJ�]
�I4�l���%����� =ͯk)����H��4�� ��S���b��5,�n�����Bf7� ~�U��r�N���U�,�J6ue*y�������@�����f���rA�R��"���*��s�\j�)�4��5�ײ��آ�>7������x��p��[�א�R�LQ�n���%K�'%%���$Nw�>�?[$ֲ�C7���k��G��i	M�>�����G���+����WkX��T�?%���	�����ޟ��]G���Lf3�)j�ә��B=��⨠��� �a����>��1��m0H��cؑ�a�Q�R�(wT��lE�4hR
?����ΓQ�"N��� �ް�@�W�{�2� Lri�)-g���8��:8� ����+)��T���BУ]�X����3oN�cwm��s�z�1�)�z��T%��B� ������5NL��1՘�q���� � �y�
��=q�j�|�}����S3�i����;���K��Z��!�u�����jiŹ��ug��)$���j���n:�(w�� /�|f�_tR[�~�"և��Y]]����HV'�T�vժ�/�G���|��G
ZU���{s�j^����m�C�9;��������-����Ux����2�:�����B딸��>T�,����<R﹡/��@r�jQV�eGt��F�>< f`o�[������}�G���3N�8����R�	�yu��i��߼�Y�y(Z�9���܊���V�ϐG��!�음³Y#��[.eUEי�0�*a�8/�0Q@׃�e�J�*+>m����i�>f<��Gg^-�#��SڄD"fwݧ���_o$DPس���@�m)h�h<�LI|��5��<`�G���p=�D��7�!�^w�Q�je�Pó�3dZ��#�Q�ϛ����u���2�b�WP�?"4|�5]�?������	G~�z�@\c�>�:=�o��U���5�|����֨%���=��T��q_hxn�����ثL�L�`��IH�m#�2{���3�PZ�d�A��U�u88PЏ��1��2u���}ɍ!��az1����Y�L���ٻ4L�G�s����q	(m��\E��M	��b]�RQ���zs�	����Em�̕T�)=5���'�D$�2��;?Ě�p��G�i�=�T�Q���l�#@�W��i�2Ոq�$ht�|�sT9�"X�2�#X�k�/J���.Z�UL�b�&RI�(!����8����/�ّگ 꼮W Nl(�Թ`�(	]�O�L!�HY��]}��֍1�4�����[�T]+a6�L�Z"�_!{Z���@��!�Ua!V�^��@�����U6�a���jc5F�UͅB�`��mx����ND��9�(��;�*4���n>��+��xu@	,t���m�3����ƥ�2G�JZ�S�O�ɏ�m�V.���?ƈ
}�ჰʐ.>o5Ъ���?F�U���CkG��#��@&5�@����>�Ozte��X�`T�z9j�q��\K[lcT)��CR0�X��I���m���tJ�~G<\j���֨��T���6ĀPڵdX��a.~D�0� ���g�rB��I�_�F�Fkc��zǯ)�Zh���bW�n�~@��VW0m	}WDn�R����
>_�__{:/[���M`��&����ѯ���?�4��ͺ�݈U��a��M`yJ#^��p�==�{M�Т�P����6)0V��l��g�ݦ�EJ����zC�q�A��Ч؀y��?�˭X��q�b����ƈ��@A�|�	��У#�����Rs��\,4XX&	�'�֓$r�F��zx�c41��ktU�l
�P �~��N����4���+=��!�9	���5b`�G���w���J�x�yā�7_H����a���u[�M���9`m!�TV�����lg�ygO�J��Ig5�X���~��.rǭ�Y6��=�>���V�1�v`9��{;ܤ���,
V�;i��<)�͈���X$z�e$���E1i���'�<��}ML����jҢx��(�P�bT��n*	����
]��#��efqXzHu5W8ѱ���8z�v�9�H��8�a��'Y��8F�L�$H]�	@T���Q�,��j3-�r�?�|~p�hUy暘S��x�^�Z�~c�\�!Woc�J'����5��!mrzoP���G�8n[�u��ig�9��y�D�E�S�"S�/"�X#nLO�I��lc��^���}������"���b��-k�s��P�{��{xŨ7�e�uzۍ�D$]v�U����{lS�����$kߟ�c��tex���2Me cl���� ��{�w�4�$`Z�t~MT�Ss�Ҕ�\7 ���Dq# �����[�uvۯ�B^�-�����gί4�şN�G��)�b8'�����8����� 0],QmSr��+���A�X%��i���o5�����9����a�eyv���΂��B�����v�=�#m7G�J9T�}�c�:�O�hX��IG�{b($U*e��M�Ӧۛ�wS&�p�T2���!X�AҵlK�/��4�ۊ['YA�������*f~���n�G4 ���7�T�1�-B8�S.��
\9EZ��'��N])b�s\�4m|G��;��S,�6��r��㌑���<�q�>�x��S�����V�<W� {n'5P�6ؘ�𹮹.ٚɫ���D�mϱ��{a������a���E>'���L!��v:����^���f�>8��`�'���tj˓���[�K�<�n?�&"r�b���^�p�$֝�3�L�����7:�L����/`��+H�6�'@r>ƅ�]I�#w
�7ZQ���L�(('�jkIk*��Ҳ���wՌ���R�_כ`�����X
ƕ_������)Q�_r�U�@�Cv�qɻ��(��bLG��--�!u�6c�L��Ɗ:g` ��6���!����e���3��yl
�n4��_5h�g���
������[o����mk�R��I����|vS�Ɠ�<F����
���:XYr�}G��'{�vHW��1���lC��j���
�WH�ӇF�߲���<����5�iƐ��';�Z��d9�t�����uC��D���|��ST��x�дH�p�V�D7�����'!�薶?+���n$�
�R4�D�����}����T�$0����&�M<�������p�:8S�������n�D�jAA�Q��O<q��b��k��I�pa)1I�]�-�}��m�=�=P�NK�.�63��Zc�f�>&0��~�w����\?+���&�**�8j��]W{.��H�̍����n>U�E�Wd} �4Y�@|#�|����)���hW&I�R��s}E-�.��p�1��N�����A
����«�.�M6����mڥ�����scl�`*���m��m�G����#�Q��0�H�=o��bԮȔ��P*�7��i��6�C9���w%���Pm
Ac�Ui^]�9��\,���9yO=����.� �m�� &1�bJ˙�"��(KSZ�x?8?��Ft���^����ᇯ^�i]���nf
�Ӟ@Rb�>��"_<B��0��a>�0�9�qו��&7֡HlrlH����,���d֔�
����:~�5m�Ջ�|I�q L	���P����,z�:�ԡ� t��S
���3�s��t1����%*��m"8��Br|�������_�.V���"��<q���gF�^N�������32gU�Q�:'
��6�q���r��hr��j���Ґ�g\�!a�t�)�������	[��P�S�T�@D���nz��L:$��r?2SwJ��K�����3w�TϠ��b3�śx�j`�<Mz,��!��,�ZDI"��;U�(& "I�g}CI�-"�;0)��#W��I*�[��)�ʛ��D����I��a������'��?������tN*7ߘ7a����."��%�چ�*8�s��/\,2�x�������V�eG�@�aq��t��~��i��v͉�k��V���t�E!14�~�9�5���E.��ߨs�;C����A�x����"����+ӗ�s����a>�$M�C����U!�3s��N&��ѩ�-,��rH,!�"D+$;�F��`]�,Y$�5V+�dt�m�n�,�I'���5�}�z�����	�}Z���� �^>�@�����{3&0&4�����cM���FӺ�ֆ��ty�O��z���(�'d~��2|x�2�)�Jpx*,�5��{�L��aW�k��k��4!�`	��ID�邝��:%�PaC��fF�tĚ��p�k����]�hV���0��s�T������`�arW�i���I���v���/�`dP��3/՗]m��I�HIE����dv�5׻���pkܒ�e
�o�q4��-vݝҭ�Kplˏ&���~�f�Ub�F�I O��\xg�qԬ�;c;�u1�(��.%&�u(��ܦ��!+rS��_��A/�T�R�hb��j���=J���� ��+;�jT��.�1���YaT�\Y�Ǻ����ن�^�G�\���P�j#� �0��]�)' �Kn\��M�F���
�v�h�rƯeY�O�:���bJ���]-�q���p��8�R�hg����v��hC�`p��<���	�?��x�Z̸���.�&�1���f�ɹi�F�bk�/mU֛���e'�cE/_I"I���
ޡ�������z���>�KP�9��6:5�����|�`�;�v��yn"��pWe_�*T��5d�J��;n�m2	�-Zƶ�Ǐ��ݓwbL4�<���\*S�I����^?nJ����K�d���5L�Ǔi$�ˠĉc�@ �zܣ�u�X�ިv\����5���b;����1M��kőd��4�iH"��H��á,j�8�h���Ϲ�m�*�i��^��4�S�SJ����� 
��:��M�u����-��h4"��5,���1&�G�3�~m��_do*���"j�������/x)�A�p�+;��r"����v�	:m���	TC!zR�w�b4�}���V[_�3݁�'�sתLkK"��;�f�V�|:��=��)�L��8H��dvٞ<MNiuׇ��,���.P���2�!X� �n�ޜ. �]>��j~��zM(F i�A ��x��W�/'��r���l
4�X-�ЉX�4|�5z,���I�Ĝ�/΃�NH{)�J��]�a5�r�-X�8r�Ԏ��ËQ���>9!�#霣�R\U�EaD�8T7M��	r�ʽ�P��_�M���Ɣ��\��iz��(��9�IJ���f�$N��=����7�F���#��S��|ސ?3�T��P9F��,�U�TF�^q_�� �^a���?��^=��X&[��x^�'�� )���>�����޵��a�ðˀ'<*�Z��K��l���l�m��8\�FEH��#X� Z'��1��(��=����E�5�W|����ȷ�ιsi����R>��ư�o��M�� 4'�:o����~Rⴵ�6�'��Һ�"����FC���i��'l��Z߭��+���2^Ҽ�)e�6�x����7�2����X�E %a��ܰ!�m���Ţ���{�����p핗Y�Ot\{��z#A�Z�u���_�|��]�t��C���tZ�ܾ�W�\�>|�rت �)
�!{�{1z��*No���]�#��__g�Q_T�C�c�-q�W�@$rfWX?�s@��I@�H�҈�@j�_��F�yR�ǯ��0�?AB#+d^+/'ʩ���ߞN��+�ûmέ�jj9���1F5O�1�^�\�E#�d��v�Ȯ��z��,-���}�"�r��>_ҿ����`�]B�׃�Uzғ!�;<:��2H�	e���*u�Nݝ�	#�
93%�w�����?h����
��_ۄHg4T��	fF�j�b�\y��O�O�#&XN�k�Te��62�8�]��Qu�>�^G.f�� ��m%��W���OE
��N�6zʔ��u���\�v���7}}�p�G����I�2���Q��>�0u ��0YqT4��b�{�x�QB�}���4Z̎�B��݉&�e�l97bdL���뤂p{@A}f��U�|7��_��@�=���a�*�㄀pU-3���C�v,�|U�=�o�����GL0La���bP����KA�ܞ��̃n�Hu�H�}d\sh��I��i�(�H�����b�ɓ�	��uׄc��o��#��hd�s��|�/�_K���^']�x��B��E�(�d���d����m�U��
ݏ������m�\G�(-�lT��qM�u�� ��	�HG�]�Qyz}Ľ`���I��Sx�ӄ,)�Fk�݆̫��V��Y$ۘ�CYl�"~���N��[lX��b�vQ"�|���r�Ir����WE�ղ��C�e$Ť��YM�e��],���<�����2� �\醄t�$�0=�O��^˗H��/���mRu���T�r���v?_LDL�i%B���F=PN$�T�Wo��\����� �5�"���;�`��ur����G����Ul�f�����v4n����/]�1꾦����.�������4q��O��®��;���g(��� $vp�~
�`�L�|�\�Z�FX��6�kYk4DA>J �Ҳ�h|��Y/�Fgǳj:����'�Ig��4e2�e2�eA�C�{n����У0���|c��8���2��س�NzJX��sJ�Fi�N"T͵��}L5$E����r:+ሯ��L��?h!�שm;(�;eC�1�*��#H���ւZ�K�������׾�����ͣl�n�Z�LCG���=u��H��n�������s��,�J�JɎ~����p��BU���I�/R)Rd@Lm1a��)��(�u�W�$�b=����-�󪽦s�r���ɐ0zY=+ r��;v���%d��� w�Iy<闗\a:M���2
,�h<��u�|Ia�����~��rl 1�'��v7�j͓�<v�,_-xġ_���ݺ��QdO����Oo�����&�����>�9*����ç#Cy��Ej�3b�sU�͑�= u�2疩ۃ.dW����#���<v�ʯ�v���ey�d�l�ZjN���^���;r��rfy���wrոwϭ'�7��2-^��0�NJd�zFizd����� *V>�S?�����9������pS�Oo� �m�J3Y�G��^ȳvײ4�[(D_�p͹E�W#J.��!�b��8y(Њ��n�D �~O�2$X�0S>�$C�Z�3=5m}I����Q˞���%��E�6��iy��튦F��z"v�@�q�5�0�:��\�4$��DTɓnz�[��Ǵ�3K��Q0����iG@�T�9m]_�4r�]ލ��%�Q��G�EA����)R�i��Ѯ�k=�W]&
�X�Ob%��P�!n��h�Je�&�G�u�������x��)�d� #��$^����������R�r/
J��g���.�`�GB͡'�m�|��m_�J����M�����Fc�P�����=�� ����Ba���aӚQ�PЏM���A�3�33�ۗ�iW:}��n���ŅY�Q�7!��:Po�����U���~�wB���eY����;��L��<(u8�a�p�f�3[_Y*��) �˽<�����N�0�*g��*YSz�Cx�� ������L����.�J +7�1���AklYp�Rt�j)`n���v�����U|��� �_9_m"	"�@�C��YݸW��*�����ē��0ొ�C�̚��<)�,ԝ��,�n��~�&�R%,���|HlN�W��zI�P��-���c�A�������7~�D܊R������Ns�L��8����02c�<<�"�� ��k܏�i�[��J����Y�l���xg�<ʃ\%qNyG���-����(N��+��!D�J�x����Rv�3�^i6�8�h��6�y��YX�5�$3{բ'���K,��~�xt_n<)��f���e����X03��A�<��(�p�~�4,�u�aO�i��eǤR�]�m�U��|�(�㨰08�m=�e�\�����ͷɛ�9�M�P���B�#��/�*�4?O<G~�zD�G�w7�1K9�v��5z��G����1ˊ6?���g-��uM���@�CY5��e��	�r�7�7k�q����9�����,w�H�EL*J�,���y/��6�T~l.�7�Cm���䥐��<�uo�0Cߩ�0��=	q}U�E����5��݅�5*W[�Op�\�r��|�Y%ׅ��3��`����Ɏ��
B��q~q�E_����f��N/��8�h}���I(1|X���0�mC��c��M��I�o#���ʞvw��HG@,q�C�y&g��YI�ʖ�F��{�W�y)+�1QpRA�\�|�E�Vfer��J���_0|A�t��S����[S]��h�m����l��(�������������IO@ɶ�����p�4ngW(�]�18��sy�HD�/�P:˝,|m�s⺥�z����Ƕ�d�ca��e6�uWfL�ݷ�����2ĜE��2-0�{4��7B)p�(x[���˅��Ɩ4���t{���* wy�N�~��=P����,a��y]͎o�`r���O# [ː>"a��YqC�
.<��N�K��cK�����J��(�pr�
SY�Σ5*�����!��L*7i��C��`<aT�˸���I�PJ�������x���b?�^*[0%�Ke��r���*+O�\w�O=�nd��2��
�}��rZ���:l�ҋͼZeC����b�>�p�2(=���m�n>����@��%!���ߏ.��V�
��@x�	�p�_`P$�xM��(��_N+y%�r~m#f�P�}��e���(�4(�a�ypI����T/�*��U�d�}�2V�7y�k�:��ο��_{/��3;��%������f�(�tVv_��m��I�20��>cl'�
3���ӗ3-f�b��������`y�GYN�c���^_�=���춣�)G��;��B� ��Kz�eL�ެG�3�u���d�L� �P1�z�%�;�Wd�r�M�8Ys��v�;�7$ȳ��5�4g,����� �O�c(��Y�=�������w�iz�۔���!|.���І���>�Z$&�~٫:(x�8`�k��E�*.�dL�v=ͫ����cۍKVU����y�͍)f\^���k/ժ���.!j�O|4y0��!���S�c�ݺz�����R>pK�=��L!-=A�B����r�L���{�|�2��h��@+"x��㤎h7%  p�\���t�U:Rp�.b�G���[�b�5�q���D������[�hZM�v����q��F|	���p}�!��lچ�y�ş�8 P�?h���o��OC&�>���-�_�A��`�S��)�t^�'[V��/T�ݗK=�){�0О�<<������y�9����뱵64����D��z���VT�+D\�ٺ�40SZ�^;���˳t��Б���
&��˂�
w,�z�6��}��kLlG*����t�!s�6�nI�5��ÒXC�F?<<�@Ʊ�K+�2;��Ԅ��TG?��O sYc�͢r_���D?��шĭLb'!�4#	��;�Kt�)A�S%#h%�f2��Y�R7�W�o��0\UY9��!�D~+;���@i�
#t�d�򕎷��{��)#؟LdFk�~��p��}P�T��c@�����UGm�ˌoP���30DF��L��%� F2��v�'U%Am�z�� ��b{�h 3�{����\�ͨS[�8m�����,�[D`�G�Z�E%�GA���1\�Cq�8Q��bӈr��8�;�7���ݹ�dK>�Al&=�(�t
b�H��P4�������A�[��RHZ��Q#i�0 N�,r?W�s��n��=��b ��P�lz,�)����R ��ft��$��ߛ�?�6��B/�h�!�L��̦N>l&��j���L+R�w�P�k�>�l%�:��ZLu��,�8w�V�F�7�͘��_X��(+Ȅ�g�Ų�
{��o�k��8�r��NG������pT�c��P�&rv���$Vղ�vj,,�(EZ�B*!$]f}���+���T�6M\=U�1c2�Ŀ�r�u�W����e!D3��0���0�j�oҹD�C�a��
9?BlmF����4��Ǽ�� <i�GD=��K@�
�􏓳����a�98)(�:�o�M����/�x�q̉$��gd���\�|��ܞ�F@���(��p%�����Z!v��|����Ge�� f���S��>;���̘-=4I�ם�����
r_7�,m,� ���ۉ�̳
#��:���R9��ʌB5)M��f�k�����}��8#�Y�D�sH(��QAw��n��+A�Y�~glb��9h�5�W���0U|ώ�t�n*{+�!��G�IR�n6lH��s���F�u��'�mY�j:[vxD��a�@�^�J�E�GeDˀ�.w�8��v��Q��oߓ��y"w<5�t:�B�y�/g��л���؛������/ˀ��M�s̨겧��N�~a�և��m�fO$�Ԭ�KHZ�/}e��5�-��<��QԴg ��.�%L��C_Y^ a�T�Y�_l���ٶ�j]	�{�*��\� �B=v����Y�7�@a���8f���RU7m�{��HO��0N˥�VP�F��+�Gn�y1� 1UY�u3�:�k7�^�^}��1Wt�|Ѧ��P��z&�b:k�χ;�y��w�i{�dՏ�C�שs�uh;�Ǜ�g��{���e�Z� 3���|Uq7�es�%�מz�IE����B~���4�cS�~0��6!�>�[�6N�pQs�&aw����D��M�H��{��J{�}i�z���v�l#vj�^~��3C�3E�%C�s{��0�FI��}��Cځ6H��*?$���j����ǁ�<����$��i�蟴�� A���ū��d��tXy��*A��<�I0殰7I���Y9�
������������BnX�,��UA�u���{Dj,u�f9o�����9+�VS(���@`%�p��s��]�F|9��i�� ���o�u����8�f�儽 S.dA�a;� �.ڮuD�Z���Z_cH�2*���zoi��@����[����q�%*�5;�4�Xq�T8S�\�J�j��h�P��.���v���(^��9*��sG>���`�aƻ��s���p!7Ø/�0��(�w� �[T���@�]@��� Ȕ�^��!9��_j\�ku6�4��H祈=��±	�E .N}
�pG��*0�����������V�������}&Gqqx&Qi�D�857�C�.od-���}��:���~G�����8�Ke�e~������x ��N�ڬn�:��~1�]nu�2�AI��l׸8���H�]�����ϼ�s\�_�O���ڄ����ZHava.VǮOR���ȃ�S6��`��R<g d�D(77�ө?N�-j2	�0D��E�Ɍ~�6��pA����+�d��: dV�V	����j�s���?D���]����Y{���� ����P����λ��i��jm�}��+=������M9��[i29���z��7���������MO.f�Ė��_��b���N���O��y$��hX[��$	��!�Ɛ_�@� Pg�#НS��f#m�	*����t�*�G�Ua�-��6������n]�y�UΑ�x��^xM?d�3�$n�~�+;�����$ٺ{}	JB���eN:���-�2��h���tr�Yw����0�RèK�>w��E�\��Xu��3����'wr�M��!�c�Г�YX~b�l�^�ϟk�Ԯ�#h��������M�V�D���s�M�P�Bl���$�
���i����'ha<�h�r4l��~<��d�tC��ˡ/{�}x�㍜�96�Ⱦͅ-�~,�_��YŶ�^vޟ	)|<-��6��d�g%��H���0����r��o4�dq��9�%XYE�G�Z#� _(&Mc�;�E�H�2������H�!P
��W�/V�]�{�ү�4�3�c8������e�s ���8�����7��6�R!��`�y��Ba���4�a�H�{϶@���?�:��N��WsA��Ez��)b�p��D���0O!S'�/�[�P֘U�N q�{�>��O�o94�u4_���vi�+���^3����z-���A�s�h0Y�M�q|�<��;L���ܐp��x�e�!1Ptn�`ФFe������YZ�5�A|��#��\���R��}䯿�d�\�7��|�hB���&���c�5���as#V�1���%.�'P�V���QS]j�<�&�>ұ������Ijw`��u�C&*��c�WC�*��8$B$���} ��=�GȄ�ɓ�ȍ�T�|���o�Q)��JS�ן2y�mz�K�c����N�/H�������n�	1Q�|���MMD����C���x�ӣ��*�]��4�����<�����Y�abVx_��L���F-���syX��=��~���Zi;��=�'��+c?��\�fe�؃����~r:ɫ��vê���_�~Sfe${M4B���rWH:���,w�|గ<�6z1��9��� �cK8�A���>$;�`���^���7"bd8�ܽ1L����.�ז����ࣟ����!M�N��O��ؗ���!�p���2#>�+�p0�}��0�P�!o8*�؈>8��Z��d�o��=p�����T�i�����_�IO���=8w, �\Bk�>`���̿��؎T��RY��>��Ts��["��9S�q������`�ۖ_��y���H��
�W-���-V�l
YQ$W���^�j埒Sݦ�����=�B�M���՝KLƷ7�\y!<�c@���V�c�w����.xp�ArC����#���ڞ�u�-�>���f���}HD�;�SHL���j6��NQ��#�_��D�L�!
�;Ŵ���w/�_��w���OM���x',!+K��/X.��'省66�F�l�Ұ�A����fo���
�!=ؑl��~�(�k	&P��J�������n���QSc}��F�"��(&��S�7��h���J:8��u�^=�ς͇kuⲆ!�[A�����	~̡P�Õ�G��A?�,!?괈��%Վ.���OZ���]�J��q�x
l�VZl0qσ��DW-ҾpEH΃՘���k���/�!H��i�|�}
�s��K]Ԩ���a��ݳ�Q%�x��J��R6����wA��>6�S���~�Hyo���L��߭�?���%hݹ���)�Iv��e��Zzd�o�x7����,HI�0��-�v�[�����d�&j�R?�Gj*�r90�sGYƸOʗcw�8�����b��y2��M�/z��dx�n��\gYTҬ��C���f�|m(���h���<7�t}<�	�V���"�Q�N�f���W�_���^�Y��|���ls�c�)j�6���٣ۇ��P�۲9sΕ�v�m�u[9������p��aY4g?V�n��m�vx�j d��.�љ����PSFeJ� �~�x)xq��N�LD�i�F�q�Z���?��!��"�4�^�J����N����m�sz���/~ Ǒ7KQ�8�_�-�_���ݘ$�L�ʾ�V�!�D�6?d�Y�㞑y�t�C�n_��ݳ�1���T�SͦV��2*�G2ױ��^�z	ӊ"�[�����ɫby�"�f�t�f��_-mU���O��`�[)�2V�V\�r4��A�%��x�E�-�����,�+7�'�F�=�1�?L6e7�d���ș��So���:�#M}<Ht�H]�̙pW�����| �Ǉ�mM��|�T�5����&1��?t�:�Yi�q�i������b+ш�OA��7������ �YW'���T�ú8~n���M|	���g�.�!B�8�����ף����{���3ག~oj2&��D��{�@���ͩ�g:�r�Aث�7���ª�M����=�n[Q��1�3��湜$l�o��[ ��C&�������4w � &&d��+}��]�����
����}�#�]Ӫ�D�����4��Y��SQ��Gik�m��-����[�=�v��b\'k�eTe���į���X��~�IQA1g����xjP{������@�G:�T��k�<#���ű�\s"����T��>�o�C� �q���j�v��3C�
��e�k~�bGLW72*7Z,�����3pH�p���MI�K�>H�v6	ja@]�H�9��U��3m���¥��(K���,�����P��9�/��)�L�����r��&xԧ�]-"���=ٓ[u1F�Y�	|�T���~$�.>�ɤ�6��R��X�a��z-�I��B.�dp��/���7�S�;%��|��d9�l�̤�r�NRXޘne���`Yj����͇cI��uu(*���]����s
s�'xt�!�cW�J��m��ϸ�i$�m��ǽ��E�bwn�ކp/!�2NT�%ITR���A�űϝ��� ��=Κ�� ���#K�l�	7�%�ua�vW���ks�}�l��T��g�D7��:�KԻ|�Z[�6�fR����(;�e�e�]�3�OE|����E�L� ^��c���V\��\��.e#g*�y9��]�_g4�𓏤���dV�3��U��pf{���J!�4u��fW	�'b#��`-�&�43H��X�� ����yz��3���R̀���J$Ȯh�_@a?F�n����M�K8�
^/@�<���1�I=6v��������2>� ����ŌI}Tٻ	M^!E~��>O�>?�i̱xseDX$��^��8�3�~/<�R�B��t�����к�ܢ�����u�F�U�f�Pc zVt�{{o�b/�]���V�z�9\�ߋjx�lE�����=0� &񱲗�b�����j��Ň|���{�*�3�d�BX������������p��n8��٦AGo�ˍ���>��ĩ��̸cu�%�P|_j@�N1R��k쓄��N�zϱQJ׭M-\�\$��)��p�aʟ��*�q��$-�+����� �Dv��J�ũ60�tK�֤�QǛ�J%�i����~b@��D�_j,O�s8�y�iu�G?��7cXh�:i��iq?�9?LE���y�$_7���|+�畖��`!<d�j��Y�'&ju�x+�����j�I치�����=��#�|j�e��>�>
���ٞ_ ��}s��F鐗�&&`O�py��!ە
Y��RN��b�w��3�Rd5SB.[GQ��z#?��7�:�y���]5�@j�Zoq��J���`�� �	EIu0��JA�k��6_��h��m��<�Z)��9��N=;�R�+�L�Tf��~��I%3|�5��_��r.j1��j�ݱ��� ���}aζ����$���*VƁ }K����A���=츘��u͢P�ѳ[�oC�V�X�`/�$D��_ysHe��f���=���Q�t]�|7x���\6���"�|��;^���$�%]v��Ά�B���'NV���_9mr-c<�p(�-�v������C�����p�\��ހΦ��%AN�k���5�췥��B�����֍�wn�#�4�u\P��NVT*+�^�²�,�*�	����:"HtK^6�aj�Ƭ�\5{�U�eGޚ�	yv<g����Kz>2Xqm��7p�)JFg�~&���L�$S���*Ts\5�Z�L��0�U˻�w(G�d�wBg�F/��r�6�45Nܠ�Ĉεk@�����j��)�1���m]��$]���ev�o����@3��ky�����q3Sn��n#x�R}-�����$��#���ޥ��sjVy�5�:�l�ݦ�>߯;}
�!�������c�G�q`HbY������i5)H\�#�'�g�:R�*&��3�M&N[��$���&�C<��]��t~1�@�Bܠ�%S*�BϏ��3���2^�\S�m��xN����о�c�L �@|�)��e個�608fU�����'��TzkMȴ,�����i��Q�?I���tJ�-��UE(�|BMksҭO7`Y.�6�b>)��X1�z=�۬��̕��Вkp�"��.�N��a|��;سԾ?ڥ�%�M�M�<����Q;��ݭkj���]�&�ౖf�@�?��Q<ڤr�D)�d
̭^j������$Q��2W+�d[L�ZAdb�e$����GM�3�VM��������6q��>đ�ȵ�=����7�˽}{���BL�jc8���G�~V��J��T�шH� _��z��-L��f���6�N�2n�ݧ�3���#���t����,�����_w�,��}�Z���a���@fJ�"fK�~ˁ"�!�F���7ce��^�(k0��YИg�=-�dc��Ք�!�8���C�m�f�Q*��F��Ʋ��#iwOjZ���?���Je�AV��fٝ��D�|:��Q7�zż���M-�Q�XBde���`�s7����{��[���'�)V��-W+
�Z6�쯽i��¨RI��k*��\fק�)�"�ْ�)Xw�|6S�.���X{���k2i[�99?� ��Xθ�vĲ����k�8c��,j"�(3*î+����w�Y�fv5��ae��z=˷zc�ܼ�B�e8\��M��9:t�K�;�R̉r��2�蟡i�[Q��d�����M�%ʞK��X������kOX�F�ve^C�C�!Ƈ$��j��B��+���S�e�!U
�	R�{-z�8�q�M)��������R��e[��T�4g���JO���F��5�P[�����@��4���Χ�א���&�Z�_Έ�u��g;����;A�kN{�߲���� ś�����Bٰ�n|c7H\��;Aߝ����S�$�~L2������H�_�`�H����^颹4؞��a�B؏ �����C���)W1��	����Q;�T�J�֦���6p�B�h��fzV��hj{*߄�ʓ�a)��bg0�,�0@�-W/�]S�ٶ��,y�����3tكAl����n���="�	됒/�o���+���ΖD�e�aڍ�X���@m�z�T6<s]ͦ��j�Gw¥鸙�0�ˁŶՊ2�f��&�D��ɮޒJùg�S�A| Z���7�]�[�  9%��n����4�˛l>�?��[m�!��%l�2/���u���q[�j�4�A�hGQ}}l��f�����ݯ���t�ذ��0jZ�;�j(L��a���5kpL��[J�D[�q�H�Sk���������{Q�!*�Pr�6��:vh�R��~ׁo�q�.L���f�����J|�i��@�҈!���Z}-ž@-��%�E0%�e�ȋ��2�p(��ێ����} �m�k�Dy�P�n��δcP���&�|s(�(��A�8A����	j����B���&��A�d�?����`�v���2X�e��hG:�Uێ��9�Hc��!��F���	Ɩ�w����IЎ���eK�TDiOn�N�h�G5��/��Ѭճ�=�s�����۹�iҤ�&I����`E�K�u1��8Vu}��v�2꾵x�%�����Gaw�dN}�y���]	l��E���v�PW"������V�����i�@N��:�˃*[d�^2kI�ʄ+�bO*r�s���B�D�$}{��7�&���Dg�#T1n$T8�JĻ���g�|~YJ>g;���^<*}Sx�J���7����f09���u�$�t� !!��l�� Y�	��H�1�Y(M�g�PCiY7��O���R�#�������(#c
ydv�Ob��ݬ�=)U�q���n��� �L\K��ނب�)��:�y�KQ�OP�B�}�[�C���z2P�����=���߂�vC������tbu6J��g���e��⌰	_Έft��Rh
�s���M�p^����B�[��ш�`f0�pθX��%�w�L�*9<�1���3�Aq�"���D�:�k�PΥ`��P@��ܲH���,��Ip� =���p�H[ͽ��������*
 Qj�2��;��l̽b��yN磷ء��������	y�?�nG�<�P�����*�uH���9��3�\�Z�l��B�ISH�\v4!ڳ)����R�0��l�y!yi��-g�L�~��>�����k�l�k�^LXі@�K����	��6��Jȴ�h2�`�>�������Q�.yqThT�1�����_��z\��}�/�
��T~3�_$��ww���{��W˖�ﰍ!�֖�B�=>�Pn�l�f[YfM.�"�V��-�"e*(B���ܿ�l�t/�T�|X���sk��7�T�Tj��8�H&�ظ���:��k�3.����C~r�	����%���w���n���itz`Q]��	��dSV�#jQ�$y�M�ػ�EK�.R ����#����o5���e�A��!<8��qPG�DV#S�*��9��\A�	*��\��V�[��e����Kʓ5	��tn�J��1|�i�'�$=���-�+5-�U��J��5�0{��x�G*��ہ�m�f�iQ��ƒ�r�\��0��(�Q�g���U�dkt'.�.5����
�������k�����AS0�sʑ6�ڛ�>���Cg���AގTPE�k��/���6 NI�w�M-W�2�]J�+@���b�OD��_� ��*��4eeT�t�̫��w:*0T�I,�_uN_%xC��u��9g5��YJT��h��LPg�[���1��>���c��J'�8����T���UNj��GG
�V���} ��{ NV7�KL�R٤d��MI���2�@VM���mra�����7�MY��c[s�	�Cl`�"#$�E�q����H�a �rZՑ����̐H�n�� xֶJ�11�Ѱ�~�L|vO��Lh�i��N9�ʻ_��=��0͚_�>��;O��'�*H��y�ŝ���%ԛ"�,�d����/1��0�~qJ�H�"±�k��O�>Fm�Tf��v~�'�F.�rcl:y	<Pݎ�
���Y7��RP����U3U����3�Q�D����bA��iU�W����v=��C�F� -#�\�Z����`��l�2
D��`��T��1�@�CD��Y���*�M����%����og�~{�c���)����G0=���'���6�j'�+(���NM�)�����'���K�{.��fZ%&8��䄤I���'�6�PH�!˼��՘��?��d�=�%�&�)0�GA%L�˥d�1x?~�[���0��U!Po5�D�0/*J����=��N�Gڨ�H�T�u��c���Ze1m�.G��"X:���J�jYMSУ}/ԛ��fm��DY�k���+�끓i���O�E��Jaz+̸��n�{y�l�jw"�4�����;�`�� �Ҕ#�H�Dؔ��s��D��'%3O	&���$�ģ8_�|<��R�]+�'�̃���������i�L�.�Q��o�E�v>���:7&�6��Gc��` �E���#��a�]���ŵ���,0pA�= W���FN�k2
�@��s��`Il荩�Y��&�WꀓbWb-��'���sh�kj�b� ���'տtQI�����D��,�a���D2Y�2dz�J)�<�8ZO�')v�ig���[nU�~D>ӥ"ٚ�a7h��li9 j��:12�J b�l������|_���v�D���� ��0���&�0:��)<��5B3:Khkm����W�q����?�j�.1��Vi8���n�%�(�f�@"tzb�8K�xT����ۥ��O�J�,��<!ҼW�3GF�<�����%?��V�&�V8�P��$́�Qɷ�4+��U�ǒ8��X椗Co���O�\�8���Nh�!O��u�#�Qm�ȷ/�}zl���~�j=���`r�w�}G�*d��*��	���/��M���'��2��.B�^8�{[G�71Ǥ�op�����Q]��E�q��{ɖ��o\�#�%&a�pB[�d$��[�]�ȁX�t����qg྘����Q�����bTXz��zуh�C�Zu�O^����ʮ�l��W�$����׆?��Hf�C°����d�fת��%tY}�g@�o�O^C��I��V�O�flH�^^e&�w��`
��]���=�df!/Q+��_���m�ki~�V�5�������S%o~���K�<�_k^��#�7�Pj��MN�eD%_(\`�;��h���|��.��?��Z�eJi4�0eOĀ�ۏ�uG!K�>W�Z8��t���G��!� ��-�C27���G/���!���6�ܶ7�&5ڇ�uC;�o�x5�s��?�z��-�h�,�p]n���an�C��=b���D)�w?Pp�z%�H8�Z������H�Y����D��77��?R�|� zq���z��|��K����������<;�8��o]�1xg�~|�EtVó�W�-傋�!lem�`k�,�@9�	�r�2)f��|Lr�`'Ϥ�zt�++`1fˆ�>y��PU�\{rc\��~���c����Q�J���?H�w�DcK��*�(�gR��M���
f�g`�鏤Z�7v�-� FP���;�H��`Mi��E0��Pk7����E����(~͢("�ɋ������'�x��)}�b~�ٳܷe�mz��p�DT�_]x]b{���ʋ���+��Ϭ�N�]�x�R���D�"�QlBcd�ܖHt$��y�������F��Ăbi��g��D��$�<:R�N!�h`E�E]u�H����>,�!��J�=66,s�b!�Js'�p"!˥�|��Np&t��{l>Lb9�JӶ��1�_����VzI�.х��g��Ct�)×��  |�;�h���`��R=(_�Y�.*�~6�n���B��A�c:0��ۻ�������ha�sm%���A4�&�����N�yc�C�:�*�^q�kfP��lG�kG��������`H��߄��Y�c��L�<���t8�A�r�&f���#���.]h�*倝���mA�=��>���lFA������R�:���ŦJs$��M��\���C��6���Gӽ��$�s_�����ਗ���Nw��]5�XV����+��[f�.��m�/@�M���',��8���d��$v� ՆS�����%9L��6 ��1�w���l�>aZ������v��v��ɗ�`�ÀS�G3�����@#}��c��,Z��܊�0hH�%l�&)`Z/��/���)9�ǡ�W~�׾�D���J�߅����U���D��&#�t�0��Ӧ�	��òi� �i: ym�r+��'��jX�/�K��1M����^�j�r��E��9n�ܺ�ƈ��Q`��0��Ԧ	�P��8jq�pt�ߔ8�B@�+i��?��Ƌ��&-�S�?�~������r��J�t\�u���j�|K���Fa�_�h\Eb�ؼc)I�q�V�B�ir��L�[�n���*Jt@v\F`
R��W���(�w-��=���v�����@U4�!���rd>��c�4��|�5�j�p����ɰSG
�;g�+t/��m��>���迼�E���J��������D7�‿�D�+Q���Jal]��ǉ��̹;�F�l�d�., 4w�F�-��H$T��/���#��j�֤>�A^9wox�5��q��h� ���Qk}�Ob8S�i����=�ri�_?�#���r���1��n[r-A~�#���OU0��v=����zd��!S`��w��62�R3���H$�_�ғDcq'mY�"N:��X	mho�R�^�\}`+�F���~�9 �[�xp��A�;��/�_�[�N����9�Z$h�/1��	���9�*]��5���C���}�IR=�R?
a��D�ic���mfj�[Yl�@����2O����)�J�4�h#_,�a�>[d��I�O]���/�z��tk�=�] K|&R �����BX��*�D݅]�����^�V����-C�t�T�o$��<��8$��Р���t�d9V�!�
�d�d޽��Po4�ݓg��������`ș�?��0Ȕ�Z:���T5E��¢ʸ�U �qD����f�R(8�[�ׄ5/���qy�Cl򤫩�@�ud������'�I��^�Q������f`\��o�(�i8�v��,t�)d1�Tr`�3�*<��-�J���%�6/TYOPU̗i��b�����6M�XB����/�i�b�{�ף���.�d���V�u�^�+�z%��l��A�W�U����H��X�����ڬw��e�`�<k���c������䎺<��E����G����95p��2��.���̮o��מ!_g�0[������qW�9Z�:��ܑ��N9�3*ĕs�X9 !���w¼$��#�x%�$��%�au$a/8�l�U�ʠ��dd+�2A։��5㶮�*%����Մ��`,��{\���2���@	���1J�z\����1�4Z��f�B,�KRO
��o�)�W n�'ؒ��>���bW�AK	7֛�u ��n6�D���d�
`�.�䦛�TRrP�`�C����4�(]&��~���m��.3�C�����KA[��Ԡp�J4T#����&�˻�g��^��3?:�u���p��+Mu�zI�IY�T�7]��l��\���qG��S��a
<����}�-��eL�.\�����	���I��`jίh�^d	�����8�~��Pe��og��td�Ε[ՊΈ ��j�u��͊OH�nP�ĊX�`ˎ���(�ka]�LIuDhTrX!�9�;E��-�d4��U�qj\B�H
�1Kj��&Wu�)�P����!�Ws�y�t�(��y�%��M�~�����X=� �Ei-����+�j���Z�'�����S�]6��:$.���*�/�N{�%����d��D�b5O�{��w`Ο�/g�����?-�)k򖈰���y	A�G*�=�Ĉ�������	�RFZ.,1��yY�<1��j]D�ۖW�Pw����TI<g�in���[��~_��^�Js���	`H"�;s��+�veqĆv)����P��E�g�S��ܟ6ߚR��Wu8~P��j�K�s �#=yq_��)�+$���+.B�*�R-в�����<xcw1��}7U3)��c����d tj(o�5 �Ri.�𖇡�r+E�b[�Y���P���d'/Y�.�C��3��0�;u�����,�/���)2�|�^l7���L�[r5�u�=���\=V���
�{���Ҝ+�����
��(@q�?��%c"�~�pt�a����}���Adw��v�}p0`���'�j3֨/g��T11�z访��zݳ�����jM�Lm��T:������@���h���uz�@_�>�Q����B4��A��J���)����\���A��b�'N�J�>��ꬻ�=|Ͱ=�^%k��~�4�J?���1	9r3N^��$��NבB�&��s�	�#Q��hI<�h��$/q��Q݇��9e�Z��^�`�{[�QȘ�bT��<��1��BgM���Ct�Ar\&�.v28��/�$��y��1�@�J�5������3��좁��S��BP(h9���g��9������JN' �FV�O��X�p�F~(]g���v�B�c��2����0��󶿉�0�zZ����W�[P5y�	Kj0�k8w��,�����Ԧ�|�����>�s�r�e1��p!�@��ẞ��Į
/`UL�X�'���,���et��e��K�߯���ΐ�2����\��D���;�ґ֮�*��|�U���xB�����rL���$��nm�1B��xPG��>����"�P
��jo¸�h����B�4��_anT��ǖ�Se?+� �]Z�@Wd�ߐl+�=t�[ �kS�H9&\�o�2
��0`%�~}-]���)C��J�J&~x����Dߔx2!P�~{#�'�;'o�//��Ly�{�]��6���Y��m�Z���u�����;����u��C�+�0�=�:*��@ej�41���sPq��A�Z�#������IO�H���|�$���p�y|ͣ����!fRק�Ce�L ,��~hk;c|�rt���ґ�L�77ax�����0y�$������G6=�J-j�xn9O��{9̢Y^�Pz��Q
����s�-N�tg��&��Au����\ӓ�l^��,�F�O�:�I1�[�^�]+��;koٛVN_���A��"�c	7N��m�-fJ�R����4`�z1)��G���7@�U6�BE��F���^c�e�!ӂ��l��B���N�eF���;i���]���[΍5ᅃ��:QA��M�X�ׁ�C���|�LKƯ	]&M��H�|���r:�4���䝯wh��(����P�j,R���0x�EA/�����[B�4�ˉ�;_%޾|2I����ͮ~-��~�����^��-�����+�`z��1�ߛO�g�QgB�Ϋ]Ё�E2��c�C�C,:��[���1�]#��8�#�-���_=�5K,����>!�T}B�Tɫ�a��O��/hØK�j�=�v<M✏��e`&24x�St���$�w��g�W�<�I�VI�Ƽz���,M��Ѝ�z��}O�OmϽ}�7�����W�����+�M��4��M�V����#���D�{O4&��s�}z��b�\a� W�tb��]	�]� e�Y3QU���u�жh��I��W]�ʽ5As���̝��T���т�c���[�-r*���D��M*�۷�MWFQiho�#];�B����YX�`T	HFg+ܠ�j]�&�s��RQ8�`�*3E�|8��ӏӐo/��o��dy�5t�.��0�ICG�Ҟ��<_��q`�[��}�@nwZ}�xD�@u�2�K�,�v�M�{�R���:�t���n��H�H�-B���&�_7��n��5L��E��!V 4zO�w�k"��ԇ��a괢 yO	��1<#���&��F��P���㤯��[���|�F�:�i��D�)��F���k�C�I�=ٗ25/+��Ԓ��S�E�Q�gȝ~�$�H��LU�o��g��ymyz�w��T?a���0�칢j�ߵ��0~C�γ�홗��NrT��+CPz�JG�I�oġϷǱ�O��6k�D ��`��Uj��g��B�
�8^1 飖����|�s&�������}�̸%ueE"Vެ�0�ūq2-&��!+����s����� �]
"�G���oa���Q���-8�YZ3���?�ш�3��%-ْ[�ҙ5-�����`58ʐ|��M��Ӽ7������E$�d 521��.����g� ֧��O������N��6iW�G�v4�ut���i%�
��9����P��[�ն8xS�;���Z�dUGTK���o�kbS���b}�
���o|��Q��ų`�ļ�{?�Qg�_���WC=-Ӑ��|ڗ,�#r5��J�g�%��vS֩ �+~8ф}��wٷ|e���YD&��`�L%���i2ۚ�~��$@Pu���ȝ��uX�^q,P�<G���>{�y@嵼����6�'�Er?�m�Fo�g���&fA�	�b�:*D�'}��	Ƀ�Q�.gn7�����v=�<'�kE�|D4^Cۯ�M��c�r���9���B�w��"�B�G�r{�E|��6���\n�aY�B�Tad�6��P�$/���;���{t��V�mv��\�Z���@��w�4�<e;)v�¨{ގ#to³4��Z|ԙ�Imm׬fc��׈��ڠG�dO���*teG�T�l�{=�"��{�f�!S,/Ѝ?a ��,���-���1R�q��6q�KA)�Q��T9!=��.��o�ް��Є�����B���K� &C>��73a-�-V�~�,�G0�Yrf�����B�e��\FSo�̆��n.�vT�Ȝ��B��#<�r��0�_l�L�7�6��]�Ɏ�����/ϋ��_a��4�N�8K���T�Y����eHҥ�E>/��k�NpXj�x��Έ(�����r������l��N��Y˾F����\b�.ϑ��z���YO0��Q"o��Tb.�0T�Bi!��
��V!�YrO��u�7;"x��Kg�$����{�}�)aV8���^!a�?�g5`�
_�r�wT�����kv�S[aPϔ�����F�)"��o+m���J�#�Z7���e�@t��扻d�������/�]2l/0��Mh,�T��t���{<4Nz��QR*�j���V�A�=(D�[�}?���n�u�
Osb�D���0��/�b��+�Y�B�b�)�� ��W����Di�.2��qh)����5�2�� $��5�^]jĄR��N[Be�%൤�H1�8ҙFs�d��c$�c�
����4��Ȇ�k�
��~��H�$�p��`��.0%���(���9�>�V�t
�w��`t�I�q��������R$�����'��J�
�sP1�E�Ҥ>T�x�����,�ؚf��VxGz��F�N�wFE�M`���\�2 �?��>H��K|ͤЁ5�o��~w�@���;qQ���?����0()^�/��W���̯�V��tҪ �V�#��1������ZBvG	-K�Ӷ���h��_YUd������0XLo�Y�F+�Q��e�y�A�`��%�"��@>�a���wA����v�N�-5�%z�8�zaMa�ΨF�lvvjy|1�6^4S^1��}��F�t�~���<�����O�y�g�jm�3��܆����^��J?��Q���A���|.��B�#'�t!��i8x��=nrw��8���3��� ��U���:h2�6
{1 �d Û�q��+�2�$�X�v)3�}V��f���X#�4�3��O^���"޴1EF�[��S�����q�^-�NUC��s����f��\��{��$�:JZ�-,Gm�2��/�&�!��P_�A%�Y��� � ��=�XM��pp�khB�:�'��\����/���#Po(���G��<a*~ge���H��!���v�iX6a�N���"[3M���W��mK�t�OK�xv�cus�{Z����nS��;�;t v�������C�A�̲ڜ��!�_T���A�B�[eG+�C�mE���>qB�#�ۏ$�����3��=A��l{���n��L��*��E~: ǥ�$�a�"(
w�O�wz��\��Γ��T?��K1���	��x�.�N="��l@N�TP@�3����NK��,�KJiم���Į7mғ��6�����F'�>�O��OPB T:�k5�-��vZ�C�`|Ԋ�6�A��W6Ɍ �$�F�&���Ӷ`�J��m ��)C�m�'�ȓ�8��j	�hT���QH�P㯹W������}�<c-��p���.��4�]�q3������r�҅� /�x\2:H��n4�F�fwV"$�M����2v�v���"x������+�sm*s��✬ m��!m&�K�6��ǐC|iy_�,$Q��a?�4j����B��]��g�j�H�E�)b�;�1�q6n�+i�ڪ#��)xO�m��]�*m�ahZ��J֡U�y9��?ق�eĆ���٘��&T+����d�b}����ۨ["�i��Ԥ?4xі�����l����z���fl�#��Q��L��z��c)��O�����oT�J�!�/�������= oe2썼�Ќ��Xn~²���>���� s�p�����3������������j;� �� {!�i��6��;,�؃"k?-\<�-<�f1��~���A3(�A^~�9~}��G�B�Z�4V��sI��O5$�
h�T�I����o����SR���h�ª�D����E�&�O&�$���[��xyʏ�#k�.�V�ul*�ە��k��u�:v=���M�#\Tl�{�
�CR�~@	{�vQWF�d!����
X���J��*�܃�~�$c��e�O��:�΃o��.H��t`�+2�J$�AJ�����sڈ�h@ϑ�4/���&�-�Y��S�X���V=�V���r��Ԟqqx-�/H�-��ax�Tڴ�����D��,.��MI�ޛI7�?:�7�Z�=4�;Q��J�=�����{�vѶI��x��"����G�J7I�#ZI4�O�<�ٖ���t��������#�h�G�Q�;-����'
�3�-�K�KS�(2h^(�c�A�+���P�,ˊ4��G��\
�-_�r��Ԭګ�Q&H�T4jh��HD �+�4�iv����F��f?����D�h��O�z1V�d��UL�˩������:Ƒ
A�~��N�Ds�x2�;MP9����z�>BT��-�u��}��76!�������Ag�2͆7�w��PN��x��l1�������E�tf�1#�������.j�)С ��R�{�BW3�����j�4PF=�Y��O�n*^���6�j��-z6���։���n����k�0�-]ц��r�p��K�-F~y�K������^(�}��M�"+s�������~�|>t�.�^�|s-����!r��&u��>��}Dj"�)�`'�^����WG��#���+lw���Z�a�!E"�uI2�=a4� k���=�O}ԩ%�;���Z�Wp6Ds	?`~/��Y[�+�0s`[����4�GJ|RH�����`Dw?D��'���Q�$V��f�F�X+��e󁐙�*r*��/ົ+ujz���4z=�"�Bu1�dr��O^���Y���)�1O+jU��e��K���ق !��p�yf�/�  ���v-�!"�Ő<��p��h��e�_��+yV��VL������q�������/�]+���9�*w���i��P��U*�/9`[����g���y�g�0�~QT���v��'���#tb����e�?���/�L�9�7��h�ک�T�2�	 �~_-�����m��+�OW+�h�"�*ʇ%V_�s ��X���5Xay��r�d�!���94���k>x�i7��o���"��{Kh��n�p����!*��\j�3;)��N\�^��=�=ܢ(��>���s��%���	�^�5�?���ާt���d&S~���7O�x'd#�,��]�Y%Ҝ�;��?�n�{�'�a�h���p�3jjײ&�CH�]����A�R�KU�N{{��Z'y%��]x��Tt�!��(Vu_�TeP�1<[��ܙ����ڠ;�P�b��@OeY ���y��T��z���T)��k�VM�b�f�C�NM{u�:���1sy�:j%�`t�����g)�~4�g�|���-�y.p���E~�.{n��C����ر�_E?+<z>���t����>Y?�b���5M�1U�'Re�H.*�x���y�`��u0�$$�#���9�z�>Ӫ}O�T��76�;�y�PZ{�H �c��8��b����ƽ~�o}���j���Cv�Ф�j�&���d��[���w�����T_��=3��r4�VX����,^�)�O%/�d����o<���R������7[ķ|zŅ��wZ�Tݭ��X���W9�dl�$��oJz
��)�u�x)4=�.r��X���m�������E�Ǉ0������㇖o0ޑ�Mu2�h���ͷ.�l��њ��,u�!7/:Ǩ����qx�Y�3O?x��I�R��Ao�SMLI߇v�kRP��c�^�h�(�F��L��0�j��C��������#��Wt�'��J�?�]���}$t9Y�_��u��cX��:��B���j�7W��%
�֛�\�p�N ϱ&���o$�ʑ�joOcͤ���o'��\���,�XۺH��<NI�$�[���g��V��/B�xC��,T�H���>�O�9�R��� �x����EW�u~�5n�p����������mx�\_e���!� Q�*�]ǌJ�I�*���>�_�Y�V�e��Q=���#4`6v6�����%�%��� X1%��͟=�A�ڦ���6�	�_�%��!��wUk�:{ 
��!�cc{���`�(]�=�p�S~Yz>#���i�pW���L�����[Jʧ6�4 0�9>*�=H��V�x� ����q/p1N-�A��[x���I��bt��e姠W�r~�v���΁�ӂ��=b�ߏ�d��rFc.�*8V� z����K�|�6&	�L��>�W^	�1mr" ٬5��-�x�|�@�s7faa��d��kN��W�O�	p�ח>qqW'�3��%�a��-7��/!Z)�g�i���'�h�U2h�^;zO�C�\:�L$�]Ks���M����/¿�-�v�y���-�֩H��$G�ޢ��w���#>��I@���崃]�c�WH͓:3T�!�e��x_���s���nѴc��FBH?���7Ijr�����Y(hq�`�.:��_��ּ&���ZP�OP-���qq��� ���$P���T�`��2��
�F
˙\E��a���!���c�v�1�z�Lc0����n��B �\'8�� ��ɏ���k�� Y��~��(��1�� �Lag�mό�h=��T�S?��=L�e���Mdj�X�r�v��3r���!os��ͦ�~�r|�M�t×fxa���7޲�(1�h�X��^Ǟ�8>�L.���\����~��'�Ş�i��c�=J�5O�"�2��Ls
����D�.���'R�ݨG9�0��m�����hy�~}�������L<$�&Yv�	�����RG���)#��u1O&�ш]�^�������i:�J�\�](� kA��}'*���s]����b�
�B�f����ч�<�7�27f��S'E؄��k\Z�v#��H��Εs�7sϔ�_mҸ���v��N�a�#�� �WS�p����&���]w�>7<�Hs�����,������=�ή���
5q��}#m��
����ƭW�ŞZ�ܝ�0�םp�|�БK2r���lqB��C��ֿv�(1{}�cl��߾���LW�,8�<�r���F�sp<���B]�H����F)DD��KK��"�_b��ٳ~�&9F�e�� I�V/=��Z����\+|@��>�����=�WU����I��,c������U��HR��A<���o�N+W�q%�zŁ��U�ُg�䷥�cQ�f-�=́����b�(;6L�����qv�(4��"삘�T_��nѳ����H$'��)vbHF��S6�����T|ҝ�����f�D��q.O'Sϗ�wO�rV�;#ΰ����5c��x�D���O�r�U�lS5���>Ǟ�:&h��aPHm��M�uA���d���x�k�	+���%+{6�Y�L�Wb�I�I�S���u�±eƬ��@⥵w{����#�#������>0{W�ϓ��ѿ0��Pɩ\-�^Γ�����8m�dR��oL;�:���[QzO~���Gɉ#�{��ѫU�'�}H�p�"�y7A)}���62i�ȴ@��t�˒f�>�0^��ǵ"ͭ��?�>s�(?��]���O�ϸIk�M�@rZ��鍖�m��<+3�<}�*�
y�`�:
�5%�i"�n�e�����jRY��Rk��{?q�M�6v�)����$
�BB{/�^�T�]6�uzOSH�: /�=$=�dN�&#��=E����ߺr!K�V�:��/̏Y��K(H-}&T�����!:���ē'ݼc~r��	'�Ɂ���^������u�vm����`ЌPw�8Y������cH���FF�%ف���u�EP]��X���0+�,���f� ���c����ѕA(��S����8�W�e��Qг|f�?@!�T���p�v�����a3\v����&1�ov�X�jw|<��j�o`Z΁�:|�9Jm��;6z��dMKmgYb�	�s�b���Y ��yy�CE��\fԿ�9������阝�Z^�l�.��h@0�Z:B>����f{�\� �]�I`I�N��;���54��I�NYR"�K�1H�^�J��n�6�t�Q�s�E-�	��m���zJ��*�X�%�B]�J�!to��>Ă����@F��������7ʞ13#��擩����ٝ�}��(H�;V���$����U����d+���]��� ���"��ԙT<��|r�BN��$�w[m�����������9�`D��*r1�=������
]+q]$VC��[1�F�K���z����Q�����מ��G>�7D���E��n�d��>���!ED�F�M����2 �hK�5Z]���pT*Mr:]Qg���k�8�������Pȱ��5����Y8�-RYw��8��^��3q�q~!�$�o��K���d�/���� {�Ps�ŕ=Y
o2�-�.@9�Z`��u0�Qy\X�e(A�����(���ЌvG�*��:
��sNh+V\�� �U3VzKyN���^z 	Ď��^t�/������H5���s�a@u�͗L:��;u��t�� �� �W&�T��]�b���Xv��8
}�&rh�R�����c���2c��_��DX�S�{�&�����������SP{m//��x��UEi:�p/Nɧnk�7$bil�s>�]o�}H	��ƌ���{B����i\�c���uf��f2�ȓ�DK��$Y��Ɋ�L��U>'�W�~Q���O#7!Uu�ee-��9UR[˞!� 0#�V4��u����:�U�+��{�̯����G)m��%��{yi(�Q���xa��ݗ��Y&���x���\t@�����AͰC��.lt���~�S�6�?��D������P\�� �B[g���פ&�^�Td�Z�]W,xح�_���#[y��������M��{�UK�J|�7:�_ݞ@r3�y'���<��.Zf�ư�C�n�����L멸r�9R���F]���F�KvJ���C��G��#>����˙���lȞ�5-�}v9,\I=��v#E�>���O(q�ʢl�ZN3�&�4|D������׮���)�T��a3��C��)��'�8Z��Ob�d�z;R��a^��('h�u��џ] ���|%%�z(�g|I��}��M�.4%�'m���ʽ-�Wm5Z5��YeB�5���'�Ҫ����m�J�B V15�AAߘ�r=	��I�xCFgK�#�=k#�5���[�?H�b8 E�օw���%�ĩZH��&�X�rOl=r���!@����	�eJ�U'�l����^�lَ���]��?@�~���p5�b��I���*֜7���y�{�<��ڛ�A����X+S��f}�Q
gU�<0K�M�>���p��C���h�n�?d��&V�3x`C�}"576����[ ��e�r���ȼ]����g?Ղ �43ǫsm=+�=@������KfaA��C��2�yl�5�?�ù�I�ϧ��\ƒ��~��z�r�7 =<ҕ���lK���sbQ��h��$Ԍ��R���Z�sV��x��^9��'�9Tu�Ύѣe!��F�s4��Ty��I�.1����`3'H"N;������oU*���I���сğ�]pzD_�'�>����n4wn���O����4q���`�6�k��&�[���o��%����l�w��QTh�}*�ηQ�+��1�0�@a^M�>���{�nF:h�qm @����}�kf�Cp�u��
U�-+����|��D���K���~��e�uDO���hĴ��6��;Fe,����1�-��C�����4HJ���G��5��bi�ܔ�R�WcqK\0H��;�}��[��>уI�"��v��ё-��19��������j�*��$.|>F��i#�?�-���%���	P����d��J���S�$�O=N�Z_q�J����S���M�;snz�a�.2�h���R༝��b�FL`ؑY�x�ǧ�������#���p*�~���q-7Lu�i�P�"<�n��^T�>�n�5���o��^����p�(�>a��r��W[Jr�}o�X�@La�h�7BU�ry7��}#���H��3��_�<�K�����Y��oQB�V����9�E�]r�z���zȑvN:=+���w�3������/�e�h�mCCD�Ci��,t[V�e�y��r���'�ٙg1�7�h�R8�N���j��a�O��E�����=���48�1�z6:�E�u}ӽ�yZJ�VHF�Z����3�Ѣ>�����<W
X�q�f����=�#�:{���S*6�ƥ���eb�X�3@4�e'���� �luWe�W>�;ݖp�L5��`�H%G�L��c�RS������p���|4S4���*3]�pd2ͧP�ӈ�L��{�N��0��c~N�f(�i��%�l�[���ܔC��{Ɣx^1�������ٲԅ��fW��0="gM�hĈ��"���M��\���]c[;JN�wԬ.�L����{�����%`���ɏ�
���6����:Y͸c�b�16�w|��9&�����9�G1=�}D$C�YFM�N�G�q�������z�s�$z�}ꍚ��Tn���w��� ^nml����5�`Tu�/�T\�H1����YF8?�$����tG�9��Xy��O��=>����}�2x������u.�*
�T��uտ0J�o��g+��z
G��JV74�c��x18��nl�X�r��'m��+�]�3j܍��_�e:�i��8�c��.:"$��t�ް�������h���P@��)t�����G闳j���(�~�j�~sM,D��:��Ԅ*�\��n�����<�e�|\�����j7�zlY���7�/%���s�X޲��G��wyEwC��p�h�צ�Ӊ�=���H�C�8zFjD+,�%� $�).@�i���x?�35��-\�}��aV�-��\%�*�m�����3FW�W�e�YJ�XC��XQ�2����Z7JbϷ�	r)���M�8>�FtZ�"��^@���dc�� <*b+:&�|��R嶺|��(HD���p��YT^�[�da6��ܕJ���uW"�Y��;�����(kР~����W�?�s�(;�����Eԝ�u��yˆ�7��_�z*��I*�|~K���f'�+��zSt^��d2�w�e��W^e����+�{���C�*ЮL�%��T��޷��|��i��r�{�DȮ�C��K��rR��R2L����R�6��1��� ;����߉w����z��>�9��g��o����B"�3��?3�|���X�)�\�ռ�u`����#���\D@�"r܌�T���[�Cx���?��F �����B�/>� i�IM&I(�-����j�*f"J̒����/Ĳ/�z����h	����!!� �I���ݳ~��N��W����kp+�%�]v͆�T�,w=��w�M��b�����`����C�4�-"��=lx��i�1���ɍv)7q~4-2��T8�8����6�Ͱ��o��'�%T��ClЛo�K���{^������J��~��.���R證�E�ܓ��2�da�ˇ�F
d�l���ȢP�4=ϬG���)����T~rϠ[��n\1�C�G.��M=i�Fb�n���5�?��_���hi�
am[�$^)�;[��p�!`�/�Q+AS>}�y��Q�WI���H^u�K�2�D��ۀe��s�����E�雌�U'�&[s��^
dL�������s�$G�ݷu.] ���2���~��DF��`ԣ1�0�R��Nų��\Bt�b���d���cxG��޻�"i1�R愴�uy��'0j�(��R����ZZ���)����,5~����Q��>��E($50����F��g���F�L�6���+Q�eͺ���:�����g�و���UdX��@fS���s><�J��B&:����R�=?G�\ͦy���9lݸ���	ރ��8����U�	ߟA�bK�0�(3��"���-�G�_'߁/<MEб��:���=�/�����m��� �ػ�`s`��&��^=I���H=�;�a8�=^��ǘ���B�(7�"��(�z���[rP~cN����_j_�-���C���O�N�#-���q.�|�ݼ\`p���~��dZ:u��W�pyRN'M:n���4����Q�X?{��Ѹ&\H��2��P��3�ȸ�ǻ���y�c���Χ��v;OT:j����"B�6�eB>3�jA����I��"�������1Z5��rp�.��C=fpa�}Y����m�Q;Y0���'��떪�NȊJ�&�↭0R�i;?�2*���ݴ��y�2�6�o�-���}��rڙ�墯ޗ�}�<���퍙�^'JlXRn��F��̈D���0�]�+��A[iP��x�3�,#K�� ͺP�&�B�Mm3�'c��3����6��:��Jȍۮ$ePA��`��N�C�kE�S?�M�h>*�Y��v%PaG�&�].o̎s�u��-{*#A��K45������U}�@.r^���N������b��Wx�]6��U��a�ٝG�`G�g'{f��	)P���U�&[�*��i&cƠ ���`��}�T�{���(^�&�(q�\�'L���^���d�Bc��;�� ���0p�1���w��#�J|��݌6�V]�G���fY�Ȩ�F�uT�=Ư�DTF�m�������Cm����i m�5Xr�"oY#��]RR��GMke4����8�L�y��$���]�MV����K'!�F�|�;��.�y�Oˤ�{�X��dNN�_��lM�5��>���(	W��c:�%t��C�>巂z�B���[.�b`�UӰ���""���=��ȅ���,�SPH. Rq�О�C�� �`�n_���S��rd1M����BQ�x��|�~�Y{�s��{�
�޶iV��o{m�Y�c��033����^�x��(q= 
{���%�
&�����/{Ȧ����+�M������	YN��qi뛉�ZUꗐUrYhk�┺p��z��#�1��*�Nk��&�:��>9F�n�)$�e�jn�ʭ�D��H�G>��a��q��j��͘S��G���=�/�(ʙ���w�<��ǧ� �y`�Z|�c��ˡA}�(>*6B���!��Q]s�'\�&�k
	��%�r�SvF=�����M�dy����.��b/�H�S�0�CޮP��fy��@�N|�XSx/� JA�jĂs�F<�N�U4���w�G�}�ǹ��s=R�([>�� qǁ�k��n��h������x�0V0bqhro�u���n�I>�͞9���}]����K���}($a�w�*Q�È�o���u��2�@�H�$c�C�[�"�����QD���ݹ�NX�	b8g�l9l��/��z�[����P�Qz�UK�Hy���6����>���+m�������~����c��	=�nT �w���ea	[7uʴ�����^\��?;�A̋J8�a:�T*��=P`	�i��J#;2��!}�1*�У}�^5| ��#":��Wc~A�<^ԟ�C�{�n58 #����˶���fR~5?}�؎H��{�A?��8�=�܋�*���W�&�CiؑV�x�gH�-8`>�"4�10%*�)�k��-�p�R7¢,C��
�%����Cj��^m"�zd��%+��x����ءL�Iy�Tx���o1Ͳǟ��!��w,!@:���"wÿ7v��G�8Gv�s5i�� H���T���Մ���۶�(�}���*�N�4�|�$�!~�+���pO	��J��w����1�����iT�\Cf���_di5��!�h�Rz��Z�Cg��i�:�-�3�Z�b��|��P:�~d����Z���'�[��OH,E� lgcH?~.��NP��rܑ�MZ��f���w�!�"�K�/H���(���RP�$J._�i�vD�6�ҁ�:E8�G��Uo��}�����Ct�{�i��>��(:Q��l��Ih0��\K�y	l��k���M<�]TU�D�B��ޟ��c��(H|x.o��֪9�_ WFw�XY���_�f�m�Z�l����f��J{��/m%� w�^JEY��A�q�CG� �U�	�9n�o-SF%��K��	�Ojm�MG�rZ �����8t�9F�/�f)��E>M�wz�*h�Y����P�>=FR��PI ���5eD�F�%��f�^�ml�t�	=�כ� ��-���6���nq뀥H)�w�Iܡ
MA?A	�2ֳ��%'z�� RG�Ң�M��Z�]�y���Ep�*����9w��]jBo5��� Hh��麮��0�*�*9�����,�τ�:�wO���W�ʯ�s�8T	$��| �¨�o^�2��m7�T��b�(�\��=u�6�k�Lj��S���,%y�h��=�3�oq�}�8uT���+�>��3�u��,���

��cMs�ު��4����
N����n�����3\vvr	յ����Ϣ��.@g��Fo��Ljt�ϾQ\�
k�4���G���t�O�z�21�)�(Y��'��~��&���� �� Q5�����������uֵ:t�5�K�� ݳ�X��F+Ce:=�Fs���Z�_��p:�:7<����K"���`V"��蕉5� �V�S��]��`��j
-r�}�"��$�JULH|�$��v +!����Q��R�$�he�P����݆�J|<�&�:Q�'����qZ]{Ta�p��{�Jǜo��/<ȓ�D�#��{���s]�U�����ҚU!^4l
Q��/����,���#�v�d+����)7�뤵V��c(U�g6+Ds��.�M� ˧B�ׁ�F�\mO۲�~W6�w��ِ�S�7y�=��y!©OWJ�k^y:v�v>�VkF�5@��:�Q���z�p #i��GYg�T��"fP�̅���������Kq��� ����(��[���n���&Ġs�c�t�������T�"p�K�|H��D�F'�rh�Q�0��3g��ư���.u]�L
}���T��@��-Eh��z��T{	^��M�)�Wꅈ�f��!1��G��b\T�H)3�o�{6��V	�?��#��X(,�@48j���(nq�CK:%=����~�D��ޡ�!��L�T؁��V"��	�O���Ƿʖ�=[��5啶��1i`���o���M\��Ӭk(c�����|���i�[�F[7,��jT�mzݓ��=��C^����� ��TFS���u.�P%�=�x]�|�3�FmU�����Z�q��������:C8{::��ON,�2��,T-�$��>���P
��U�Ui>K��_G2r��%~��K���L�H�G�j��<���|�i?�����l�A�C���?ϒ��Bw�Z���3[�m�s�b�T��d&��lގI^� SM��:��.w�x��G���%H�)�K�,ʮ�dq���PJR0�[
�"�E���5@���
�[ ��z(�]'��H.y9ns#U͂!q�V�5l��ņp�ѧ�?���AnK��'-!M��~�eQQ �Ue��<W��v���%\�܆��S�W�ݣ��I��m`eǳZ)�U�|*��{��&����=�h��m�y���܌��U���/���k ���T�I��|�JYT��+Rr�B��/9�%�؄w"�G��^y���%���c�� ��X�2(���)�,|��cp�3���[�Z�����&ot�E�8�~��!�~���7<bہ
�_@���w�54�����l�a��&QsS�A#<���K�.�JJ�5��/����-�mթ��f0�)&�(��5M�/&Ú���F���ھ�0�SR�vD���ȆV����~
���˷�k]�u�p�C�2��;���������+?q	��F��a��l=��s�&�4�o',O.�+#r���akY��0��Q�z�Qa�	���Ĺ(�$��f[z��'����}DmbM���P����UK��~�.˂�h!�1�0"��t�y��<I����f�<G�j�C�l���f�Jt�!�剴��4�h���m���5h�_�����k2F�(Wo�V�6�~lg%*���HMt>�"�uv'[ȵ;�y[n6b���Z���MoM�q�K"s�)~�f���*�@F�Ӳ&���A}���9�(ãvBm��Q���0��3��e��4OiA�$iУgY׍gbl�	0h��ȩ��٤�l�Ue{(k���q��u\k8�8���]S1�$�?_?���:N�?��{e�M���d{����@=7�7ΫF�7����'�]����'�K9+����j��;�6N��ip�3@E�TBU��C��O3���b��G��gRo,���;�)���It\ﰰ��'��,�"��Lr�L�4#228WD��YÔ�F5(�]/��r�lS�L�'�����ļ7C��A��]?��7E�Bl�_�I�o80�g�zg�6�;E	$*���ю����Rq1��`�� ��ْ�ٗ�{B�Ш��ej�rV�JcBЀQ�K�ҼI���U����}#�i�N��5$��Z��0Q�JH:|9n���s������|�*@9}�gu��l�P�Z�`���,Xr�Y�C~S-�Sn%�N ����ל���Vp9�K��"���3�|��nG\I��%���v-Cu�� ؜���,@/�#Hp\��R����ġ���W�T�ϔ�.�''�^D�������m�?X�d�9^�������YY�Jd�:*7 ���Jx��+�k�1���9�ŊC�l�ɫ|A4�S��/�OX�� �Ӥ�-ߨ����UՓofe.�Y�(�9�/�}�>�?@�#��4���坵#��ЏpR��1��n��ٯ