��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k�;_�>6Hl������t��Z�$ �G�g�Q-8V�6�������S"�"�M7�ꈾ%g��^� q�ۃO/:��[f:�'֒�%1pLP�~����;n�Y�o TS�ꄣ���n���/�H��CW/�Q�Y��ҿ^8�K��m?�t�gm6%��>{fY���>�Y���Xuj�$i�MG`��  ����k��L�L<��Hǿe�o4�Y(2��Y65�'tǠe+�I5�:�&� ��N�<���4���U��J
��� ���D��e�.8�[ū�Р�,#�U?VQO��8i���O��*XոU�\l����c��g�6���b�9��l�~���״m I0 U�5���/J�{~�p�j]l���|C�"��S�&NQ�"y���M�[������z&����v�J駜pR�k;u�>�(������[d Xwon_i|��mE;j�ǯ�r�q�j0Ө0=�bA%&�-M�|�N��ߛ>�¶���T3~��u��Ѿ����勲r�K�n�On1S������OO(�������ػ-}K���N��2&?�g����!�����e�':�o xբ�&�N����k��p����Hݠ6�ũ ޘ�cT�,������
�\�\d�9f6Y�΍�l��(gTm�r�FK�<��}������`?I�Lw�͟�(�G�C5�}!��U�ݹ�E]��^o$䀅�"zoh/U��rK��uG�1s�[��G�+����9Ί{(����E����>����a3�o�wC	����į�z�u"��`SX��c���h	)\��N�I���;�2�;wu/���u�:���YN*����^��I����vٗm]Jd0�9'@Ī���>�NB��j)��6��0�m�X�m*��y������_.h��sD�a9�Pp+�~m[2#���.,����7zG�k�c����77�b��k����"�]���/�%u@Q;n:�P+U�����I�U�v����ʀ1�SJ�����2aS�ڡ1d!r9��J2%�5s�R���sL_��@��Cz�i�c��i�K��+��H%��Q����غ#���y��EC���MSb�R��S#��%7���n2� ���鼅�ʵ���XR�O��K��N&���ޑ�����-"�����/��~�$4�K�|> F}���w�ȴq[� �v�ȑ���*ᘅdAv�{������B6��P��_�9Vy8h0�ӧ]�&�E��0�,xM����J福��V��]�Q��`�z$r�ˌ4���Ғ�����)M���Ӊ��ߪ��M9s\��ʱp#}{ٹ� �ix���3/?MbD��Sb����c���i�y+��Ң�����s2^F \:g3L��ƶ�������#_D��:�T��
vP�r�b�L��Pݹ wlf�^1=<����2;�~��B�W�&Nd�Wڥ�	�-	�=�5\�4���ύN@n[_��M�F�/o�sY�X(j��y�	�x
�B�El�����Dd.{�)���#adI��E��v?g��7��j�.73q�
��)GJ��)`e�	|M��姳
X�o���O�	$��C�s���V��LX����r�DΎ*c��{���`>�#o��:��0)8��}*�1`P���'�ɏ��8���s����b3�T��s�����v�Re��'�$Z��I���b��Pʅ�#���ƈE�]H�T�!ѥb��$����ן�Y1z"EB/���m�
f y!�D�Z�|{Y��P��Ě$�-�+F!4D����aSv�[��L�_Iܬ�L��fP�l`��A2T�d�'g�,ιl�\y� Q�Uvk�:�n�c�%�2����I�|�}&x#�$���([��/P-L_`]W�h$vR<��sJ�n6%��Cs�q��"�_�V�>�aS8��|�PsL{1}�5��=g:zoa���V)����d�<�z!�1���1�K+�1n��yMѦF�w�d|M����H�ŉ��v�dI�׀M��9t =��^����@�#�������K�)��$�b��!z3�$m{~Y�lqG<H�Q�LZ�_������3�'���n�J�l 	�Մj��,%���,�U �<��H/��>T2x�(zJ���+��� 괛��[��#��.���5��U%��e*ϗsҵ,�+�NHj G��]l�����G�����Ś�a*�_A�$�.�b"��wh��?��K%��]��*J��5t����)��^�R+�P�M�FhNZ�Z�`O��tK�B~P���r@��NpW	:8�d�(�����:H~<]=`QQ5����czha�x�)h���/e|d�C"�d���@ؽW����:��Л��T�2�?��+�)�OM/�]%vD����&��~H���v�'��Sp	�
���7��̌?�V��j�V90�[�j��
B'�e!mr�+�|�y%T������o����,���r�*M��cen�	�kJ����T׎�=��x�}�2I�:�����r1\#��K�������-o������pҤՋw�נX�����rN�:�����q(��p���Բ���
w:HS���G� �E�<���i�W��
����]ޯ����D�I�WLS��=7��u����{3W,��׳c�	��ka�|$f����e�c�p���	��`B� ���1��L��cM������T_͢a�����	]�*l�~V�_['z�q�viu��������?��lO��܇�VA���+��m�^>&��aB|�nK^Ll�P�I��چ���Eu�3F��L��{p�k/d���}�Rz��XvȘ�������Ba3M����v[?�����8&[����Y�XuS}&�Q����K��:^0I�K�]�}�����COv�w���q��͇e���#]��m���o��eF���"�\��j�Z��١��(��z�|�W��<���bt咧�����fT1���Hoc����V��_�.�Ս��!�Lkn��ή�U�@o�k�<����uF��c^3�~��E�ш]��_7�3%��\��U�E�×97���J��]y�@ǁ���}0�=���h�b�}`�c�w5�	�F}�F����V�BF�
������D���f����|�86D�N�}�����Ł8`�� _����0����ȿ������B�)e!���(�,���E��j��MKtN,��j���'.U�|�애-���SfF�d�M(��b	 ����K�H��=Z�j}{���vT�3��|��w��q��b���	&����yJ��}1l����a>5G�dF5y	gW(��T4��٭W��
��%(����R����p�)I��cO�ʦ�R!���e�d v�r|���)B�T�d�"�~B�c2�D�V#?[~�͟?y,���5��
3��WV�W�Ĥgq��H�g�~L5��w[�|kߒJ�}��*9�K�� BC�V�D�}�ގG[�nKs�(bel�b��Dd �Ux��1'~�{ޥl����@x&Q;��:Ez���b�L�+ҽ9X(V}L��b���� S��������_e�r��Q���Y�~q9�11Xxb#� �r$'&W��K#�-�y/G�;ـ�!��|֭��p>��i]n�*�P�[56�����ص'�yF��,�w�v(����`�7���
ϟ���R���@��Y�r��`IO=�����!j|غ6��p����*f�R��S� 0(ģ��i�T��
	v�
�p�o;��|�:���n�o8 W(�%�C���I�/On-;�1pG/ �-�ߚDXx���?+�j�^	��znވ�[� �XM�ñ�Z�c- ��妮�/h���,KY3��c�gY���~�\�)P- ��ȶ<�����Ho���d\�ئ��!Ub��&y�O?nү�f�c�O��uR�^��u�]��.G2gXtcbXr�:��l���{�&��#�n˚��+���R��UWvȨ^;n�G�Lq�����X1�8�f-������B��@�l�lM&�.��?�����&j����qOH��?��m�d�}NK�������[��#;����mN|�l��,�Nm�s߼Ե�5�9�7�ؽB߹cB��X��!L��4'� X��49G���& <�1�JIg��W��9@/f�է������}��Z� �T�0=|�n֐���@�ϻ��A/F����w���w�G�k�4=
�y�ha�R��+2T]���.K7�S��X�Š:7�|�؆v��{z`�JE�[ki"/B蚸ݟ��;�G7&L�(�~S���$�v��"%�1�U������	����J¬ܹ��SaЋ��������]�S�n�,�G*�e@�J�"X/��vQ�ZuI���]U�Y;ø��⼑[+��>�]�dg^P����e�3w�n�p��>X-��*�QILD&VHb�e�?� �*��.sﺆ���Hl}������ �8S������N=X���r~5U�&�G>�sV�`�Jv{5�H����[�#�bp��4̚�©��eC���De���3��14����5]�9D�m3�g(������I�bhb6��J����#����wqYp�`��6�e
��s�婪���q� �Y|�y������0~�=w�c���$���0l�q9�����a~Ä��K9�}/�,84��tz�/��? ��"���|��޹�^�2�}]�m�c�z-����]V �h�o�Y鐃�Ƃ�w��e�>����t����wl,`�y��4Eϰ)��R��q;���b�jKK)��'�Oߊ�f�&�X��d�17W�ΐ~44}�D� 8m����r_Q4;��Ð,p���+�R���������{�Q� i�("!(��$��0��_Dt�-��CV�8r�ӵ�����'����2��W �W8C"3�=�RA7�ތ���$������e��ōd�z�b��;���n 5U��E$A�GE���&�+n��{^t*DU�Eiė$qf]�Fܓˡ�� ٛ->���Jwht���� ޅ���&`�HyXZ_= 򦸽��~���`7uic���.#�+��4��K�檠�R���UTY�\*�
I�hN\��{�B����e9�F��<���f�u����N,e�a��ο�Dt��gN��󕤱w|x1z,)w�7��������W�I >��F�����j��n)!��h-��Mb��9į	��J,�;�6�Gi]!�4'�Z������I;��#l��s��t��;��Ry@l���~�}�m.�Q��9��WCR�����|p�E���H�l��x�Sr�$[r�_��֒G
P�O}G�D����]�/��G��A�0��0q�`��HB��$:���qS�7�V�"�h�K�NP�*u�z>�c��2�y��SN�b�͙&}��z�͑5qT��e6�y��.u��^�Ħ��PwMY�S�C.��H�B�t�:����4�lJ|>��*/X����J�X�\wod���7%g��)\�t�]c̚v��[�ѩj�3ZP)���L������.
�]>��u���A
fU��m�z�n0�ݮ25�GY�C��T���b&y*T�&)H���F4��1�ǷCH�33���@�Te/��&@K��$-E�}3��xA�ݓ�����6��-��əv��>1�X�7�ć�2�H!�ZM;`��d��ML]I ��q��sMl�)ou�Fx:��+'��ոq���T�n	����u��������dq���^p�#�ʯx��t�zː�[E������˂����+tR���
�5����}��3��HI,xL,���"��#S�����&�VL���>*4�|\ͫ+����!E=����[x��~����VSZ9H�<���Q���o�E�f���Kj� r=7�-F/I�#e��\�G^�cv�EKlA�e����FR�c�E��[��ax�*R�'�{�D,�x��MNJ=1��T����&@׈r�9���q�����6�wk��i GM��R���Dp��C!���Y½}j��v{I�i$os��;�����reѺ�O��`&�x�R�(���J���t(���?��?)�`;�Ą��0Ƴcp"`�D;����ǡ��oT�ժ����e�����A~�q$�U�]d�ʇ��$�,U����G���t��p��OO*���
8>�*A��y���U�P �b!�����<:��q���-�4q>���P���e*�
=m���
D��:�V�7���/��!n�c|N
�c�+�PZg>):k1+մk� Ꜷ��݋f�����N�ӛ�jw��rs���ՇSa3o�P���)�7���n��b���ƒ������8�wi��݆������#f�o1�C:������-7@�>,7�A3�V~�ݤr�ׇ��� \h�e��/g�-��y��;�h��&]׬�B[�N�p�~�-~̆�v��G�n��"�csL�6W~�^�^�:ױ�xQ�~U�1�sk�).-	@W�Lkط�n)�J�H��0̷�e���2�?X�eL�t*#�2���w�%=���K]x�̉��~��-�J��������NB��lx�8�vr�{T�H�&ۅ��m1����)�vx�;�4&�砹�hHY��Ĺ�>���v�&X�9�~���A`]RA��âMguP����Z���7�hK㕑i~iF*o���0'��B
���V����eiK�O��F�ǀ��*)Bf-ϯ8'&bϦ�IA��,�<����Y[��{�]g>}k`fo r:|L�qA�����(�l��B�$ތ�ڔ��$l�q��Ĺ���g��12��xfJe��Xnv8<P���A���u
6'����Un4�s��$`O�@&�J�22�ғ2X�G��)otH�"7Ҥ�����AF�AC�ۼUw���ͥ{b�u�M�:�������W?�V�Q"����{�xe�P� ����]�����̱zM�,a�{8�f.��3W#U'�< V7�y���S�[��1�D��觻�2V��Z��^�@W����7`��U&��|�9�
�A=vZJ-�A2w#o"��Na�ixԨ�L�	��V"}�����s��NS���B�����.Dk��7G^<w����sxu�¸��ɯ ���C��AG�[�����>��Us�������K�\�"CQ{ �'�lc�gK�k^@%}��tJ���F-7k�|�ٛ{zC�}^���JV�b��^\ѱ�ǐHV�u�6�e�����(��n�݅��\�C�j	��aMk�.��hH/�X�� ���X�y�T^c�)�`ܧb=$��n����1�V�!�:���1)ey�?E-��K�;��6C�D��{�=U(��c�7���it���l�]4�M�f'�p8��d���x�e�K4"�wU�{Ǻ�Sk?��蜽��ۊ
��	��I�#w��\lJג�l]=eq�zٙɕ�6��.}»�|X����>���q|�#q����x�������*����<봁�z:�|�]/ʹ����͟�2���sK��i������.���,��"|mA`b���a���~�H��[��pD��b;b3b��w�S�f�Pٻ�W����ċA�H{�-cN_=���j������S�uϫNy���V��w���23�h)@�nʓOV��^�.�����s[�Y�|D�����
όҤ:s�|]�O/X��r#�tC�z�eb���3�5�v��)�i$�aqz�3�SZ�X27��r#�����j�% n ѩ*��(�}3��fb֙����G�	�['&�h��|�������":�f��o����-.�H�sʏ�*�����D��	ͷ�*<�e���[�:'Z��!�U�`6��W�J�Ԋ���p��H!&�F��������B�zD�#�vSŗ��t�З`���̿,�s ���7r������(:m�=��bo�)�;��*���ae4ph$]�6��;�:u�=�C�d��=DEK;H��vu#���I���Q%��������i^|���m���P)�hX���MO����z� �f��Oupy~�JsX �;h�ܕ�!��}x���O�$ ��w����`�MƳ���EC��~I��V.K�N5`�w=	��nT��۞���h�IR"�y���Cv��8��OP_�v����:�J�@��9Y�]k��+؆�ֶZ���E��}��PZ\�ě�� aʭ-1c�	1G�E�kX�i��|�UM�1��E�Nߪ/��{�=��G���|ʷv|v ���'�NAw���vK)O��	d��{��5gS�f`[���A�hH�6m���b��Yơ���@��������]l,=(E^��hl�8=S)��x��F�r���+N��C��rƞ�|�N'���v��X��Y�p����d�����X�s��O�&JA�Z���^�G��Oz`�����:!�e-�< �ڐ-�R�HXJ� ෤"��]�*�ظ�v'�~�,GO��9�{i��z�֝z�Z<\$��$�Z��)s~��~\'I%]z�iP�sB5�U�#���Ll!F�#��;���{\��C]�����l���0��zs��;b�ƕ�>1a�`���=_��aZ'!���[r�,�����|h�%m�pb]��/��,+U��i� ���
vFe`v���O�Z�2�#�&��*b��]h�+�p��py��q�|%�[��*�S��A0�ھD����_4�꘲ �qA�f�hi!r-�t�U �1��.4���f�cs#0#�ƸE0á�(�p�Tۊk���у ���E�3��u�$�>�@���EZ4�f
%ș�:H��G��Jj�����{�������133|��t�aQ;����F��>�1#q�.d�S�0ñw\�΃��PV�p��+ݚ���L�������v�Z�f\�|�hD��F�� "��[��z��(��B>��l��^*}�o"M:����3GT��B3ѣ0�_vK�8�)�a�\�F�_��t۠���Ho�-�K������]�KS�M?�%~+�t`y1^Jf����4��D`Q��1m"�9��|�i*��{@�s��i�,�3�e��y��\h�w-�啯��{ti�Ɋe����t�k4�2'-����M�K	�k!4�Z�?{SpI�M�O��W���d�ܖ
˿<�	��Htl���mΒ-3D8��m��r=�i���V���ѣ�W_\g��#�%A��4;uo�hL)$����Q���m��������i�0c�kq�\��@*?+y�9m�u�@�̕��ȈU'��P�0y���jd�0T
���
�V\�:l1���3U-rs�#���4 �X�c	Ɖ0�^�+_x8���o8��wAr��ڞQ�=I=n���zÂ�Tw�|{���&SSR���,���k��(Nk,"��P��8�W�2��sQŽ��2q��ԟ��`\�%Rml��C�&���Ps/�dۑ� �$k3��M|��8��Z���_���S~���u�O�W�V�~]e��1�Ǭ*ĄG��q�Bl���DH��hA�Q���g��`�F�юDG���5�uߠg��}Gսt�ݴ���j	`v�/���~1�}�8��+�3��=��K[��9�o�l��;Zz%��0 �y��쌠@k���GN"O@�<���7�����A�Yu�E>��F�Z��<�}3����_�'�:2��^o���{?h�*�$G������e�y����������E����2��O��d�Ѫ�|��	k��� �JޟS�L� , .񄥒ɿzK<4�AjĒD�x���u��u��NT��M����~?��ү�>�a�O��V�����Ɲ&��k��|JvI��97��x�9Of�G`~ojv�L*;�B�澨Vi��(ڈ\.`Ӝ�)����K��gx�p���B��8�g1=`AZ�G�c6B������a�s��:��7;I!e^8~��E5�5%&�N�����u�Cx������#��J�4>,�r1�!�T@:�,j�U�n���J�i8����&��qu�-�26�v=���?�"���8g��O�ȤY׳��*p/�uA��n	�k����|,�T�NOm����ɦN�.MPߨE�d�&0������*ۮ(���9�$.G׼���&I~������]?w�Z�͐���3��`c����ٕ�[�u߂�N�]2��԰���!3�k����d�@�j�)í�-�⪣rC�oj�M�5�1�i��MS��4Ɗw�5C;t�"J�}^9+>��/���ʒ�I3^aܮ��Ȓo�Bl�i���_!vTy��9�u�ݣt�ͷ�.3�b��]`<<�<�|�O�����~Z���k�di�|+�u(Ա����䶤5+��X\9GY<SMPb�3KV�F�v�|}��X�j,+�[��.(������p,�)�����t���iB���j�Rg\�{}n�#��If�"#4�%
jٽ?�xGC���j��q)Kz�=YN>�QIp�?n�C�Ż>@��������C��nŷL�'v��b �c�Q�݊�i�ld.�_��� �)�^� :�������@ Q���j�Ȉ�|�p?�8���H�|`��{f��䊖��ն�y��n��w���gۂ%\wAvt�x�S$8aU��[6gaA�@��K�� ����ז�p�ɟ���Hjv�9���VLu��!b=7� ˋ����o����V�Q/�e�?ɮ�^ ����eF���F�^I�����  gu�+eZ�y��M�6���N1`��-�s|Y�@�u ����Z�c��gŁ#���7���K�rf���G��![�W�ͥ���rPஉ"�i��� ���\�0*�qSr�����4��	2E��@�Q�`~zjIO�c,s�2^�≗ڧ�_��?�r&$��ny�LQ�`A�l(G�L.��y)�MG���Eױ;tpZ�Z�����5/-�ު(�t�d��C�hÉid�dQ��To.�	�̛�ьtL��N��M:����H@��z�G�Ö�<o��:Z����݆��Ʃ<I�r�u  K�� �җ��om�աU�z"���p<�~0�_IB"�׈"�g�>�����G���Hz6����ا�(���Q����o�3�hQ��0I���(ӳ��d�0}_y�#˜G[��3
Q��KW�	��ad�`}�X5�At��DGI/�LO�盀��G�+������`���b�*ھSm��w���^��>H��1.�"�$��~ԓ�%����'������s�T�@f��hc��T���q�:�i5��GD���.V�JKvr�M��G����D��~�9�ˬF���5���7��E8��><��CtK�qX?��~�W��F
�+ni4��Ͻ�q H;�znN"��,܃V�5�&��LY�%�-�������w��h!z��GI.<�6|H��+�E�>�k��`��&�P�?!�.cۚ���{J�bvn�����`br�c�H�w��$��3���#�Q�j�Dmx�)p��o��q&�H��bu=z+ɯ1aJ��0ywsN��QO����y#}���V4S��9�l� ���[�ʇ�L{a�"����-����'^nγ'�]fK"|u��2M��e�A����M��"D*bmW�d	݂J!�BrE����$m�<�m�fj��з-ra{�Έ����A�1L$F
">����م��bp�@R}+}��{L����4�Hjc��7#K�z��%�z5�)�<�K��u
���jv��@8��J�*�
�%y>憫פ�բ�ޤx|�f��fG&��QEV)GQ��+����D7^���
�*�ƣ�k-�K�kq$����6׭�#�P�r~�A�S��4o i�� �s����ǜ́+7�_ۜ��ׯ�NYY��;5�Q��@��#�1�Fy�&�{�"C����܇�B��,_$��JV��{4��c=+�N�����qYS�*c�1�Y^���E���Ѫ�	��HG��9��@��\�}[�Y~�>%�'Qv�ѧ7sg��@o�����-s��Z�<�������CыIƤqĳ���km�Y�J\D��U9�������0���7�A.���A���Z3�-?2/�0r��s����%+�-��g�bE�sc؊��ѐ�J�/�Fc��<��؊��s(����Թs��"J((��g	q�5E�MXT��\'~�D��ۆ��":B��yY�ׇ�
�Pz�g't���Lk�|D!��Mf������������"ʶ����g3ꄓeã!��Q��䁷��(<�y+<UA�P#���Q0�$�Ϸ��_�H���rm�g?w�ˉn�$�BOu$��-:�2��+�vA�z�3����N�M"��O-l����'�K�Ő��jo������m۲�Բ��sS��C��T�����H
����h�W��K�؍%���������ngRM��=�pHu�A�c���E��	�7�t\l$ȱ���$���3�Ou�/�Qz��1���c����XZ�������Λ��T�Q��kSMr�9�Q�kRW§��q�����7��ѡ�q��1M^�{t<��k!��I
s�,�ώ��~���ƙ�I��E�y�U=ՠ�ʤ׺�+Ӎ`�ǒ"{�[ǩD0k4bv������"���lڝ�@l�����6��˽>�o�q"�FH�:�^!��%�Z��6�x�Y����%L�<����$S��M�^��9qYY'��.�$�0l nk=,;���_�:���r|*�.���@CU�ֵV֍����&9��Y��E�;J.;4rbscrm�E�[^j�w������C�m��&�
�_��W��LZ��Ú3 1�	�9Ls%@R���/��p|�� ���\��#6�x�Y��Tg���j��vi���L��y���kt�"����؛J�WTܫ���� �銟؊��E��8k�ՖsU��g�3�49�����2N������[����,]-��L�cGE�@ht}աT<�,���zK=�$��AO�A�섚�p?�}X���
��%M!�.�`|��:��IW�j��<�W�S>���о�oG��E6'����������üSmL�!12�VDGpF�0ɴ�'�KRJ��r�6���&����f���"AG����>װv�|�H�e�8��l��4ȩFy���Z�B��(�����(�/EO�~�t̠��C�D���E�;���<l#)�����?��>�Z���lrΏ�@`C�F���J��r��@�;�X<.Y6�Ȏ`Xq' ��kb��*��Ŀ�����%��jBѶ�ٌ1�%�y�ΏJ��I�Hl&����7T���)w]�[����/�����!m!S�Bj�%";���^"�5���)$�a�f�b�B�<���X�F��?Y<���AԌ�"Bd�P�Y�V��LOE��`Q����2��B8�XRĞ��kd@��9�C�iǓnՉ����i��,�o���`R���G��6Z�?q����8ew���f�xh4g�/[��Le7:���4J�[e��dzh�a��k��(
[%�;�5Y�Zo����{]h7Ak�"o��)j��F���Z>�`�F8A&�O����I�!M��/h��J��O����Q�n?#7&G+ۤ;)M���<�g�?�� Z��'�u�\��W���ơ�)Xo'<��2�O§�A������W�"����@��x��q���Q�ě�yp��������\<�
�L���Q��7m�
*f�/�NB����گ��xP�Qe�u�!�(�C5L��'!��'L׷�N���]���]h�l�5��s��1��R�:SHV	�[�Q��0����9w���]v���,��t�ZC�>]�B2\�C����屙EAt�?�m�\����[è��b�l�|EI��*�_���xf�È�W�&r�l$�ߌ>K�r2 tLW�~4�O�q�*�y�̋����Qg��aT2�>�$�0ײ:�D�u/�U�b�ߑ�K�ZtkE�b7��gqb� [ZDRL_+����P?�J��:="֭�`���V�D�=hM5�j�GEx��~]:��]��R���)xx~�4����to��_HC�V���'�<2�px�b-�ĵ�2bC��ެ�oe )�q�R��=
u�AU�˖i+��X��j��ŢG�;|�A��\��k7�᳾�L��O�Jc���AK<v�Y�I�����~#Q�Me����`��5Y ߳����X%=�(Y� ~�'K�g�f�F�	C���n<L��_�.՟�*���bn��㣷EP�Њ������I��Z��gɟ��X�/�$��C|���x%*���q��DRL��bqC3�E�����{ƮUߨ���/K|�~���N�cTr� ��O+���yY�&hڇ�a+��	4��������و���0�w�qpXf�@�\��4a�磱yu�� �:�X|��fv��7���dU-�.H�`|=��=+ilD.�҄�23���31�Jr�TO��$��_� �:|Y���G4]Q�he~�T��t2Y��!{ʘ�$9��ݸ7=W��|���<w�A\���n?��z���2���-,T)��Q���ٴo���3���2��q�=��W2`QX.�SK�,�א�:�Y��L��e!b���k7GR���]]�|ۭQ�u��:��y�?���G�P&�.�ny� ��43�Ew�uOU[w7IsHr����>�������< 'h���i:UX���o|�#���ɪ�u�Rǩ� ��B����CI;?���̨@��A�Fۅh���}�Y���B>`_u/�'p�^|��v�W�k�F9,�w9�.�B�)�B�驴���һxY����'�a~)�r���{�����I
�����p�X0]G��u����+جHIц��tFn�9s ���y����ۈ�:`7[���6�7'uV���f�dg���c���D��4�Q~�?�P/�Ȥ���}n[l��~F痮Tq����t�� H��CN���� �K���Z�H�.��$d��1o&��Pc���ɇ�L>�OHL��~��-K�ìuS3�`���⣩����W6�?��Z�mڮqP�e��bH�,[G75��8�w�'A�ׅ�$�j��,q���U��Ht�/��X�T-Ak��E�8�2�/HxI�#b�(x���6�	޸q�=D#�2ڻ��b�KTu��ڇ���Ђ��
V�׺Ҝ�{\�X�c]}֙ڈ��?��G�w�%v�����c6��|�^{V�afz��#�*�]U�U(��V�#���v�N�&���S�X����P若���~�B�zF]8��m������O����Qew2D�x�p&j��8���&�rA7���-[̜�㛴��R�"��P�|���]����u��E�&� t#��t�����5�
���`�{SU-���"z��A���h|~#�-4"aۡ2�P����ƈ�Zk�hb-��ӄ�_]��Iޑ	�ܽ$�8�37/��(�BRFʐ���GL�;�T@��-��)�	Z���b�A*��%�i��T�
N�k�ׅ�D���Ġ��8_Ux�zy�bV`�*xg���g���⟍c��v��y�2#a���`��r��p���ဌ���}�Y��sQev�:^�.&����)��Suљ�~�S+�����5X�����2��#�4�RBk�e8���p���j��[W"���6�TI^A+�Qϭ��Ş�@�%�z��"�n�^S��<4��{�V?F��^�u����"�9�k�h�ys����5�H�9��Y��Y)����R-���B�i �=�r�׵pCh.Cy6@c�\K���ek:�6�2b$����#/ $g��ox(��H�%�� �Fd
%H��0?��v�#��p��p2��l���g'8Ǚ0_���ψI��U��o�����%1BO눀}���2�b�ӌ7UIe�x�����6}z�'?)�m��$N�C�BЀ���a#:(�Me>��v%½c���.Ƀ��hN������}UNð���Z��{�d�MW��r5��Ji CdH$��V��"��D�5�q��@?!���'Z07��'���  ����*O�w�7�q4���W(���7g�R�P��6�$�S���ԭ]\�T�g�.77k��� �TN�Z��/t(��������f	ѵھťG��A`G�����4����������.���q���AMLmݰRY�2���K����'�W����kX�?�`^^i��n>�u/��W�ݤO!O����Z��i��V?�h����`��Ʈ�ˑ�����M�s�x�8}�B7 ���E�')��WQxWJ��ܿf��w6r� 9U�K � ]�U��C����D����hR*��5�8$O�/>z]O���Z�����/Zj�9�s[��%���L�L-0��υ��Cn����2���'=�L��y��/�=���P�y�h��h�8x5c93WSmɻ�U���`����LR�KA���z��K�k�vh�x��v&x������Ц�oy`���)R4}	X�e蝀9�
S�7��INž���`Z��Rty�Z�3���|���n��h���wY�ϯV�J>�a���g�)�0O-�+��ߝ�#*F�]�ۑ�	7��]=٦�N���Cc+3��;�g���x�е�Kyl�I8�G�O�-���V��V�{.����b7����\���s��܄m���%�$>"D��'싾���fP�7�Ab�f1tj��յ�����E�]����7��%�SX� �D�d�x6�	���iK�}���|��=%�|�Ѷ����e�Q��G�-�=�0����<�)�Ņ�%���[F��]�t�~�&gs���,b����p01�Q�ۓ=���v�"(=��ܑ-$�u�f=D�a�7�sGmS��C��9�=��,J|�d�p���dە�M�`N?G����;uE�ֈ�#���9>9�@©�@ư�d6��&pP�v: ��[m�*8��b
'C`cյy�ᓠ9����ڳpk����)�:�y�fV����K���/�*�}��n�#�M�f!$c�\���ÓVX��JZ���.�'<�C�d�-���.���ش��(Z� �Ǆ!,�|زrK!Ñ�װ�W�t�
׼V�����Yme���=䱶��q�P�zg*I�n �<��}��圻�60d� �~�sܞ��.�xM�N
���Ѹti�m�J/&�w�Ռk�4<�VIw�`'~ѷ�{�q��*R��h����$�{ͱ~�h�I�J�������]�����V����e�MW6����Ξ���Q-'Cd�;y�R�.�]��u�a��j� �S~�o�ȑ�3 �܃��-��g��t*��d��
I�ll,�f������5,x
Z<ɖ�_Z#�*�s��f��wP�w��ן�T�!���Z����wE^s��TEu����Ao�o��W��@d����-H�+������iv
)��:���*NR��Њ��IG�	��J/��$��	B���%m�=9��Sn�]��3�#�U�}Zگ����ē?V)RTi":��8�Q�Z���t��/�8@�Y?tX�иT&Ҹ�������&d<_&�^��hm@�b�?�4S3�n��!|��9���@�&߃�"/�g<ma��~���pp��z}���]JK��-SY~��	��q�P:�*��n7�^u���g}������2�x�`��n��G�vPZ�r�����m&@��n�F
ǎ�9��'Z�=S>�!5?w�gaaL{��%�S��*P��{{(��c8z�)P4"!KW#�}��Du����Ū�r�-��k��J��oHx��=�����JU���p��ؑ��-.M��������|�TQ5z}�c(lo���N��&���6����R	�m����׈XsN-�ێ���O8��R�|O��)��(����3^��\<�c�|�G�h��a�)x:jf5���+�u|������~"O��<Uت�S}�e�w���s;1A�}�	%�*Q부7�O	�?�}m���i��y���$�]��pf��E_؂�7>�}���|Z�Ɠ�b�E�����p!9�]W�_[6����4u�!�����Q!�$��a{�g�T��(�uh�����2�5�pqK���h�z�h�x� �x�"7�~g�Y�D�ߒg�?�&�D����-��Eumv��J wև���/�dJ��qǜ��'*�]��K�P�!m��:В�EI�4���F�� �J+����#4��G�S��A�lً�$Ló�j�e�a*+X��$�E�좱���O9��a�O�*�����7Ud���W;�R�ni!�#�lӕD;��Q�F�ítM��0()���wh��xv�;�)f%ߞ߲{�8AK�ot(t����cYL'����n�.O�"ɯf��N�җ�G�&�OUC�T�X/��|g��5]J��H��9������x���(��+�&���E�xn�Q�7e��Id2�������f{����p�ց1�,m k�am�p΁�.�N�CL���B�.�nQRK��@R�������$����z@�N���9[���{��A�u�q �ٽ��v{��`l�ENyU͕�P5�VW{��t�J�)��{2S=��ٶuؿ-�������{G�?�{���#���>���ȶ:�`�Oe�tG���C�_T/g~�#{��N���P��Y(�܎\T"w�td�.�̯�)��bp��C/ ��@���J��b�A��& 64{@֒�P���:��h�������t����4��˟1�C��ɮ�pzEL�������"����*{��j1�`�^j���ۿ]��L9�vvК�����
��Nl�3�C}^Ɤ�)�
a��λ��c�����z��n�#C:�ZVx�'����'N��h�	��H?�qAq��Ҕ�N+�����P�D�p�4s=��T]���F��/}!�%�G���t���I�ں(k����~���`w�8A.Ū�T��]�R��۶�1LP|N�G� \�d�����1�6�Qv�xǇ����=j~��f��Ng��sô��n��Vfq<���5s��W_��F5�a���{�F�CC{�j�}ϝPe��H>�����Ň�`�ͽ��}PP�ƛ��P���a�>?�w޵���ͭ���$g
��}����_��A���2��\9�Y���`�|è�ĸ���q�1�b#\��}���G���ąE�%(Ζ���z��@��F+v���wMoNj����!Gy"cY��ɂ��7��y�ʭ9��i!� FP�̐i_��W'�Iپ�%�|ɓ����Bl�/3����}��&�◠F�/WJn����|�2�ieҋI�����s��҃	�K:Z�+J���Ek���Bp�I�DO0��B�EڲNwc���j*8=x<� ����Ţ�����}�)7J�n��bզ�j�tG���<�C^OW�mI���o��q�s��{�@��	zW��jJ����! �Ho��B���w��;�-ݪ0�,'��y�IY�IE}e��d7�UG�[gǣ�/7��Z�P�:i�c��j-�!�A'?&H'���I����q��Z5��>9-#T���l����Y��{�rv��7JX�2��n���!�
N�L���3xKt>�s�e&�_��T��Dc�H�E�)��-�2yX)�� �S�*Ŕ;
q:8��������d���@S�Iu��Ҫ�u������g�ҋ�֭��#)���GE�X�Rvm�N� Z��D�+�cv����(Q�e��&�c�����j#U�	��������(7���c��o��2 �콕��˥��	��̖���n�f�\�G���4ѵ6����\�1�l��}|�Y&g7�)r��ҍ�V��#`��~K�#w-�R$�&-O�n,X? k]�9_'n{m\��ɏ�0��2����	�@X�H4T=�1.Α,"�r���d��=(9�E8R ħ=~�`Wl={)�B����ݼ��%Ɉm ��ύr���カ�$�Z��U��qD�u_�� ���窖��XW�\��7�Y2b+�0B��˗�!i��w	��{��s�Ak��xQ#����� �YWܨ74/�Ң��_����H0CDU ��v�w�dSL��S��	��EG2L�B����z�11�8��V���������C��v��m�����F���C�w�}��qU�zHτ�{�O��^��R�	�>h�א��9?�,���5s�u�U��118k�nz�?��_,�������E>�hX����BoɌ<��}%�,�P�ǂ��a����u4=�P>���Nv�1���uF(�}�)Ū������3tV�,��Q�
�|�p90��_�����
@0��n�G1�����A(E����攲�T4��J��3� -�� f�0XG�kJ4��*���O?L��t4�,ɖ�ׇ��R77<I��$�,x��[�j����H��K�� 7�VA�'KPS�cٛ(���q�ڂ���IU�W��`׼W-�<w*%�����@�쿨��}�C7tk�G��B�TM;Fq��.aY�,���z���EL'�cmا,Q��`Zc5'�Q�&�ğ:"�^�܏�|gn���v�iG����Cf۔�?������ؗ�+�����Ǎ�.`N�<�y6��������@�Q1�ԷY6��.�m���X#�X�U��Lm�N˟R!������%(T��BRI6�ˆR�}M�\�߆��Z��p,����W�����Ζ̈�a�f�I�R�a��C+��,��k�O���)�U���L���C6��Ώ������ ]_c�����6�}�-:
=;a�u� *��*�_=�<7� ��d��t����	#���Ⱦ�H������a��o�]�;/�b�S��s=\W���ﺥ2� �a+�oEC�Y�=���lp1�A�@W���8.dש�qF7j\�0����Pm�fs�D��_��]2����_hER����C~�3�;[3����}������u׆��MբiU���RGP�-�8���`<��@�Q���b��Bn�SY���cVs���0�c�@4�����k/�#!�z����O=���8�3s�_���+A��0����>��w����@}|���ۼq�r	���oO�i�S>"ym��r����a	C�Qɵ��U�Y���]o�d��W+��0�#�?q��Gj���7��wd؇2��Ώ=w�;���Sl�di��seoy�6I� ���,C`'�1=�h��l�u��h La�!�xeF��ނB)�>Т\�z��`��W+���Æ�%ԘyNA�9��~ �m[�;�����嘮+E�-	*�G�d�S��6�[��|p�Є{~��Qa�Ou���Mu�Ʀʺ>k��^�g��O���P��A(>Ғ#���;M���KR�]a63dh�a"��fp����q�Vy��U[f������L���'��n.����&7�yn���Bu�� ��F({h�S�E��v]�#I��|�}u�O倿b�E�mE:+<�'�X�K�R&*����7,���w=$��=�F�5�c��s{W��ye5��T�h�7v��*$3��E�gDִ�%/Y-+.�oÃ �v�-����u�xb[/���#��Ū#���Q��;��00=&�ꠐ��|Š��F����l�j$��}�j]U��i>rD=k��()R%h���	�x�[�7�ͩ�9�'���a���+��X~�T�D6��	[Ҵ�I!�#$q/ݰ��?��N7!�q�IF��}�!�*�!L�N� qK��y�)����cI��7*��-���:+w����~L�S���:� ~"�HӘl�K�VŌ�&���@���('R.�RIC,��e��눫T
Sa �d���3����(1�j��o���_^}$���rUqh��٦�X���k
Z�A��O�W�-��?E���]��O��W�n���3�&�h'���$2���诟�ʡ��?5����6�_�V�O�6i�TD�`bD�!p|k��LMضe�`";ޚ�#ݫ�����a��۟U(}s@�lo��X��ֱ�'"�y9�.1�Pދ���e��#�ʵW�]�6����<^��/���3��
ԉ̢:�`�|�̘b�-_��a��M�'iuG��/���͙��I:bu3�y�}5jjX>�W�X�Z���\�ʷ�����F�k����灃�C�c���w�/Ac�&_�RFXi��3�_�'-`�g%����v��n�څ�7>L���!�;߼��>�!9�cWꆠ\۫�m解�ێew�*��X���&5PP��+��w�[X$H�Z��v��*/���3�"�	'<�
f���G�gV=O��,o��B�9@_):^�.a#����>�K1�|w�P��nZ�֌�s,�a�+�F8dসDK7S��|ͽ�� t��	"~��>�K�����l�^�<ܖ��;A%k�3�k{����\��0���
�%5�����S�a<N�$ź0%E�#vA�ho�nC"�Ѯ3��pm���M	#F
���j�"#k-�F
�Iv�|���� �1���p��z��نTjY
���F�m$�*t=7t��0�Nj���}x�x~�$��,�BJo۟��lv�3z��V,���V�\��Ԁ*9��X�=��[N��Oo�w�'���	�Q6b,�~P(ǭ�(?��(r;8��R5�϶(h;>jI�A`U�X�׈��Ǒ�Ϸ�=K�|(�O΋����(��OrNh�kd������Y2~��P�ȭ?�Mpt��z��3ޑ~� ��?l3G�9WO������6±�.*%҂AoO�R�� DR��*#͏ꆈ�\^�f@��.�;�����[�%h��%���FD&����_�t��{���c�WYZ\�Fr�N�A��0E}|��;{�w����[�-�}T�| JǳޫۯӨ`1�����չW�e �N*�� ��۝Mn�rQn� \�O��~Z�_��~��Ah��z��Sx�!5/`��|���D�&���j��ۼ~,\��R�7������ ���n4���fŀ�xl
��O�l_)�,�+2Q7�Mi�V�>M�?�%�~��9�f0�r�u���E�bp��E�9Η���{������x5L���j��-71��C���]�~o�&�JݝR�_�A�6��� �?��3CL��&����G��W���Y.�W����N�?3�#A}O�)֙�~�h��r�Lb�3�7�Sf|�,۠�_9�${q^����ύ)����k��b�؊�7�a��sh���G���yӋ�S����8m�%�J��+@)EpP�G���y�x��)�㪌��ޥD��:=u.6�2�ﭧ5�d:r����s�w��V´3Ȏ��v����W*Mw��AH�X�%�H�-�Z5�9�W�\����Ϙ)x|�RPiw#"ҍ
�%M��Aí�q�X�l'cG<����:�z�{ON�*mc&�r��
٦3;����!�8�	�DЛ�ډ���S4ؕ���r���&��l8���+G6�v�{?Nlx�iLߔ���S�Ȗks��c> Ԓiw�dP]nw����8ك�F%#&k�%��ʽ��3A����� ���r4�b�� ����zq�}@2}2�}�%c��� Pw���`��H�P��<$���잘{�l��M��I(e�F;g+@I�z���`�N}WEA	�W-����q��H|uAI9�Bc"�U�b�Ty=(؟ljx��qev�ݚ�E��������e�����v!��ܥ�2Y�.�3k��&K	�����5躣Ap�9�+'�Ғo�Dr�%�$�w�ci����m�gcc�>�Шt� RVy�K|��GF}]�g��=1P�M&ɨ�?��7��ÖgF����0�Ԯ��A9�w�����RM�<Po�%܌��d�n���ؙ/�����(�H�phY�;v����(�\��-Z�"��+��5f�NJ[���E���nzjD[��}����0�ʓh�k��<�-���v��P�f�R���#�i�p�v���[5"���cC�H\cs)j��u�N�H��V�V4b�`�ԧ��4�WI3�G�הA>�M{�K�F\BњZhL�����(V��pd�1��?M��y/�T3��.a}����B 7lX�i����k�d���3T��v��#�ɮ�8��NB���i=}~��7%����U�
n6��F�U����"E����H�\A���XɿdT������ѳsr)���g��/-�� ��{��Oa:�aW�eUt����;������k ���_/�m�⒙�M�vG�B��h��/�َ<�X"`_>1��U/�m��!D�C�X-F5n��BZ�h�k"�ha���Z��y2��[��HhS,Q��p�d�o
�7���V�7��g�$�|���F�v��%r@�!�R|ǁ�K�+�ʆg@|T�*��U�Ώx��8�*|���+��B��u�xb�f�1aI�`��^%�·�!ї��u�zh����Z����5dz�X���[��fڇd{�j�S+�w}�I'�.��+*�N2
�9O�N�h�n�ʖ�20τ��䬟��j��tP��I������˄IEV�;��SON:�S���g�@:d�;�Y��$r+BF�	�3O�?Qą)9}���%�H7dv��{�b)�cR�J`�+&�;�����/�-v�4�K�� ��X�O��D��a��T��V^����+{�S4j��j)!��xqGp��E"��m�m}Br��6�;Z�:w���Y���0��R��:�odî�*`oTa/�}�Ww\�9t�����N}|H'\;{h#��EI-����q�c��UfMlB.�ۯ#O�#�5je�;��ry@37NR Q��D˄�_���ԃ������U��� ��{r:�څ�i�_��ٓ|88`�XiU�4`�Q�l�DR�rlF��N
NDC�(��_m���]����k^:,h⑃Mvǣ��%���$��b `���B�=�'�;���נHXn��e΢��$���L�h'e�k!7B�2�ฯ����2�4�3�\�m����:�iv��3�ST��%��N�W}n��*Ő~8�(�M�� �4�I�K��s��@55��I�������|Zg�¾�J���S�'�o��;�f���{NsU��� 3B�-׍��m�3K�&��h3+���sC���i��&��m����]���򹦛��g�?Yw�;��@��a��_Dz���;���t2E���}5�l���t,v�V�@9����}5o?���"4hۮ#�C?�+!�+پ�53��,)�������a~�7�Q\����OVX��@n�&2�&��6)��wL\2�A�pw�X3J�����%��M�l�HJC���}���_�`EP�B�p<[|\����7�[3���VCJ/�@ 	���I�d�N�o�vV���â���f�a��'�"o
��,�Q��� :衬��>3�@u1�٧�����k�p�I����?13�
���aq~:fo*���*��G�W&��%�c3�P��Wq�A�]���w���0g׉�����N���q2@��-��<PJ��#��c�q��ՙ�gD��ϯ��?���~s<�
�i�[ P�=E"����f���+��<Ȩx�˪8ttOQ}���k衩5�HaUf��zx��o�!PJ\%�;�8��n�͊���7v�NR#�sX_s}y����.�l�֐�UCk������_��i����B�{'�Sh���|Q��yA�U�JI�[[�PP���f�d�	�z�|.(L�w
��}�f�	,�5E@���s�����+�ۺV��J�.�����*��M�y�ǡ�zB!$]�W5*8����>����B�R��c� {�1��<B�K����8�ս�B��>A�S��4��n�DE�3�H�1�b%l�*��������ܚD�N$����ģ�L7��J���(ݾ��I�%�2AN/a�x1��ě{R7\v��#0��Ϩ&�qEr��lǇ
U5�
�$�N�Em�$`wf�{Į�̼�R}V���N�;�D%�p��`��S)�����{�e*��ǁ'}�䃰�i'�H���#w�v�����d:�^9����;�?��6d���u���� ���J����ށ���Z��-7�f������w!�+QY~��P�l�8Hz5�+U5�`n�^�x����n/G�[+��������+s7�5u�V�7��>��R�|&�������7��|��^�E�`��1�n��"q�������!?����3o�_OGddM`�D�S���`�3�z�ꩍ/�;u/�@��L��`Ĝ\,�.]��	P��ҼB~ls�;���v�����G!���I�L+�n��99��M���Z�ɒc�u�8$[:�^�Z8�N,'e}��W��æ�Ql��ϻ8^E;9&!���fk/]`Ծ��S=��b$���ߕчN��q����re�d~�5���C��蟥ݒ����� ��lF���
4Y&�*���E�Ȥ0a�FF0	o��=Rk����G��� �����KO�=�Nh���b5Y���+1��X�����\7l4m��߸Ն��ߧ�ܟHT܎���*9ך��'�u`"�p�CDP+������<$sH�qVG�0��d�h��HA���{sv��9�8��\�w}ֆ�:=���Φ$ñd�U�����q�T��3W�W�F��z�t��j���z�h�qn@� ��Ji���� ���U?���I��@q�(�YNg�s2��pB��T�vo�6'�q/���aSj�OV��~�'Y.ZP�g˕U���~�L�Kߗ�u1ƥ��d�s=t���.���B߃�Y��.�[�j.�����ta(ц�؜��'���K֘�]�M�,>�@칱���x+ځ{���S�����ډ'O�85�N�^ƙ�g�s�ue���������Jpn���2�C��-[<Fq��E�ody��Z�"�Pu��1;�YnTx)"�Z���z> ���4CC�5�=k�h(�ەb�F�$�tc�S��$p�%W���|%4�XO�msPF/i��0�	nX��(ұ׏�ݎ�-HÁ�g!��S����Ӌa]��|".OD�8`�V�I�=�X�S�6k���i-*�)�h��8x�(t�ќ��lkvt��N�,�a���t	�^H7�U7�m��
���XĆ���s��Sd���<C�l��:^I#���k?���h�ݰuB��|B)���z�dEL*1p����t��6[�o�� 1�7I!_�E>��U�,2G�Ƌ�k��	Y��{�R%;�aLe[mq����O�C�y��ne_�	�"ir,D�'�
�yQ@Z܍�� �"u�'P�ӌ����6��ܘ�9�L{rh��쓶�������Pw2��� F�OQ�3��H��|��BsH.\�6�X� ��D�Uv{C%[�Z��S��Z�H���D��j+�[���$p��Ce�ӕ�#�Ñ1?�X��e�f��"��������p��ιsǛ�x+��4٬� >�DAB�z�U�k�M�h,��W�� �S X�`�Z�8jQ�D}#���[�ȋ�p��GЂ���� �y,���!J@����y@�%�A�>m���+Og��m4�:����(Ԡ��[���\aU��8i�a���jB��T�תb�)V�����Q��3�pLN3M�����w,Z�W/���o����,�y$��yfQ�~,Ŧ�>9P�	����`I���V�A��Tt�H�,(��{"��F7㹰��٦���y*�n_�u�M^�g
~���ɕ(F�� ؾG���m@��O{-��<ƍ8�>^��w�z�/o�d���2�s�x�C\�@�a� �eM;��b�e��X|�z�$��WoX���R;-{�)�XR�q$�� QL��n��,
���0tQ�T�iDZ9�r|�:ql�T ���m��f�w k$�ɍ������ ��,�f��3:R2�
�m]��n����y��s�t����%x��f���n�����D�*��~��́�'RU��Ig��` �|�ťo_6砆fS��VB&�r�8r�^�0�F�'�Jq|��K�:w�{�OQ;�r�+�pt�O�J��z�xs�������^b�T��~I�@`�f��O��M&W9g��b&-dG�/Rd�Vڝ"���R)QTD��p[P_�)�a��H� �E%.H�c��ԯ��Zu��#���Z.*4e��8�-1��I}�86zm��K�b�����vq�>�����/ujf:4>"�t�0��:�;Z+�7���#��\���H��}��R��/��Sͱ?$�y���!lc�p;Msl�Hv�C����u�J;t=��V\�8Њ�^��e-]����S�m m���ӎ6,t?ْ�brٌ��2kΎ�����A91�"��H�V_	/�K�!��!4U"�h$62H����w���|É�h ��ͼ����PA��ႏ DQ���`��Sm0�Jbg��-����3VPs����W��
��^qV%��~��S�-��H����WV�,�p�[�i������X���������}��n2X�)��d��nUp�~�sL�i��P��
��>z�]	0��p'��S�A�%�(� `�$l�UkK�m2�t��(�tDg�l��v�'�8���m�'�՗�)��#�#M��~���x�)67�-�QJ�P��nz���/0L[���۰���"��|����Mj���X��X�͑	a`.舼L��Xr�s|� �Ը�Y�o;��5L��'�;�3�Ѫb���Kyvt�p|i-��0h��p;s~���N��T��m�������}+:�;��>`�
m�8'~��6�գ��\��̥ѢJCz ���垦�w��iH��4h�����4�bY��r���h�u��2 ����3N�_��C���f�!R荭���υ��֙��a@�M��q\����+�7�Hr�tl�]Gj"�����̝�@G�ȗ� #�u�nw�aw�fV|3S�mY>6��i;�k��ʬ*�T���)����c�t�[��&0naI%5�=�>6���B�{Iz�_�y���B�]��5��a�ftpGyP=���:���@���?�'�3�i���]\P�0�p�gwJUu�������[�9Yx��$�(�@_���_+u�����ι��j��,)�d���"���\�|Y�%�4��v�<=����=_������*��������[���-��4x�Ώ�L_h4�	^�����7�g������߄��a%37����PW൪�ց�Ub�y�#����U�$y"�F���]�\>�\�_�L9�OA�W�kA0��~'�e��2���Ik�<��q]3��J��nH�.{��+*�Y�����Z�Iq�����|�*��&2�~t�m
�sr�$�����	U�GQ�� @21�l4�0Y��v�e��k�� E�~���������Q����X�Q��`�p�"#Op�<о�Y6@D�a t����N�7c����i#6�2�'g&@�b���F���K~*�� L�M���3Ý;�����J�1�����/�B�O�)A�`�]ڎ�%�a�8�[e(�:T[��Fr����(�V=���ʉ��ڹ��Κ�	�;��lr��O�5��58�=�%��;��l�+U�y��ifڡ�9<x2DlLN�0�d	n��)��5����Y�-BK���n3�,; ��o�@UU�"���v���'�g��R3��	���4��}`Ц#��Tg�wF�`3D�"$=��ϛ�&{ti��k�=pO�~�=ݯ9�1�_Ո�`�����x���T%�n#�|LQQ:����w�0�N/n?t�_�4�%�e|���y��;�W�6�G���
&�8�J���P��{�JF&���3���C��c�D��3i��OV�7F�L+oG�S.���4�\x�@0�E����@�`I����R�a�C����,�ƅ04j���ڐY�����y�6*���.e�D�4n̨�S]��U�G��P`Z����L�TG�y��ɂ�DhO$@�^��Ū�Ŏ,�e Ѥyg���}s�?qkL�Q�w5FM�RU�]P�|
e�ɉ�
�T���t^rWT��J��q�/ŕ횜绬�\��f`��{�}�5�7D�lp�X���c��#����,L&�������*Ժ�}W�gN^�.	7�5���	�R��o[FK��%9�7�hfD��n�/t���Q_�C��L6s�0�F.q(���y��/���_('k~�a����C(U+37���cM��jx��ô��tMbsQjE[���^���r�����K{:�A��楢��3��D�탾�Vr�a�D�刔��;��vcp;��B./몷���M�'��)��_��v����@��}ʧZ�LU1�#-[�-��ť8P�(.F]s���E�r����6�2���}{����P�7�MG��qqr(3�����8�}GZ��2�Vg"־
�/@�n�R���^G�dJ�Ց*`��~��Tg��U0o<9s/�$R.����6s�g�H�O�R��Z_�Ƴ*G��%A�Z�UPa��A��Db����)b����&�[�������n
ʈB�x�W)�kԥ�b���_���R�����@z�.p'c3��;�7 `�@a?���5ع���6�j_;!��oc%�~ ��*O��5/���<~���y��&���^f���w�H���	����M}ʁ����N��~#^���sn�w�^�ދ�����.j���ނ�M���G������������PD6�'�y~nV�̫��jP�r{�5����=���6���'A�zy�$��+�ɁJ���ͅu�#�ޥ���hj�<=ޜ}��	ջȊ��du��j��� �YǪ��g%k��p�a���YP�_�Y�U�x7�Xꌏb-t�~����J�f#�\v��h�磑hh�}HAj����(%m��9�����S�Id��*��]���[:pj��������{��ڐ&7���>��J��֔U10!�.�B�o�~?1�����B{��}��c�����'J$t��l��G��v�**�Q��B��7���Q�r������q1'�e+��i�-*�>��kȨ&ڌev觑 ���/nga9hv�`��z!t �c�mQ=#��K࿜䠞��f�h��B�%u��>t��Ǵ���e-x�z�S��x��5��KgRwGϵPyqX*rl˝����G`�
����KVidk�]C�'���T�\�%=ڷ)8z�Œ�сb�"U�DW�f�0dJT?b���$s�q�bw�B�ↆ�>����R��U��)=���F>��>u�u'��ܿ�H���;����|����]c��U	�UypA���Z]�x5���Ic�x.�-Zp��<��q�Xm�d�:"��/6��O���qY�kZ}ٺo�Jv/��+-t��$�d���@5���\�l�$�Tx!�����i	2�������vn�7=8�/>���pS�s�u�U�F�<}h����f�y;���a���[Y���>�=|���ŋPB+�ORc�w�?;sl��b���E��e�o＞�~"�1?�츟�69��B���,z��,R�����la�j�Xk\��AZ��N �R�[��[�W��������"�>��d���3��Q�Xte���(�M�!|e`�t)�̿�̝��JNS�*!d5#�2{�����C'��/��m#�̯QL,�:�0����wG�=ݴZWaWc���aP�]�s�B���cT��!���X�F�)/R,�"�m�Ω���8��l{֩]�Q=գ���G�qa��M��)�=w�m�oM)�����*�;�����k���cI[�xs0p J6-+.kf%��^/�����\�$��8-��kdQ_V:������[���/���h���!=�\P�� �_���J��������u�"?]�����m��R!SN�V�5n�X�2�}qKo�����t� _x�H+�~D��u�.4Gqk���=F�:l���1��HIl�9 :�(K[��/i�钟��#&g�_�:��&�(5�����F� y�'C�r�V/�wp��IAku��^7�IGT^� �Y���Ea��iAlsv�%,;y0���;}v�>vN�|G��� Kk�����3�zr����"+P#�WU=��� �(��:���֘��||�������(>�P2-�-����J��ZpŐ�qS� �q�?��ws}�R����d݊#%�Q�\)b�1��`v�̴�Pm���VH��nD)@��u�f��<� v<�	�B���"h��
��/ /2�٢~�ސ7�s��^$��HJ��0'Sp9#���������iA�8��E\����5���?���]�<Wx��H��E�(�-BF#J|Q��	v�=x����q^	}
�.�����q����a��qE3+�⑤d~.p��d��/2&/�8��� �[�� x���EG.a�@��iv`��c6�	������a>ta]QQd�԰�!XҞEE�R_����/Wz�&C�%��ޢJ쒋[��O�7��m��؏ݢ��8���ym�@�n���*@�ȤĴ��Č����.���.��7��E��W^㕠gLBEf�V4��1�����f����Y��B��!z�� R�$O��ћ�a�g��w�d�j[mE�4~+7���#�,1��2��u����{��#SoD7�Ct��_h��ՙ�
�Ә��ҝ�������{���#z�0=F_�����v�,J�\�*�oÈ��vy�3��N'����Iy'6�&Κ�Y_42��
��8�nW��(�=�N�k?��k��2�RZ����Ӑ��'o�v,�[^Ν�"���l*�ƥ{�Ԩn{���hr<�/ݩ��
yg�p��n��l2~�g�[����mzGo�h��ᴘ�?J�!(�:��#�1��\���g��!�n�����u�9e�I#�.�G�r�	��3C/��J��������IQ�<[p�pY���a��%�)ۉ�<h�ᅐ|��(�����(�ݗkfs�9^r�%�e|�e�ڧ!B?�_[�}����>EKK祍��}vqi	�vځ^Hu���/G̃'(�Ş���f�$�x�H�LM��fe�/�:q)(Ϯ��6,j��{���4w�Xڤ!)�-KP�K�"�f~�}Yĳ���� �\ ���t��"@DT=�V��~��M�G'Ƒ��F�f�k5���*���}�5f�$J\|>�җ���6ekV�C��O���Nxe���q��E��<��ՎSQ�髄�g�����^�Nȿ�P�sB�Fι�Q�wL�g�p4g���z���~�C#�O�"��e�[������8�_k0�I#xқ(X@%�Gӄ;nn�����@�Dӊ�a�H��
�=��DV)��]�@MBw��>ڷ�)�����՝M!��Ć�|���MBA-�������ۭJf���ueF��'H��h�R|���p-z&'kNʛ���">�����!d)����ڳ�����ܤ��C���y�A�(�V�R��+��C��	V�Ϯ�T�N��a8��l�F�� $�'=Ue��eeR\B���r% 0٥�h@��X�����ٴ9�3n^���G"�3Ls�,��tiQ��2[��hUAV?ߒoX�>��vtd�I��>璍O�� Nj��0=nx����J;�&Z��-h�\m���8^_8�C-�R�LnD�Q`H<�;��a|g�R�2�@�n�1�����S!?J���`��Q�̋���xTAc~XIH8�����r8�'�Ų-�ƶ,	st�Lp��ż��ʢv��
�
ʖ�]NY��m�P�+�ϐg���%'N'@2�R�3�b:���=:�#��+�U����{ا��nVgN2�R�D���ǥ\�����7��Nl5 ɑU� �s����{�N8�0��!��Y��_��n,O<k�����TE��G�	��b�:7�2�'z=�gϧpB��y�oy�C����@lV���؂Nx�'���Ŕ�o3�ZxX�$�{�z����;~�AQ �%/=(�>4���o�G+��T :�ipۼ͕^
����5]��NFqK���84��5��D�%(��O���Q��3hC20�s5^#uS�1��L'DH�+��E��|w.Te��Yi.5� �IlBj-�nU�^RS#㰌�b�t�Z%�R�5y��l���i;}���У�)~�� s�/b�yg�Y�#c�`F-~�&�������ęK��K��t�͟/"P�Ⅽ�C4��G���Ch�9��k7�w�;*�C-?��F`al���'�1��Ѹbl��(sd:S1����q����.���3y�]rp�;�w⛽5��Kƹ��Muc��axp2��T���=�o��#���uRȁ���O`�f��s�b�M�L�I��k��e3 �)1�� �\Q�2Ѵ?�¥�U|H����/o��k��<��N�
)�ʃ<P�)F�&��.���(�BQc�ZT�G(��wTv��Hr��q�a�\4��A���X���)�,Jz�B\���q
�	�0_f�_�������/!���
Pϙ�c����r[8v�ib�a
�����|�#HL\{�P5�������P�9۴m�8a'���M�7����/)ft�-9J��r�߸Ƿ��+!{�r�I#�lʦ���f��]�~ŌW흅[�A��6ʿ�j��@�� �dn�hrz�=�b�.	�B��niS��C���R��w?�"��"����ఄ��)��"��	��"��	��b�nE���fB��@w���w(��C���uP�ٗ�����&,�ŗMZf����])�w�+{��S�t�v~���}(�9�;=3�8������G��~��`����_��t������i9,�F�;�� Td�w}�Ń h���[�˱�܏'"����/�a��*���.Kڍ���
�%�ѧ�\=�����E�u7���,/qwt�s�Ј�k��؍�� GT<<���#�<�lf<M�{�ߠZ6��.�D��2J�߃�tQ�=�Y���~��T�^dv-L���"һ�}��l� Y����S2���:Xb�F���-�F���)�s�Q�옆�?>lb��u �{���i������P>ӡkYF�K8�茛�"xY�kY��ӡ_��	I�4�fXyV�{t���^M_��&]�������xH��&����='3+�%�\�͓��S�"�A���m��/Y%����'��4.����Bg3ܳK׸[��s}���+[�����r���?ܤ?t�;��Vc����^<��"�!t޶>��]��#s��M�u���Sa̾�T���;ֽH����2�(~Z��z�2�ࣼ�� 0�y�i˶�CJK,�+�����ݢ��T:���T�jB$,�J�L�.��K{}(z�ּ�PU&��Ґ=fcP���'���(���fh��C.Y�6����c�HJ��1�y[zvf5Je��ɱ[�m��;`4�m4�|f���HIn ����ڷ?'�(1��S�)^a�d9.h�0x#�� �!b�{�Dm�b���.����n��+��u3o�r;a�����V�C��O�J��㗂�lGk��d1<����.��j;+�ŵF`FT�� ��*�1�u�n{���t'@�/�����M�m�|��j.�|���P���K�U�^	�*�>�c�@G:���Q�$~^��-����8mC��l5�AB)����ѫ���̟���^h�"q�G�h��.9p����1cI�}Ɇ��1?2�=�O$us�&�pm���N�zH�2n�z��"��O�Y������a9���r���v��/FD��9Eub�Ŕ8�Q���z{���C�g����bB��V�!W���$�}�%���H0B�cD��_����gI��2�l��*d���yc��FB��O��Uf@Gj��w�H�\�#�uw��ǔ�{ '�2��U\Fѓs�88�!� d��.�7H	6���P�p��R�7N�jQs�~���]��X�!���Et3Ê���n�pf�
����_Ύ��܂��+%F�"��!�l�x[�D:���q�&�|����lj���K�E*�L�����귲��"o��2�nA����c��o·MBq�˧2<F�0^o��ʃm����� �1#+����$}�S�[xٿ*�cY����� �Wu��Lpc�K(��7���]}gtʓ��6��/j��F5�'��O���(^w!�CKX1�-�喰�w.'����桼����]E�>)���L�S�G�O[�����X?���X�6�CXx��32�L��T��M<�U��s�Y�i������Z��9��c�oR���4(�TB��2U�pl��@��#,�ڂ�Oa�j�\��& ����� �=)�%�a�EHS��D�i�k0S�Ҳ�WB�������'{g�݉g�~\Ѝ*�"�W�r�wZ��2:�(�ɿ�@��y՞=��O ������8�������eR����8U��2./������O�G�,%�c�Nf7 ,�<
�T�fSGn�L�(U= �b�;m7�¦}���h�����p6��,��i�����M����/hv��~�� ~���������<�/?�5���9+�ԓ_�=�8��.����}i�ez+������Ҹ�m��J�-��w�����$��M`ܡ	\�ߨv��9#���T��uj��*O�|΀�-$�U���%!r�h���$�e���=�3%Z"�7è� ԑ�--;����dӋ⸦��<3�t`(��s'�ņ�,�+��Ħ(�'Wl�"���/���d�[:��^EHYK�v#��`>tl���^�:V�"cf�{͌�_/�}3ӑ
P�z<�`ň�Ѥ ���*R=�[e���d���	�T� ��ԡk���a�{��	׹����$��|��%�%Ǆ��ژ��1`Q�n��L�~z��y�k�hp�W���,��b�l�3/�fS,j��[����h�W��#]<�`賘�ߢ`l�[��u�k�ސ�D��"�ҙ�Km��S6n����08uB�;ŠwcO����4ƕ�*���ܟkN���clE���c�U��5�r~��jq�puŉ�p��n1�j�%�1�׫�<�q�>�d��x��#�WN+Tg����I�	��s9M��8&!d�z��8�˪/��{p�G邨�?"g����}�힣�`�9�V*�.Wv�ܭ)�W���ݠg7�@l;�� ���c C��fX�	_����!��0]aS�4�,$z���T>� ܿ�!8��p�����QMZaGK��qwW:�`J����fj'P�߉��F'���%��A�(�_����/�g!zq!n�%s����z�f�=�X����[(l�)��q�����ثyx�'�����@�J�g-��x0��#����G.�&TBp����ɼW�B������qT�^{�zb�s�1�\�u�Q=w�d&��Z��c��!���h�ޭ��G4؆��^�jS:��g`��A�j���:�N�����eQĥ�
����&�[��ٶJ��gMA5��ytSTwr���ύIYf�����u�J��n�u�2>�h?O�'�p���3}�Cb'�M��k剖��k���\i����jJ���#�NnQ�-Q�c����f���7���}�rez���ʭ^O��+ �}��B���Q���L�jo�E�שro��A��)�m�H�9 �A!�;��yo����,��~%t�����J*��9q��Hs\�zB�?�g��Fg�3>��d�) ��o�+H�tU���r�7�����0.�Nƿ�{p!8�_��G� "�r1!�t��")�J�o�϶L9�i�4��A�9�q~߷�Fe�!4Y������\��^tct.#�6��v��ηC�>�ܲ����<�[���Ň���5|���� |_}���V����Te�x#O���e��}�X|@�' ��H�{�	��7�9F��č&-DIy��}-�ų�,I��\�;������'*#��&��?����_������_m��4������䲱a;���pnV!�A��5�-Ƃ5�&R�.�<�&n���#�dK6��js3@n�� Y�"೏w�±/\kS�T�E�L�;��P eĝ ݓ�yy�R�
X��)Ǔ��t!���7�P	�eh�D�
�����:{4�/ij6cr�B��Ȣ��2D8pYx�撳^e��s��C'|2_�{��&��񨁔�A��|��b�K�rq� ث�r(/��O��8�}�olD��o)�� �jH�A��M�*��X�n��l���=�y4"��#��A����-ɻD����i�1-)P�b��r��\�\֦��5���4V��n.{޶��1/�<k
۪���O�"=w1�|,��Z��G!�� 9u3��QniN���p>*�9c�{�2�������"�df��é\}`����%��X�t2��3&t�^��z$�	}�� HH��s��X.��b.8�n�N���ߏ�W���@*�=���|p*$6�b�򉷤k�ҋut �B[ۧqհ��W���8�i���qLA�W��,ھx��5@j������P��*}���@|��>��J.�R.9��t����S��d����N�t�LOLy�a�ډ�fȿ��ws����A��l*_oF^�r�����g�x.�߬�wj�L�E���w<��K��?k��]��F�Xp��ekQU=��m�"/�4ˏ�8�x+&ݭc�{�IZĺ��>�:q���OX��cT^Fƪ�/(�F�����c�K���3:���mӻO�H=�e��B>�+�Ah~f#�!`�h���8Z;��k�� �5����#_�ɏ%����D,����w
.�F U���T��l=l�gО��~�H�E*qVN��p�֑�GB�u�Ha�۔�>�>&bgh��fo��h�T����t���Y��*[�F}�M����s��>�M�����:��Ln�~.Q3=g��Z���]M��y��V㐪^�:�2S��9&�����4k���+a)\I�d�=�	߄�𵨤)ݗ��p�p{����Զ�������ޣB;
m3�=���~K�W�����rl�s�����pEA�#����#���Sy� �5��)rlR�4�\�)� � 'M{�(�T��@�(���F���CE�ta���S�2�y1�_&�!��x^x��Ue��w&�n7�g��q�ii��1�>ot�h����e	q���*�9����hl����?C�A��4�M�D�*/^��A��0�L[��4�D�=l���YZ`RT���^?ށ ._.�v:6��q愜#cظ��[�Q�K���m�ˌTݘހ�Ɏ�L�>a�^E;�7�/�35��4��L��d�������k�����'�i.?=�/�-̎���JT�ګ ��[O�]w���S���l+Gմ[��k|Å��ߺnͮ9Ĩ���F?ݳ�*�]x'q��F���I��RH`^���!�0��T	%���mo�de�s�������N�
x�槞[BSʋnY�����;����<}mF!9q�}>���x�1�Ϻ���[�=4Q²_Kꑀ��_W�@z/��O �������<�HTx�卝��:6 &��.��PSᕗcw�0'�B��p��%��J����} r�b�i_qm�ceYg���&�]P���x�"����#_+�����?�	7�T*�B�W�`����ɶ
�u��j�����D���Oˢѝ����2�#��Ȼ��L�l!�`�����u۹�|Gtz&���5��_*t5��}�e8�}2�p�x�p\����%A��8b}=-ᘞ+E��ج.1�:�{h'*���;I6��Y������ �
L>�k��7`	��U���~pj��x���z����_H??eA|�j7�]0@Ż�k��T:�*���6"!��@@�
Η���me�.ݣi��5�u�& ��ܪ��{�Fm��u-�'�� ۇ�6��6�׳Zm �i��߽�����VQ	ӝ��ȉ3�����V�R�j3�˯�艙�3SQ~�#�5�"�jA�G=�P�f�yj�AƋ�Y#�a�;����tH<5�z%��d�+ {9��x(�_�h�*ʤ�0!�8��`�-#=�����5��� X�CŴtı�0}�%��s0W*��D<��x^ИD�zi����M_u���'��a4��4�%�]�LU���YA���r1\��P�cXL��e��J%��Ρ�=��֢[-8I´�ژjJ��{U�R2�W����Ӻ>�R]܅��'�aE2���.Ox���*_�1�?�����,�ɢ���C����*�Қ��LC~L��O�n22l�.^G[��F�!~2�x`��{�2�U��R�z��57�6���U���Vc H��!���Ğt�W����z�܎��g�jc ����ˬ��-�Tru�DPS���c��0�����Q�	/sq%�Ѳp�6��S���=�Z6<�� % a���	w��;4vX����vi �-_��|���]4���Y?�A'ا#aS�d�o�u7}+�+���Q�FJ�l��J�p��I����[���o�bM�/�a>�3N�s	�X���J6/37�,
����Dj��wg��V>l�:��1u6Tnk�8��A�>�������$L�9,��l��VS�(J��5�K��=�4&���P:gL�|�4��M��x��ԙsՐJ8=�����z�K�u@��>w�iˬ���!)r�D��*c,U�sQ;qq�j`*���I�S8�JE�8( M�(�mw� h��Ɯ��C���ؖ����=v��L��ݍ�e�`��=�KD'��t���(p�������Fɀ����Y�=�����6.�P��!�뱸Z�ޝ�>CO#�,�I����I���^d�ίz���?.�����
	�'�/�N��*��o}��+9��B(B���Ϳ����،9��[V��f�&P�<+GH��\b[9ݦZ�e|���*D�6�ǾO�ifqv�ǑQ�BG��U�F���fq�GK�;�h���,� ��4~��Ỳ2�LU�qGQC��6q��2���=rJ�^�{}p����1S�p}�b����o����:��@)�aw��U��љ��W��!8t���{�g�<c6�!�lDY�m�����_\yk�2f��ÿ[!��u�O�%� �[�F�����u=\Ɉ��ےՑ�]xvv�s�\CR��˳�l�{�t�"�d=�kAYUUIv�AI�q�i���t`f�g�&7����	��Tc���C��\��5�����2���K2�8�P�����	�)��������j�#1Ql@k������&��WB�p�Ϳ�~�YF�6Kg�Ir��؄���Ǩ�V�'����nK~)꧃m�1�'����u"�5⒛,�9:�JU���%ت7�H�/�߫�r{Bxr�V��D/��#Ɨ�w��%}p���*{j�&�d�Yk~?.��n�zEQ��9�"�dǃ�}���TM ��=(�c(�lN'4�� ��N���GxE��qoMPYȸ�'�2n��j�r�BꮛM�������Y��x��ܪ�Z�2�L@���+.2Z2-_;���I����b6�5J��&ڬ(V�c��U��:?w�L�:��z��=��֡xW����tX�M}s�-��L�`��Ƈd�k �uُ���2\�E
�DG���[t�O�'��|x�3�`M��i��{��3i�@�;�o�}h�>��_6�mm&\����0�UHKЃ�$-�s�P����#v�N'=��-�C�C���%e��>��1�[!��Ĺn��<:=On9[�K��%��C����`�%n�c�.�<6i-)1T������L��(��Mk��h��./ȼ�݇2���V-o���� �R��>A��h3�j,H���A��G�'����e)�*������ݝ����`�=��
P_��R619LQ��*��W�����F������L;�i346��Ʀv�<��`�2�NV���P{w�Uk�o�b��Xx�� >9[�W�PQit�ޜvs.�oIQ�cۉR�~�a�re3d�;t��2<��k5�j8AYN����p��_����M2����2�;�����)��!V�3��9��7j8��F�u�^pIƂ�4��k��o���N���	�y$��XA�-E�1i����{$A-����PC��:�����z�'�Ꞇ14p�����ӾZ.OX�[����Pv��7�#5��l@�t��n����7������z�� XZ���O���(�I��኿(�5�T��j/�<�6_���n�愤���ѥa*�V���i����!�X=��;&�d)b_�� �]��mn^����Bߦr����8�Hx��[p���@II�2d�p��5��t����4v%�фp�s���.��ժ��'��&a�]c��k��f�}�����f�U��X�b��{�+���4�ρ��('M���ОUf��n6Q�fU����G�4R�̊41�f�s4�a�lE��Mh^��T�Oշ<��#��cf��KrL��'��a��!6�z���Uh< �w1�<�#���~8�8�z��3(����{Fu�i,=��z]ᛋns���)�Ҫ�)x�O�GdQW�����5����ų�D� =�)����ҳ��s�����3j�E8|��-�	�V�O�Q�KҬC8��eK]���I��ί@�i?��f�p+	�� ���� �uѿ���֜���<��S:�}αU�>�tKBt;
]W����*�"����Q4���DojG
6	#���k�:��l.;��fms˺�%�p���'� �ǧ@�T�[x�;�[# gU@��FOI�U�"��L>���;9D*.��P��:��#,����]��?��1NOy��8Qy�]�Gs�S���@ی�֙�Y����|m.���	�@0���ґj--b�\��"�^���j�޶c�C~���%sqxpT���[;u��Q"*`�'�i���N��Z�^|g�+W0��@�u�)�v��kk|f=貯~��[
ǉOQh�=�P��9���d��D�誊�=x�l�C.��h>oQ��w��l�n�E�����R( #d��R��5�Yq�Z�㶘c��S�\���{�9�ťy8�^��9ʂH�J����+?ܡ\�XWU��\��Uq#���ggd
{q�T�_���&�l,p�
�yG�mvW!#UK���ۥ��(ɉg�U�[�,@�{����OL�|�e7/�����:6��y�f�N��5��A~-�w<�4X䭲pK;3�eH������iߕ��c����.�����W����)Q�����Q�}������Y�o��s���q��eFP���,�Ӣ��w\w�&�s.?����K$;��� �W�����c5�䋩~_����فU��8m�����B�7�P��� G��k!�'�������#����;u�XT`�T�����U~�+Fw������N��3�h/14��}����;|�(�q�������k���aޏx�	��K��L��*,U��3z�Bviȁ��'�ͬ���e �|֗�H)k�0�:׀c��A����C.�c���*=����������C�P�xeu2�K�-f�9�y��paT��^�H�U��d�ha����Q�ѯ5��ʷ�-�L��h,�m0Kz�b�y4�ߕOs�:�-���п?+5z}��kLa��џ�M��l�Q�2����P�ˎ�Ϻ�;��U�	�飯�T_m���e5e��{M�����Ȍe��	N��A�T/�t	�H��%�t��Ly���"o�����j�+�p�����n`��ꕏ�\j37�6��~w��vk���L� m��8��D)�`�Z�������ډ�P���W�p�M��Za������mO��=J�f@�{x����G�h��P4�W�0�W����f��hrɅ���a�q͆/��pm��Y[r���<�{�}AB������[)��[�� ��Ƒd�z&*��k�˧�hY@~M��γ�؎�_�y�8��B*��M'ul�W� 1ߛ�pa�4�Y'��;.��+h2k:��|-#��8�N�otk;��G�H��x!p_�� <V�݋�_��_\�u�e�Rh4]�!bw�ފ7�����.ޛ3!���y�O�-���-����BBC�h�(���
t�3-�l5����Am
�>�ൢ��S�\�Wem]��٫D����jk��]?�W^1(��ᰡ�����S
kѫuA-(	i�;ϡ��%Pm^տ�nFz�އYщ�=z!��������K^Q����H��7ƣ0O�0)������&�]���+?��ڿ�3�����Wu�	��00!�i�u����m:���*!~���Y;%ȅ���ۏQ��L��\���XA��|g��	�����90�t�Ә�R�M��*���ct#�	�F*��a�m�A~���/��
�>|��ِ��������;_����+[�	�5�<ܚfqH�њ���Vd�?����@8!�;�4	/%�[���r���ͱB�u�#�]���'�����x隤c��N�¶�/UV�N:��4kf�o%������c\�T>�v�v��g�ۃ�Py���J�Pџ�P9�
NdF�d_�>d+v�6�\�������
\�F�o�;@{��,Q5����'�|-V�9�U&'2_ݼ?x�o�ȱ���]�8���W��n�9�S��p�>Cs�G{ğ�����A2ԩkQ�Skv?�'�VBz��~>�G7����ڔ�8�(w]�n�$%S.�Ѹ�W.�+��Ke�������'��	�V�/8
t	q���\��Y ����
4�䪵K���6P�]k�}�_�&m�چ���G�� ����xg��.r�-��P���tT ����
}e��AN�qN� �%�ִ)e��+ �Mw��!�4�	Φ��i'�[n9�;'0?Ȧx��F����}�#
��{�4��|���ix��綤
��d�X�M!)5��G��-�zw�aU-�!Vl+��˓�Ť͔�*T������<pq�I>#����f�u��%��Xߐ�����pΧƘAo]?��B�&�X�N�A
�c�=���
j;�)ʜ�����u��C����N�$	uخ����Hc��XE�ۏ]���qHsf�p5��=�&xTY4E����ג���"����̪��������!�Ix9�U���)��A�yu�H��{���Slmꀼ{�X}�|�IySvT�;�)��X"o��#q��s!��rP�F{��QB��ȭ��Qՠg��� �))�D/�y�
��^(Aq�����݂uH��X��X�ad�����:깗� ��r^o��R�/>w�ֹY�������d*I �������˞��3��]�7]�K��( ��w��JT�RQ����jf���1Ɲ�GDzR�^V0 ��6��K��L�:rP��U�E^E�p��Zz���*@*�M{Cj��>�B��;�>L�P{͘�}�KxB'��7=�vp�����,0��"�];?�Q�[�Ϛ�g�7X��p���Y`oJ��:���;�ͬ��3d���{��@]rs�@)�4�v��[�,=��_�]�R���n+% .'?[�i�Es����a��9�#�v�)��[���H$al�y�ԟ�~SE4����}!l&a��c�v���B�&^'��5���p��&LgIa`�sm��wz����c��
i!|���0�e�Y�Dú����8s0�s�4���$�Z��J���j��S`ʪz��t͉j ����m)c���Ҏ�b��s76+5��|�K�34{[k�������s��N]t(夨�N�8𙚛�}ujAHQ	�'��]C9@��p��TA��a���3H����K��[��|9��+�������L�&�cf�1cM���* �ݡwwl��������R�x���g�
P�&N�B�����w+�DR���~�oxx����tU��f�P�hS������a�	�J����a�m'p�)�'���S�Ħ�Q  ��;d��.�a(�ӂÔ!�Q���Ŭ���T�����p�v�C������\U���ί������-�Ғ����G���? :"�&)t]��'J�d�;i��&��������N��35������1�� 5?�����WL1�	K*t��ՖyH[���z��}Wݼ����.Vg�a�Kcd~�t8��
�
���J��ƪ�>���J�y+%�|���5r�ӺGݐ(7���Z&����V��S�<9�}qک������+��SOq�y2?C�-��Ry�e3h,�9?�{̘��%"�d�Rmz�X��x,8s1��0�����"jSt��"D��
5�!�.
4=ڿ��I�c�E�w�6�q3I5E'�!Pff�2��"�N�*����E)�Ǳ�qҪ���I.�<��k�L�kZ�~qfr�x��l˅�yD�U�^�z��#BJ��pXL�����Mq����	
��;���A3��#��iUsRsl�O���I���*�e'�u����ne�����M9���4����n��Ր�nnvt�	$\s�ˁ���M�t:D���� ��W4
�`�wP��vp�&�o(U"峗�޼'�]-}�$-��m+�J�z��2�����6,�3�=l2C��=$O�z7�	��2L�?�1� TBKf��k*�o��\AT1�hFݲ���8�O��Zx�z�u��#���N����꺌}�o�3��ص����ᔠ)�um���:�3̀��[#��L�;;�yΧ���p��E<�ֺ#��	.�W^�WxUe��qǰY�F��^9:��I9��P���f����`a��eD(=/Wu��11�i���my`���O�/Y3�}I�Y͗~� �����7~�i�`.�ޑYʄ(��Of�M�*X�UA8ܹ����=���`� �0]�����Ӊ�j�0�S�b�uA�q�:%�uGclk��jG�T������������Cu5�'�B{��еǐ�I)�\���^ݵS�)@op���\����|�'�Jvٚ���A���}ɩ.�{�s(73	�f��|h�d[)5��~���%�y�M�����~��\��G�y��5.��;_L��� Ҫ���TpZ���b�%:Ep��c
�(J��лL���10=�
�赽NUk�^Ю�/���Qy��:�BХ�I; �1���IY�R��9V�t�/��v��(��T����I�f��OBI��R��C� ,��c!��!$��0^�D�MD{�Ŵ��Z��	��o_�^^�#
�f�a#��j�H�k�Mm��Y��S�h��ųz�P=葿}�o����d��Pћ�Bn�Y�������Y�8�E��W����S�־U��T�|6HE&�����Y��ɧz�e�e���<�O��׬SҸ�McR*��!�n�n.��;(k�����be����9p1R���o�	�f�����n�q��).���~�L��� �)��d���Ṭ}�+�׶��w��"C�;0��~��	��K�{7��v1���L�1���P��D3>�4j�㪙^� �q,�lS�hgQ�T�v/��%��L)����`J�6y���x���-ac��!5{�AE$F{��a����ù�R	�������[�#)����?.��;&1Tq��qUW�?Ƃ�/z��[LA�`�Î#�0��2�^:� ��L��8��2俞�'�������~�0���/��1r�g�1�܌-��� }���0�]���R�R�J�� LD(a,Gzx����<� Yw4�+*IA4W�G��c���{�����k�����^D�%����U���&�#ojK�]�tɄ�61>�}��N-ȸ�7� �
���@���CY�Nw!���ƅ��� Z�ٗ�8>��U��m��i�R=��`I�Q�}�7�]C$\����sq������g�Dr��P��du{���t�;+A�����y&��4�.���&�Fk*��B�rSe����n���R;h�ḳ�EkXd����D�>O_��[{���A�
���_���Ѽ!B����Z��Y7ַP���|~.��0(�e%�q���Ļvu����T ����ņ��[b�����%��$��Meo6f�b@��fR��ɬ�����Bz�9]����7�O�b�ˉ�_I�_���d�E��W����(�^���YlOL)���80�i��R)~氳�I�BR.�Y?pjߠ���(,��	��nW턥�EE~Iw��d��d��p����'�e�/ZR�Ȝ����'��D�	�w�[2�R���,�.w �[����}m��e@S���c;��>Qv4|7� D�O��¯y3W^�Y]�e��b�E@�o�Kd"yxc��o_!��	6��Y1��A�P|��)����o ���#ܧ�0�4����zaw��ڢ�k�����D�yKr����'4�0����)j�]Y!��ǘPnp���o9�M�X���\.p�ȼ�Q���	kd�mˠ�1��*;�̇�Ì�A��aCv�(?"a[�k�3@X��p�s�ʧj�S�W��aH+ǒ��l�}�ʁ "����qh�5�gѦ3�<��<p ��<-Ib��\�>᛭X��={@h� Uv+�o�.��i�_ �DQm�9�BLa��&3f���H(s�E,��4�O��/N�(�6q��Z8a��X��:v��9;��g��%,Q�~;CF�c���ʘd��E����#����?��52�;�6I ��ҿjPyT��Q�Wb���_f��Gd<�lc�o6.��7�k.QO��\)eX\�?)}
MI��dn�g�5-��U�pA�f(/q��5H���ӭ02��7��L� ��փ��LD���n��̣(i#.���jfh��Hp��7��J�t�/צ���'����ʫ8k���`���l�>�QcD��j����\iv|e;��f"���-jTZn��1)�3`�"	�����[�R�g��#X
?��.�\�Z�*�yÆ�Y��S��Us=/y�K�́TT<+�q7�ֳ�\m���K�vA�u�e�&��zvo4��ǌs����~������ϳ���A-Hul��=��
�>
���TcE/(< �ID=��x�і'�{�጑�����.=��$Y9�,d�j���@��h(H�M�G��Mꮦ/�5:E��U�X�f�i����-!�z�9f����� �(�(�*�N�6&�#�`��=�x<������K~�^�W�K�+�Y���4`�/*1�}vX�ݓ���׸���ׅe��㶇�}ѳ�����U1�)1w������AQ��k|Y�
�.Mf�h�Y�`*�1��Q�g?�?���W�� ѹJ`�?�E�1�us::�,&��N��Yn�q�א~)ę�l.,d�z��^�*�����a�s,C���0��	���a��u��b�W}ce�١�(P,�(D.��b�7Y�s���ˢ�ݎҥ�`U	����W��KŒ�@������Q���v��,�J(�?��uH���)ݙ[���*KZ�+X۵qr��f�=:�)��s��}�BL�hO�����@c\�4��U���+���I�vhT�������&�Z�ą>��+�Hū~��`� �V,��z~��I��⢉�W���`��ev3.=����W���ą��w�'����]�3�������V�7^��JUl�����`�ߕv�}�X�{����O��~����ChC����c÷�w˧q �A�7�FuG�E�Џ($-�w�|��m<�t���mea~�ȡKm���0�o�W9�{��\���}s�	&Fϥ�yEb���;͚��I�����E>D�v�7�ͷ�7��(.`ˎ��Xa4�M\�!#�7���9�TZ����1]���>����Ά�/m�7���r������%ElDuv� ƫ��ºY�J�e7� �<�P���y6So���o�X�2Ӕ����ͯ8��n���0[��F��|�i����!�I<�׌����(𑀳���3��3l��°��VB^��1����6��w�,�B����`��6�x7?k��m�����!٢��H�67��Z�̂��"�қ���4�bQ��
��\�;�v.dzW���
R�p�O���c@��<��¦햾'g$~���)����Z�lfYELn}d1=�'�l�]S���r?t�W�n��}=�Y9�EY������-�}VDGGH����~PN`�w��z�7{ �B'	)�r����t�%逼�{|[Ɖ�MS�[�o ���n�eL�𩁚�o���R�F����Fq��̙1[>�eu�\_R�bH?^*� V���������eژa��]��0p3;ALs|vVv׀�NQ��2	�~�+CA�^���u�A�䨷��
#��s?^�����I����"�x���)f�C�t_�2�Qf�H����d��<~	��jS������H�b�5��ֈ��c� �� �~3�8�@��s�m��c��f�� �Hz{卂���B&k0F�D��Γ�𦢙~�+�>�L1.��E��o����ݢ�[-V�#"�g�4��!��M�o��G�,�ii :�C��2���~osU�I�e���Ź=�k)h�P�j�%�0;;�`������������k�c� �5XO��z�"�c�K�M)4J#�Z��	ۜ����-A޽�o{!@�,:m���o�mg*Gד������?��j+o���3�]�2�)� ���=�j �.K4Oq��p�{`�/��4���ϑV��2*�BQ�h��*�=O�A��b�R�+���|���Y��}���|���7���'�s�$�?�D+� ��"��8hm�f�|v�9�N��8sgY���=�x4cDHX
Y�.�=[��1��e���-RNm����m6k.C���O��&��vς�$s�ir����7\�?�[۳��&@igj�#����r���?�Mi���K�����_+��%H�\$Y��+&]��� Ӱ4=���7�e�8N�*T$-�OwD�����BM�c�hU�w���G}l�{hC�6�]�_��k�N\Ff��^�6�`R�1��B<��8��xc��@�`��c憻�\y������8m����ٗN4��\:�n�N�0U"����0��$�g���~dm�j/��0����J�� 	BXAY�V5�Tg�)�*��6I�9���)�*���O`w���ko�.��l� ��B���!�jѪSGD�T�.h�Y[��8�r��X�a"#�D�-�^�;���G
 ��-�����J�H�+�Gv;q�d��m7�3� �m�)��`�����D��}e�,�O�V��������c(�@:�R1q�JJ3���O�m�ҳ��V�O��������(�)-�ld=u��i�˱����$ ���}����d�PR���'5�1	/��b�K&t��垅�W����g��Nb��̆΄R�
�xB�^T�j�0f�.�x�jNG�"[o-���4����N��3�/����T�cYjI��Y�V�ںȫ�t�'�J��#��	w��oq�B���R`���3�JzP�2�L��)��X�kAt��g�vd��~�Ym��|Z3l}!��C����\������<d!�0c�(�xO�xe��g#�&��z�7=�@y�]@cd��5��48��&�bn.'�b�x���ܴ��3/IP�K�;���MᎬ�������J���^5S��`z|��־}Oۦ<kI�p��G*��,��	������*/w��l���V�M�4Vu�GRVK��:Z��/�
��zcNjz�s��.L��s�׃���s��qP��D]���+�<ӣOgP�}�pԒ�Ca)c�Y�4�A��������O�,��d�E���v?��y�TC,)q^޼n�T�^��m~�EB_�O�<��(���rF'�2��脣�iv����a����Q�4��Q�oQ�On`i�	+'�G �����h
�ьp^�MJ9��{WX�5L�𞄘�Vy�
�srZ^HR����M��Yb��}���b���'���t����K���o���Uu�|���+�?��;����������ގQ!�	��U�ݨ(-�Q�����f�3F�kV��-�Ȃ��@
,��S "l��4�'�1Fǧw�����h��O���T���N�rI�Sf�����nQ[�����ۻ*�Md��U�I�GӄY��� ˢ�����LS}��b����nU��Ԥ3-�^HQ�.~��F��f�/ߍ��e��R	�e.kL���B�`_V��_���mA��\0\�Zn�#MyY��.P��?�\Ͽn�PV_��њ��g�%��s2�d���x�(�ѿ�%��;$��P���$�{av�[��엚!Pd��o�B�Ug$	8*I@�<��O=N8�Ӳ�4l�Cn��:(߸G��m���ʃ������<i�3P�!��#��}#4�|�V�]�ߚR�l����yT���+Ɔ���R�W�3T��˱���K�'=�ϳ�hJ�������}`l�	D�y�I�ѹ�$֛��T&�i�p��
��u" h�-���u�<4A��=fKGKٖ��l�LpԞ���;�FeDp��rD�� k�j樂��-k��h���W"�,'GY��m쯷ȇ��P���K��.E�\mWm�Y셞ꇜ�v�D߇�}R0k����x��,�?�=�F�e��,≍f��|u"�֯���@da%O��B�E� �}�~���<_-Ğ�8�i�*�A���m����q��"�RT��`Cz�SQ�^t!D07�j5�;V9�k�&9��r7�GG#�w��P�	��uS��%�����J;t&�~Ip�b`f#��^Nh�> �&����cp�b��-�&��"�np�sH�3�*�>.�C��1�	���Q������+���9(?�k���Kk���M�U�4��ng6�:	���FM�Z�)� s�W���Nf#�|x� ��|w�}�xdobU�{i��ޚR�o1�
&�_;|Q���]�N��ֻmh�䖿���2��̝��������h�-l~<� az�,�	���5Ȋh��7��Ϩ��������>�w�r&�jx=�dț}�_G�w+��ii:�뗡� �t�?�y2��-5�Cq_��8+gޔ%p�b�WW��{������{SO���	V��"�O��f����>���w��B�[nWwHq�嚛�	H�������0m�mB��BFnY���>����2,"kE�U�	N�����`k�<�E�ol�_@]��8��+�/���j�/�#`�TC��u]?�+1Z��ٛ�%���ҡ4��E�F��<!7��`�q��Y��~sfE�"͐��e��N<܁�~���l�;@��BΟnZ�X��f�i���a쪲Y�Bc4*X�$c9���5C* �U�gi�sІ�6����Ǚ;���o���j��7vKt�/=#`W�9�������R1�P�j@�s ����eݿ��!�T����*PU�x������J��l�L��@S���q���E���N����\���t��{��&bm�麶���1��=���7Cp�����j����DWx� r�}��H� ��\&����hh,ׄ��JO�r �{\���N����;��K�C̳�Fco�q�	��-�Z���
٧��;]�./�ګh'54��ֿ���E :P�:�;�T�	�eF�U�	'���T�";��g�P�|�&��Swc�%d�qFbC.�$D&P$�i�r�� p3F!�>�LU��/�ٺk0�U2DÜ�VB[L�>zi?D�/�
hF�+{[G�EH��T�1HZ�"�%��m���6r=��6�q� �?㠨��o~{8�d�P�bU1]����u�
*��)w��~�&xRA�H:L�6D��r�	�7��\{bLx�3�������mH����ɨ)�ds�������[R������{��Lʺ�\d2���ܪ8�sk�6��5Ҭ�Rs{2���w��k�
�ز�o-�LͽKu���͗�V�NA!�!����'��oN�&��?�>I�s��ܑ1]�x2��҃:��k��Z<�3�
v�J��]��<S9o��| �J8�^$R�(tq����C���Bn5k�'�{Pt�<�h���w���<@L,q��H{"=�	��;D߮-ҧ�d|e�J�p��x>��l�`H�O1+(똩S�c`�t�0<���0���SH����.wE�x�E��Sm�߈���Q��Vx�Jm���:t�%wE���N엪���=
�0���7}�ү^X��x����\�m��(Ea]}��@�Nk�c�]���u����OP+p�Ѻ� R�g���8�k���KWR���ϛ!�7kOA: wq�g�w��aGS6�$�}�@���^Wo`hw@.QXF>�*z��K��b��E%SR���u�ԆRj%�����������kl<z$-��(��a�����gd��^Le6%�,���K����"�DH�G]c��9�*|Á�]�ןf=��C��}#�^����u�����u8W�h?�����#pأnӡ���.����C&�D) ]���|�p��
UKHn����;���*7���%$�Bx����̉����O��-z!�y�U�G0yJ��Y�|$�+��JDC�碍7�2��/�EY����Y��!`�A����|�Y���}���F�PR�r�7q��o^��-���?�i��������c�Ɩh�0<F���̃�k��|���d�יr�[2�J	���JW������i�U���N�Q<g���Qo�;m3XԊ�����aǐO'R�8�J��3�z�Ɂg�|YNO�k��Pdkw@�ҁb
��Hx��ûjƸ��M9{��֠�AX*�����H��w����j鎜� �$�<��-k>�V3p�T����i`Z��n��k��;M�C$h�}-��Vf�"�A�Mc�������n[�K�B�k`b��^K�_[��n���B�B�x��XP���i����6�O0-x��\����,�34	���s�r��툊ܠ8*���2Ɔ�m��h��d�3v*j\,dE�j�<�0��C3�i��a \7O̺�j�&�D(��sވ���zgIge]m�z.^�7YW��㬄���q� �*QND=s�E�4W��O�S�� �F��7ȧ�T	�k��������m��V��u4{�̐�:8Δ����œJR����P鉗W}�)��ܩuq�#/��y�ʂ༥Mn��u,�z4:��G���j��)��%(�y�db?r{Sab�\�=�G++��7��A��������]d(��b��D3¦7NԔ�m0 [���%�ɢ*'���RP�Oc�:Q�XΖ��6YI8���Y)����+�˪�������,���p�50�ΐ�7QTV�t�b	�a�kW�Q��}��wW"�I�Zq�
ֹ�x
�*�N��W]��YΥ5I��p@�=�p.t،�9"�����c�ub�� ��tx�����⩍�+�`��c8YSʀ K���#�k�cF�>�:�"kz8��F��(D�c�)���@ǕWE�L��$��,�R��0��\��)Ћ���|�ޗ�/�=}n�PH8t�wjX�P�^��^��쭸����̓P7����H��jl��z�6�z�2���m���ʔ��Z��|p\s���ײ⼐`Lh�g1�ҋ����d�W *(�?���~%! �[ ǂ�]��ݛ��Z�¶�����G��B����M�5`<:���!����F��r	�]G�x��&awo8��m<iB��2����m1Md��|�I���Ū�]c�j�c�/�M���#R(����?��$�Z����N��O�t���^�ND���Y���]�O��ֻ�o��"� J�SY���K��/�b��7ۚD��kʍ�jf�Gc�������ޮ(/KO�4�fudѫL7	+'��.��c�U��-�BtIz������6������Z%�V��ê�����W�
��:R�x��]J���g��/����+ݨ�� I��yuK��*����c�	����k��K�$��尮����|�ȑ�V6�
�Bx��P��ޠ�Z���5N4�R�C�L^.艼�|��3���.>�@��xh|����8�w\3R��8l^�����-k��y��1锯��
I�E���`��y�R���ݻ�2�C4^2�v�7��8��^��EI@{@>VS�Ӌ-�r*�dbl?��\����^F��[/����oK>��]$V-P�?yᮨ'�xL�^ABG�p����)���\���0��ƾ��8P~���7�*�U���ݻ�S��G^Z�5�(��+���|"^�3d^�{o
�K׬��"W��Y�NS^T���0�R�g8Q������%�~qU����%�����H�JG��^;3l�1��w�GaѭGAH���{���� �"�J��(��Og�"!b�y�R�bY0BIa�2�8��1ﲡ�ҥf�Q	�4�֟��l��G���vV&[MB|Ƃ�MC����Z���^���^��oN`{�&�Wm�B;�pt�8�<%_(�"Ѱ���gH�����	�����7����՘�L��37s/�#����)��H����!�m�73GM�?��� �/�e���z�"z'2P���"}V��w�yŝU �y�΁�->}w@�v-�ҥ����;A��5Ӻ5.�Uɹ�N���i)		�R��b�R�#������w�U�F�����&����>v�+cJ0F3��^F?'�RW�)�xU ���SSJ�RAX�A�����!#BK�^�Ơw�S�'�L����,7�N�C^���#�B��Z���
q� �V/�����o�WA�L�&E,�j0e������<�Ԁ�Lok�~�$�����{��k	��q�K݆7P8_��h��9��\L+[�J�joߒ��zr���e���[�@l\OR뮉mT��=�+��Y"����v�y���T��"�j���ȡ�-q������<U�ߎ�t)΂c�9ׅs��Γ��%�<�K/��Á���J�c��(<�kƢg5#�xd�O���� r����Q<�>�:͜�^z�r�%�v��g��DҷW��F�B:�1�]b��rR�Q��C��Ϡ�D�P4sD�oO��z����A��p������:���2N��'1z_ܳ��5Z����	��s��]�{�ۑ��Qf+�-�L��JLo$!F��S��9]`K	v��F�N���.�I��͖B�J�߮62�>�-L� � �li�>�u��D(�pJ�Z�J��&s��-�d����kӅc4��z+MD�7�x�|�e�t����`�@o@��L�����P��g�<)[�A�����X��E,i�9r�\���O����7������2<��ޖ� ���w8��H��R�^5FU�F4D0(��H��~�f]��3���?����L��k8�m�EI��a�?f%�6���vu���T����/�&�}�@��[U[Si^�M�]�
l��4"��!�͂q�}h"���������`�"<�kCP���DpmN�R�0g=4{K4�p��~V|#�8.\J�J35��pg�ƾ'��B��<����OR�`[a�ʈ9Hr.P�أ��>�Q���fG�=1��`3�w�����S=��a+��L&�23Է�С�a�1�����NL��w?����fٲ"©��,�M9�ř��ҹJV��vǅP��H!���ƏS֐�+�
4ر�?h���=��TÖ�_g{Z�J��)�$��$��8�}�V�*�)F]xlШ���8I�D}�� f8�-5��D#���q�k�$��t�a�PJ��N=i�t�bZ��FOcso7���l��u��`&EoѱM%����(V<�+F��/�~Ef�H>\ׄo��@���vOp�x��붮v�kh�~f��K���Vfe$,��[�����Q`<u=y5����[_N�/��sY���6�x�P�h���,|U�<���WA&��ҟ�dD飻ҡ���0��>7�O�wU��@�D�����_��^��� h������Eb�! &��"�E��Mj3"�̈"�*�����^��[�ϓ��6���j�bw�����ě*�=U�M����q)�3�8��ŉP��s�op}��y!���̜�b����u�6>��%y�܎a��'����g#�E��$�ш1�!���
���S�Eq���7\�S7G�^�m{�}��u =֡�Y�M8e��#p�ژ������EB���oڂ��(��"Y�쨇�*Y����*��gl�u��K�0�7x~��Gs'/Ġ���E-��Q��w}4і���!�whƙ�T�:��YKX��	mںo?ۘ���&�ܒQtO>6�$ؒ���㘣x���~�d�x��}���#�#R4^X�������=���Ғr�^	�}�rcI�%���Ј����*̾��j:���E~ﺽV�H��
��u��WxM��灡�y�1�ю3}�`U���'gp��j9R)�`ػM��q�'�P��Q��f����=
�� �X���?/��Φ��B�aJ��@3L����E}�OW�"gb�*�;�I��3���p'�!�q��d�J	~��%�p���K{�c��ɥ���+]��/ɅoU0x�M�ʰͣ������M�a�*����(#	���f\b�l�����c*�N`�����Q���j�_��}l02����Kaڞ�|������*yC÷�{Mk�x���ǩ�Tc�؟R�_h�KO\M��Ȓ!b��B?���Z�/��2��mC'��"lz�����S�I���N	H�T�EY�;�dq�V'�ږ��³"�ld�S�Νq��砠� "}�p�;�C��T7��#l��荠�؄��a�)y%(��hH0�ݛMv�qW�+/�uz;Y��d�ᑓ1IX��=��6�֌&Z!��`���{�>~tbO��x�B%����y8���!��Ю�2U�yk���aC��j/�����H������ef�%�g��n%c����;ҌB��Nq�������v��o�NL��p덯/+�����Qh��)�ȨB�RO���w3���q��DdgC��M:~$p��ǰ�yY3Qו�op����/P> �L���/�h��ֹ����-J� ^�7$w�I`�T�A�ʮ4n�h�I���s֬-49 *�w?V7������'��azr?c#=�����R�u=D�����w��V�!V����@���\	�>:J�	���14�˕pf�gS�~�csh���s �d�����]`O��[n8p��H�J6)����QF��ظn��`~OΤ�40���t/d�XL��+�hKw����#@k�!b�����>v�YAл��}��ɁסJ�~���u�')�@ڴN���P��w3������ِY�E�0�B�m�������ݤ���/��T{��X&2�)�S%�鍤 d����Y<\ⱔ4"j��R�:�jZ}��OU!O��2�,J�u�q7D���}��?�}�;)T����ϸ�g���J%�*q��#m�ۮϨ86�cu����RM����{@�%�L&吷$�D���wd���G:e6϶T��Oc���!0�瘉�I�G�)��"/�7|׋:�����aw ��.4'���H�&�D�P�Bjj&T��#�邟�����5ʹ4�Ul#�Yy�Y���$�A^�ΐ���2}�pOy��P��J�G�GH��U�np2b^��-4��T��Z��W���	S/�Q���~M]Q&_MV�7�[+�̱I�����6�$�L��qzj�Q,�D�Wj`(�m4c5��<[]z��&���K7�une�Jp��q����+?O�rc¨�P�:��*��jw��=MF���w/ g�X���pG���M��n��)g%���5_�Syrw�#b�������R�+�s_��<W>׵~���6���G��զx�*\@�p��#@#˾�@Vht�[sU?���ZN��m�e=\P�X%%�w#�ϧH��*4���!��6�@i��K�b��^�u�8���f��zvd��\@���V��Z6�7�7/�X���lX"���P`�M&�r�}��!�Ec����/���M��mD��X�R���k��x��1��2u}�R&|��P-3��[ZJ�꺢}�ک�r�eI2x�g2))[k��B�:��N?Y}�/�d�Ǭ�´�ҷ��1��9S��%dS0I�9ќ ��!�}X���H��.��_�jFz��Y
g�O'S�0�N��l$~i���ݻ�8�(
�m��F
m�Pވ�s��UY(��wFk{�������_l�����oy�p�?��N:�m��g~|8���ps�/Vj�𘉨	���x��l�ь8�{QA�!�g��a�'~��NP�CU�W�����K��/���#F�T��fء�9$��rA}��E�}%p}ڣ�h���0��
C�'��>I�K$�"xd ������I7�>toY'���+4ү�|v�ֲϳ��;f]����H.`� m"4�K�-��菳�E��t��5����ҫ
,n�@�a̲�,` �j��,��杪�q?w6ԇ�Rx��Rt�I#	���M!��w�u24m[�}2 <0��3�]!��|��a|��)t���K��W�R&�����{yF���!��b�XnF!l�@	6����3��Q�3���Eߚ.i|H��	r��~���@��,��7	��?׸�9#�j�3�8����܍�J�B<��1�ٲM	@U9j�S�̺x�(e.A���`�N��z�s�(���,x�zB��n�|�~|5q������k�g>�M[|�B��	y!�+e�e`7SG�}���a�s33l��Lb�D�Z4H��y�R�̯U$���؆\	�d��ak�i��̺'�8״�D#�mOT��o����5�!Ĳ�(��W�)ϩDT�E~|o�h\��x�ҫ�@k6a��E�K����\q�пV�E�-�wv�vDk�%q(	N�j� �i����@���$���|��TlBC�(<�=��uIk9�|2��D�vz�<?/	���9�}�q���V�(�	MX�#��o?�ưG1���u���Ɯ��;C(���?�8�6�!X�o6���ӄ����'pOgZIz��F=ws�ÕUZ��`�B�%7ڷ����u�:T�����/�[��HCi�Kͺ�d!�u���\ ?��K�c��Â{�M�Q�8��u=�>`1�z�>��q;���Z�9T����8akȡ<�b���;��&=B����`N}@Ʈ ���l$���<nR����AFq��7�,�I`���DdQ2�68����B����
!���|ba��õ��HCz�g_kd���!�MɅ-a�/F�"˱4�n`�B{��!0V���gr<�����|��ы��	UK�>ޢP��q̾���HW'K1�K6���w��������?���uV�� J6R��U��qڴ���b����A4�%�l����B<���0�ʑ?����wM��z7S�*qI�g���$��~��5W,��aCŕw;��P�@�󢿻-��:��g�hn����	��
�{QX)˦a�� ��v�L�w�Q�F	Z�)�l�6��1!>5*i�l��w�RX��}4�����jg��8����)�� .*�sOz�Yr3F�D�P��%�0�F�=Q�"]�T֠v�"�)/4Nm�2 D�Y�(�N@T����d֝(pg��a���\�Ӆ�d|eB���U9�8�z��F����i׻��#������V�TقV�d[ڷ�_8	Ҝ����n+�	��ܫ5�0z��ՏP�:�)��t�\�_	^�T���!%���C}z�6L��L��K�2U���.!���`�+$E��m~�oB�Ua�CmT�� �Zv���0,��I�ڳ3���?h�x/˳�'V,d������7ϟ��|]��4 �"�H��dKy��&����MoZ�l=�1����(b���E���.K>��G��(���#Z��5���#�N��ٚ�`&�ú{���u7GX��%��x#���:��u��"��S
}�C+����p��5�W���� ���
��x̞3 O��9�� ���$�ࠍ��M������,Y�T����f�5��⑹k5�µ���\�@��5��ג��W��>�a�|�� ���s��#{b��:h }��!TY 6�y��O��6��XK�Q{ޭ�;�v��P XGL������N�u�1v�t ϊ��x���9q}��o����C
:�G�k2Ľ=���N��<a�#���(
��2?��r���ݯ�y���\5� �F������1/2p
�Fk�5��-H�䄍����(�⨜(�/c�:��˪績��S))y���K1�2�Fn�o�V�����?-/��2>S�����C�OطWXϚ,
��F���K��f��|>ߧ���:� o��o�i�	Bdd���Mf���+Iܢ]�.�
A�Jr#��_����bi\-}�� ��-����}Ս}�&�Hx�l�7���rd��(�*(��ꜗ9!J�������w�Ψ�25���e>f�/�`ѳ��؏���G��d�NJ��h������YR����u'� �:���{3\n�Ӵ��� /?�*�5�^Hv<o�,H�ܚd;�Hd�P����K���$F?��%�-K|m 2Ndk�@�T�&�{�y��j�=�u�D�9��k������O�5�A+zY��O��)k�tfo��]�i��P���DTM2��O(&�w5pݬl�-3`o>�i (ߨR�a�3�3���y�����p�՜�Z��"�T��L�յ3 J��аRd�V��J ���ԭ���
r�j�4�MI*CY�*%�Ws��)���f-�v���u�5D�2��M��Z��H�(�U�ki�53/�>n3 �UƌQ7wX5zѥ��㴁�<KyW�-#i��
�i�,�R�k��ǽof�=k��4cj��-%L�T0o��X�AT]���vF]�ٛ��F"I��*�%���=-��pȭPb��L�[B���j�%n�b�6��E�k$���餠����$x�/�haz��o߸�U��E".%��"�V�Tß�d#��9Ւ�+
�8j�ɻ��l���f��	 ��B�ԁ�1�kF`�,g�o6�J�V�Pn��nJ�[{9Yo�7����������|?���y,��so�#�wڂ�1V=yq�_����U��T�Ά=ş _��'�6R��eDN���6M_^wr�F���m�Z��0Pz�oOI.D�'ID[�9�x��[���J	���"���>��F�g�-L��G>��Í[���&�ʡ��o�]w����Y��.�#/4r.A����a�٤�?��T��t�UľdL�4��ރ�Dlj�l~!��]�k���9
�xBNi5� ����������>K��(�A1:**����y�3%����nv�����FÎ�/�QG�Z	^���ƚĤs�l�
�<=��̈́Z47e�O2�U������z�&	 �pK�<-k�"ý�C�<�F��_�ڂ�j	���i��$�R����hս�Z�w�M���|Ҍ�3�M� �}����8#�Wu������	�����Ҙ�n��T��]�j_��d���ʳ��ɆF9���$���I���
�p��i��<��F�A�k�v�#,w,�LI8��d�i5��˚��.�Zy�Ւe��!��	4yۼ8|;`,��BW`u{���_�_�{s��0E����htD�+Nh�t�'R.�O�P��(��m��ɉ��b�4�?#�%��?�1��>&%��~/����va�-Aj�p�ή�}�sQ��ԉ���+�G�1dH��,�c��L�a��T�2�Z�Ǵ�������̽����u��q��rn�Q���i�RX^�^��gC���s7>�b�������?��*�n	"鮹�
�_R����ɰ&1d7��a�4J�u��d,<YW&n%��Ͼ��̌|$q��*���ī���G�=��_�U��n�Vw�:G�x�vxn��^�Ia3E��2n��l�A�����(�v��G8��I������!��ɈY���m[B��v��Џ�?fJޔ]�T��S4�V�ʑ� ��"^p�9��i}�k�Fn���ֲ,κ�^�Ǿӹ�VCC^���S�<���)��l)B��~�.!q�oO3ـ6����$���׵n�E��{}A4I���m�H���}?#B&;�Dǃ�y	Q�r���K�պ)pi�1��g���LWo��m�B�]�dt��i�$V7b�2�p�wj+Q�`m���r��^�U`"%�y-��K�j�_�(���/};՞�AM���ub���$�����h)�a�u�$$��x<NÒQf|9)��p�5eAI�7r�N�D۹�M��d2��� �w|�꺍��)�h)��f
2N�0��u*_~��
��U3����D�]��>�1$}��D4K[�M
�����2��v�z��L��U��|&N�'+�S��2�-�n�A��8|���Qx���e6�fT}�F���v���@B�k��"��֪ ��d��"D���ƞMP��7��dX�f�'ç�Գs�<Fʂ��{~O=?�߇&��hE�Y����=��_��cY�<����?p2�S�wT��Lx�j�fpd��M�3�ǈ3B��F��k'DZ�x��*e����ž�!	Z� %b *���ia��7��m��(O')�8��Py]h!ܛ�2�Ԛe����p+�(?����SZCn3Ǩ@Z�D��f����*;��Ϡ��T���� ���[ҫQ���;���m������{������?ߘ�̃�8�Ф��cUa㮺�|������F ��h1��̣��e���|�`1�O�s�3w����Y1T������l��̐��S�LX�(GYf��5U-��kG@�>�b��1��2��J�1ө�h�e���⳦�Rf�w����0A3 S��_
��U������΂?�$r,�P��γtP�@���A���?u�u��]�Q:E?k���!RCO0{��p$���e��3���?�_�ѧq�� ?�t[�"�%Ϙ��3ـ��e��ɷ���
_,{:�t��~�w�i�B��Z���{�7M�<ds_�d�A�"��2����i������!�l�8+I_}�P	X�l�@$���X�FL�G�oЃFW�7L�űȸ�u���"Avi� �sb|Ek>�pK�2s��ii
 �o
�Uͨ-����W?��T�/=�kg��~i ��I��+ǐ��+3N҄��B�^������S��N{�R�w*���ܼl��[���#��~�b��|:���;>9j�n#h���L)��97>|C�6)7}�Su���>}`/�\;���V�J��z����q8Z�v�m�od��i�w�x=��|o���� (��N�gۇ��*�#\ܑ.;I�1l{��AD��u�){������*ǻ��߅)fJ����vnF�Dq�ٖ�i�$��u��?����F�9�1Sū[ C��e���0�W~�z����jXSx�v[���Uߋr��7�����O�A̻]u���񅵲���9RO@�q��μn��:�󨺸������l��q�'�O�	#UQ�HW���d��&8דAԻ���7�W�>�/��v��Y�b��>Zed"Qg�o=u[x�`t΢`��6��Ng���(��zĿ���d�^�e�Bڙp��{Y�hye�c��|�21�̗�����~|��/��+oj�xr�(-����keO�߃4�[��Y�ׅ�����JbkֹXi�X��V`�I��~��8�?����~���%��CW���Mi�SM9�M��'a#�;�>���Y�/�!�%2�ł�p���z�C�4�?#�T �f-�n$?A9!"��(5^��j���݆��	�^F��C���F%��ҡ��	�6n�VM��B:����{�@�4�وJ����m�	�P��-B>�3&Q��F��0�夞U{�3m:��2�Q݄2_Z�#��*O6`q�CG�!��!Nvh��t8\ߑ�j���d�Y�ntä����9Ih�l�8	�h|̉�iʇ��l�kX��k6�����%'�ݗ�.�[&�~���q�f@��N$�>[i-{[P|<�rk~�긊>���t_UQ��W�9�ze��Y"�1b�����0
�>��3__���I]u��z�ݬٔ`�hJ눍��׸y-8jV����w�`������3.幊W?M��fL�%�(���|(B��	5��3:�~	4s*zG��3_��,N|�n;B���+dI��ҿe���ֻ�]� ��Bo6��t%�auB)���7'�d5��׋�k�۞��#����}�ۅP�ۈ掿�&�#|��]Fc�+�<P��?�1k���/	>�W�3����T�tB�S��R<n]B��_�L[�������)�ZB�R��1$�+� ���C Nn�tDm�ɰo���"t�������o��'�@%&�Q}~�^�t��N9E4���!�6�U���=$J���Պ� �u����~"��л�B��Dj�U�J���U�%W�F(����5�/f�B�yc����Z����Rs�G���~�����bǃ����Yą*�,.�=J�p�n���:}h�zWhPE�rF�k�	��Cn8-�3�p{Y�'�a��VMV:�UE�6���7���G�&��.N��n��gk��,����^�tN�F0�(�1.;�o[�����#�r�����#�6cn�.��𙟢��;��c�it���<���	_{oJb<�h����Ճ�u{_}ȝk%�N
Y0��i�u6��?+�@��]�N��`����h��
3�G>M��[.A@����?@���Da�P�	�)-8e�X oҿ-������h{Z3��&^���Lfre (ɯ� X: Z�>��{{
֪��Cf�cu+퉑�?���Dv�Q}�/:�i#`���\�q��_�s�5�A��j�r2��;��5��Nd�Zi���	����̫��VB�3*�EA;n��$��f01�"TIu毳��R� _r�W¸f6�ۢ2�@�C^,F<Z��0�6A�l������ķ^���5m��@�?P_��<�t)~��GO�xb[��V�s��VU6�=����2�z3�<��J&���@�~�q��U<	TgA��&n��NM,>٘����z�����g��_ܞ��ɧ���+�yظW��|��:HV�RΞ���0F�~K��:���-�>$ip	�S�Z�D�̟��i�HĽ{}R�����;9H����K��h|}3�o�'��m*vu�8a^Pá8))pM�3sMk�B�b���)���֛T<78Pѵ_�����ٰi(��6F|.
��W��� ��T|�z��8]�K��|k�SX�O�ٺ���T�B�~�;x�Lj��IHV������g��Z�jj�l��.�-��Ly��U�&��>Esw����|S�^����ئ�y$�%P(nB�1�'���v��-�d�9jd
H�Ә�\��,}�8�T�~�i��'d�OqI ��9SM��TffIJ��8�"Um�J�	|"�/�t-�H���Щ�u#��'n�.i����=O��%M�E�1q !T���3Bs��@���LI��Y[���)*h�U�3^�	�;Pnu��]1|Dsp����&wF��R��r����fi���<�Xn�ƿ���̣�s-��KzJ���G��<�E�y,U����������L���,Sݰ�WlMfε���gR�Lq7Sn�$Zw3�	�1��ȃ�'���V�O[�Bӵ���j��u�St�.��o.�.�f����)�����D;��V�.,l;=�O9��5��M���D�%��zo:"��L�Y̗T����ZTգ��ݚqؒ��*n�����������p�N���P{U,.�=d��^�ƚ-�݋K�f#:̙}���ԧ���� �TWN/`0���hV��k1X$�~=A-�.����r�5b��fD�5ܮ��ڹG|*��'Q��ӝd��y�K^Ά���t
��3SO�4��'�ɛ�Rb)$q�%�Jj�0�R�g��"d��S��i���h����P��<]��Q�Jk�zl>������%2>k+!�#X��H1�|P��A*h �:VۨM}!͍b �s��k�I�H�:�h1���z���N_�D�;������@�t�I*�b�����������!S�F*Z`\�:�vtLzdR����4�'ʶ�1��O��Q��6<��\�����r5��
&�j��p���	Ѽ�j�iH�����`�Xn��,e.����w�6��5����zR��u|H��82fڶp�1ԥ�%�K�1�r�/ݛe��	g񒪖8u	��k������&5�ޮ��3Do���m�g/���$l��3��~#K�c�ϐ�Ĉ~=�c$����Ȫ[���=ڡ�Vu� ��E ���6���
D�U��y�}c�� Guu���j(ѩ=��tI���� �<pX���7;�X3Y�z!3��u�����}��P�X-��S�ou�@Rz�}�*'���
�́L9�����=:����b��e#�p���,��2��Ƣ\\�Fq�! ��(������m!N���J��e# r�Udl��%h0?�H��,��U�(�7��>a$P��v�e	f�ҏ|!�Աel��{ս~���qq.K�%;�v�s�RB*�$'kEB@�4#f׸�w�����G�)�dXL V��6�O��ʃ5}��HO�r�{Ԃ��*�]�j��H���p�6�����r��x<��t�5w�U����ƴ�����$��vp�S��;����!g�^u�y�{�!�g�����%9��A���Hq-��_�?��nb��yL���	��{��'���o*[���Ie��<4�^�)�P?��������v[�fTfaO�O�����k�^T��ú{�B�f%wPm���ѯ6���uI#gs�I�G��n��~~�2��ub�W8-�cj3��ABZ�Y�Է����'�~4�'Q����X���S�q�t�+`���/ď�ue�����e�b�>P�9|�CJF����	�T��	�D��4d��MIdo����G�J)X�t��컗�J����8pd�K��;_`���DH���,�Rzf3@��P���M���gGئT|��.��,�Y� 5����R����Qw��Y����۶c _�mi��?�jQ`-�H��f��T��>qI8.^V8��5���,B־K�ƚ%���iy3�_*et ll.c��4���$Rƍ�i֟r(38�7Z$��y���&6t#�Ξɓ&���w�B"P��R̴m]p����i?p?b�.Ŀ�����b2�gk�;�ݟM��Dv�2�xvڡ��E�Dd�W���&ϥ�E�6�(\�7�����02ي����[����9�癬��&�a+�;��`��Ak��<��;�*� �c��	��cCx^�a�2�y
bI��2�9��kJ�RGh)�/��$w<ɼ���Yq"����$ Q��BK�^݌#�Ř�7�TM6��X�"EM�g;��Y�Dk��vd�܁��}�5�M^Тo�`8��[n 
� �?�<Ii����!ơ���@;�s�L�A����V��J7x�DY�3_������BJF� ���&j�AE�6��)$��_%j���j�gch�*GV���GV3�?M������s��x��5�����1��O��A.tl���_���/J�}:2�c�f��0��F��Xm�h�C��!�Luv&�������<	|�I���G�,5M]�vv��	-��U�h��N��_)A������ݷ[em�=p(�_i���!lך����E�y~���_ �d�m|6#��/k���.�E�����n�$��Y�R����S�..�����{Ay�Y�ҿ��am��7[�1���QVZ��JYH72]@����	rb�I^*�%jw�Q�0�r.�ƨJ�g��]8���M�������~���~���l�wHG$�>����M�r�k���)���RC�f��,9����I���g���=�^�Af�����Pۤ�r����b��Kb]r��q�û{���h�M���=M�wu`�f����dv�e��)���3�<%8WR�AD
�"�:	��o��nA��Vy�ᨯ�i��ve�M@�������9��쀠�ݿ/��ݣ`�ʛ6v��_�k��%hճ�ϭ�ַ�y��D��+�6��2V�����SW������3��?�!5vv=O�W/�s"���W��	�1���u�u�Qq�(�U������ݤ9R~��P�"��p�ȵB�0
;�2�ai�����g\V�^k�������@�yc%Z��I���ag+�'�>}��`8�(X��rf����t�uK7�SQ ���񫱂EQ��?˩�w���V��a!K/�w+N���f;��w��G�
������u!��_�0�e�Q��1��8u�eiÔ�VY5CqC%.@P�"�;��&�f$e�A񇕣��wzwO�Y�
1������Y~Tk��}��LQ΅k�D����F%	%T�|1�	�#�\̦d$R�F�Z0[	uG3�� fˢ��U�fL]C�]6�KnK+U���OUI���E7Z&SIWK��]�������qL��e�8�	�擧����M$��u:T�$����;V��t�L��f��t/5L@��3�b@��C�����\�K��7��~$��ɹ��T&��,�Y�s��Q��6ݪ'H��O������OS�F��B��!�������L�`�b��M�qS7Yw�L�����3ʓuO��v�^�`%���b���W���"|�E��,�6�>E���YU��Oߞ�1x���˯�T�<P�U��jSt��[����Dh��
'���((�{󝈏���%�@p��!2��=�C����Μ^9��l���Ț��"�ơ�7��%p�hӭ�ΐ��#�:$[����Rǫx�������+�X%dۈ�O�]K��nꅻ" 'ST[����T��`���׼�������[��X�Q$�;TX�g�	ntb(�Z��׷�������7�a�B! �4�&��7b������26U��e�t��M5&�=����w�Un�����9��AZ2D��xq���ؗ�ce��<yR���B���dtn뇚���	���W&MN���xo)	�R+m�z�OF�.�Ak��v2T�o �=c��]P��e0A\Z�h|�L�yF8��R�Ϙ�bl{s<Yz��q��5W��_cs���$�� �
�1�w�WI[8a��_���T�@Wg��-�ZͰ[�ۭrM\���������BD
�:܋��X��N�O� NI��)�YR��Õ���6����G:�W[�ut+�Ҕ���B�T��6QQ^t��0��8]���P��ä��tz�W�k�8\�Z-j�~�6�"��M ��E��dV�l���@� ���s��ҙ^��ii-��דR�K?�4F�8^�.V�	8UZ��aI��v�NJL�
Pt�CK�u6fj~�-��u�U�Gs�+�x�&����A�19*��h��A���k ߧ�T����I���2(\��;Y6�e�&x���3%��ie�0nF(Z���(-De��X࿂�r���T�+�V���o5��|˛�-�pi�cY~5���[!��D)��F�U.�K�����q�Dҭ���oBv�f�/FkV�#甴b@�L��\ :���'MWic��~}T���݇�X@"�T^���{<�N����G�9����|4��#��Qqj����]���MO	�j�=�Ew;�	��E����a�EGN�m�w�l&��9�	�e�5�w�ꘪ+$���.@�J�@�o�$!�Z�_�ܓ2j:8���@(BM�-P�*!���>(���`��K���ت�4v����0'U^:R�Ⳗ���Y>���}9�s�{q����RҊd��4�$ ��Y$J��s�����l[��xء�~nd�B*!X�1m�ƣ��A�$1Kqo�AL�|jEQ��z�*������ޖ�o'���>W�e��B�|��Tx#�̔����(���t?�� ƍ�����(�p�i�it�ٟ5��"M���eT?vy��ٺ����L�8=�iDW�X���;��xς$oyw��]�%��"a��p�������<(�&���V�\�Ӏ�s���������������#��-kU�ČW��^Z7H�!'��^B��n�_��C�2�����(�_�DM$>䁚Ko�}D"�ߚ�v���ؙs|ԃ.�W'I���q��Ň�璈��WE�1�e�=u������P�-����\��", r�1[׻�D3y��ꪠ�?���K�t��V�� Sv[���ҖkͪT�,��Y��'�s��߮�jPcC�V�-�3F��l�r%��R������u	�>�T�`w�Ml
����)j�g���B1^8�R/g�f�&����:���~��_ܮصժ��V�2"�Մ<�dy���̡�[d�S�Ý��+?��禗�q^���̬*���0�(c��c��
����O���I��[�ن/k�YC�!��ֺ&%;�k�+�I�,����(�_0\pMurq�z�W3^=�c�M�	M��Y5A>l����S��*b4Ә��Z~&��Ϣ�B�$�L���6v�2ؤ�g7�i��'0��~"tv�N1�Te���ǎm
�m3G�y�d(IVb�3��,]9�w9�-�8�u�1\���s��!��Ve8�K뿉_^֥���a+V�ljęX}x���D�+��?����ݶwz-PvOM����S[���h��F�����H��j��&��b�䞻�n�������Ӑ�Pe[Č�@�c[��p�{%��E^-�m0(�%Ԩ��ǟoz�|��M�H��1l�h��ǯ���o��:eHr��quSx8�4t����t2ξ �C%��[Ծ����!���m��~~$K	X��BK�%�5Ĳ���-�����x���%1r�傚��TKj����7}S�߾ ��!�^0����\C�������}���퓱Q􂨿(���$%��2Ϯ�y�,q�yN<�wO������v�τ��>�X]�����Nz-�|��D�~ʵ��]�y�#��r���tEį�r%*�Y{m���P��:��:�����i�B��[��v[�6c�$��s�!�R˞��aY��qN�ԸH��E�f��`�N�	�xp�;mFz�иiRI�qG3�@�IR�;�ߏV�[tj&�=,��y/�$�+TG8���,ɗ�kSu���v�N%͊|���G��+y#|��=1�.���
m+��7�@�KE'�W�Ҋ��$t>�?P��޸�u���s\�!��U�`x#ռ]��dH���L� R�Wȯ}��IWZ��PO��(zU����Q" ��U(Ċ�yBQ <XE[���&+"��{�>ڂ������$I2,���φ�Mb.U�����ӕ�� �|'���HUy�H���nV$��|��Y�.�P�/=X�U�-�p�C��i�����,�J)u�?Ѻ�d+("[�)�������f�Q*b�D�*=L�O��0� �t�ޮ�o�c�)�B��o�����G��ؘAސ�ޯ�|9̭�w��{0�����UB���A��Ս��� 	��m�f@;�7��X�~�)�$����~ D�Χ-��3M	;�R-���ġ³n�_��BZfX&���..���Ƚ�I��Ѐ@���-y�J�9���T\_ �M�5�o$�uh����@�0vw3#	�(���&|�7�e�+P�n�Ѯ���ΰ8+qV,�A���i��[�G	�d�ꢭ�q��.�nη����!H��`_�T�-1~!�H���v�H}������7��'���n8��ok�)��rbN%����z�-��u���_�a+\o���.T�H~��b���G�9�M���;`�\�LQ3i�,���������?��q��ۊ`E�/��"p2�Gpr�ҕ�M77%F��5V%���4p���j��h�ntl@gЃ.`>'("�x���fu.�'JF>��y��WL�`�\&��s}�h��g�qu���G�i�#��S�7�r��/�f��\�2>���ʽHu�ʰ�h?<�2pOꝛ��K1�'�|��t�E���=b}t�j�;I5��\y����b[ե?��'՘��c���%h|KWzP�(˵L���e��.M@U���S���w포W�Ch�� ����v:�w!� (�oh��m�S��;15ӌ�K�ҷ�c1���e�+%���,�V�j��� ������%���B���F�s����Q.?�g�r�ˎ��y���*	�As���ZmA=0�|A��r��?u_�?��������@��8������Fqa7ΰ;YG��r*�\�����i��3�X�!�?��m�8���^�U���^�������
V�ciV�E3�J��n��V#NW5�)�Vj2�SP�N�=Q�g��aik��H�K�]2o�p����{)��������$.�AG���[��pS�E\eî� C@Pu���m�	�j�3��1�����1�m�T��?�ͺ�$��|����nN�eo�7�� �!�m�[���B�-��lyt�8v6@�@D�h2^n�]��.w}������#5����kHU�g�!(�����7/�U��A68�8,�7J:��OB3V{뿻+p��7��H'�|Dt�C�:���z��w�E,���:�[�%Ģ6'M��N�3�y�����/_u�4��$k
��@�o�U&�6�k�m29s<?�`�=k˰�mu�;�(:6��m�@��N��߽Ws2tы��Y;yL��Ϊ������S���tux��}I��hd
E�������xD�����Cx�s(r���-vÖ �M�r[�s@ȟ�0���d�ƹ�ٯ$tmV+�r�O�-���Q�#�Hl�]�5У��!�5�F����@�r2}w�X~~��w-#7���yi�Iȸ ��ҁ�<=^�����T����El�_�N����2�!�+�K�pP�pX.����=@��	��%���5yl��!����Zʏ��F�f��.Ĉȅ�
�*�����Wm��i9o����)�r�����r�N��	l�u��ĈAkه�lc����4/�hE4޽v(Ͼeں/��iRM������WmŹM�c��4�Q7M�V{j��D���5 $����*e+�?8���:2�{�B*I϶{* �"���V��K�u腷 �U`�y-���'%�Xr�����A!����^�'0��9����Lg�}]���ݍ�<������vq����W%�s�9�����#{����5�v��[��[�e���)7H�5�F���o�io��Îք�vu�l���m$���D(Y8/g���p������)�}�m0gP��Dw�QU�� �n�4�4	�l��*�%����?𤉀�+��U��,�w��)js�:�_M�@���m�E�Yywk��WS����u�Z���|B��/e��'1�*��lw4�^�دt��NCԉHmL��?{��XFGb��o������g�!�����z���(��p"���Q�u���-R�|�ok����B�+wQ�A�K��!��>�����ҷ�e���}�ǃa*�s�{xW���R�''� *���-�&�{<�yƼ3�O��v����rk�2��\5���9��"��8j�Mwj�p)Ξ���&]֌��U/�+t�Lr{_�<���EHPG87U�_�QvO�c�/M����d���̳}�E�?#�`�M��!�"
�_r��vη%��o��=8��ʎPt�!��Y�V����������gA�Y����6��D�dK78ko������5@z�4�ش�W��_r���.���>�tV�fݫ-��Ǣ�5_�`f(<5��i=ܝ�b7��L�x��	i�z�"�
�I��;OmX��Ϣ�:#�r��W�z ����4E&��tO�밒�د.UT��-��i��/']�JԄ����C���7W������y�(��h��2��q~����ߤ8���Ľd�e���v}�)p�k����;��])aJǹ�-��r��=Ny�e�g�/ky6�h1�X5H�H�q4��/8A��C�^�e{�8U�Ҟ�����}��-sb�{�nh����Uʅ�4�1.w��|p����m?�ꡮ�c+_��?�F���,���Ia+��d,��fn�X/�7oV���(P�r��ri���o�#�N���PRٞ�'>��YQ��|��6]=Q=lH�]�=�(�Nډ`��JXYbH���6�$Z�w�Y����=)#H�:�X�v\���Ov��;���1+���Tvf��W�݌�\��˼��cd�70%�ʑ��̌K��m|�Y��08�t��t���].O,��Xhj���zD���7}��ϗ ��� ���'��&}S ��a+agF4ӛ]�En�Peg���_ռ�m=L�P��7�G����	R:�^������;з��4��H���a<���B�t��m69�k��p�X�W�K6�&�(-�C3f���)����B���� �.S%�N�˚"������z.s�4�V�s7���4�]�;߇9-�?s���٤�c�e ������]�o=V8��
 �5�a�q"�0���\�3dq����sV�H$��t�(7��<r�xWua#K��D������~u�����/F�vUbH��{\�������+��7�	�V��T
R�����8]�����l�$�<��vQ1��0�!i�c*��yF��ǜ�[	�}ҳ�v��� �5 y�sU����#U���@E�3�ع4������ɋ$�����5g,�fP|�d�y}Ï\���~����\O�0R|I���t-��+_���ý"��ҷס&D�m��?j�-g��,Ũ:�7IO�Q�ZԐ��9y�il7��`�E쥯��w43H�j�@�#Z���CC��c���_D/�3<
M��*� �������