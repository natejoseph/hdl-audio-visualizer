��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N������ư�_X�[I�y͘R<�X=�2Ӛ�'Mt���Dފ()���9^��S�,�v�p�y|�����w� �C����{��j6&6�tb���x�'�$2=�7��/�D-e^2��:}����l�~�*�\ۇ4U*�q�rk��C��*6R�WT^n�V̨<LGZ��W]�j��;	��r�5^������z���"W��� �$�z�0x����i���1p�����W��bV{��_1b���jTFؖ4bk�>p�Kd�T�o�Pf��)�z���PS�W*34��+ x<�BU�/p")&8�q3�7�������\D(�y�m�?:o�e���^��RKQu����xZ43�Q�$�:�S��������N������1��~����8ӱ����	I����A�!lղ���YV�Ѵ�(
��k�coѳW�q�?���﹮+4-W�z��]�\�nKD7�Ȧ9~�I4+W��2O��aQ�g���1��tQ
U�������MH�x�Na�����<ؿ/�yߌ�M]1x9"�y��@$6� ��� %JB(g�8E�U `f���i���/�7��1$����ءCŭ��=b~L�kp����%(������^UI��86��\]����-�=je�;R���y�԰oP.冯��ǳd������ybnǫ��[!���e���lEfs�"�B�u���f��<�0PuL7����L�ٜ��c�n2����x���%��}!�M!e�g���'�b''b�oZtȤ�� (�2��jo�AH]f�hs(T�/2�����#'x �u�$�u�ۯ�nފLE���h	p�h��z�(շ�*��6����Y�!����b��^:��(W �<�!�z;�7٦!�N����7�W}4�/�%` ���$�ء4�_2/��rՖF'�����m��)�^��KxD�(�;��K���F��.�>k�9?86�3��(M�~+�El���G؋�ʸP�6h}��v)i	��ڋY}g��{�F�U-�GQ/Ah�<�O�_>�t��@�"�)'�	b���5k�`���#�&��h�jr)Z��:���� ����um����ы.�#1�M��o���!j�R��x\�9TB�`�&>Y�rn>цɇ��V�UmD|C��?� �P�K��'�`Q�=���n�2��.���cA�W��kڴ��Ĉ
�.(��`�<��D½����M����3ǣӉd�"̀��c6����_3�n:2��+����z��ap�K���YK�!��O�W����S>n�����R��\Ш��ҸW�$���BK�����]���j,��q@�f����&�8׎m[2 ���E.�A��s7b�V�4���ǲx��+WJt�:�q~�����׉'��w�N�wi�����܌�u�t�S~ƽ����������ؑPԵ��"!j�Ep����%3J�����7� ���I�ڄSF�7>�Ȼ�V�P���dU��&*�|:���-(#��Ґ���(���)�E'P�}�	����A�"�{C�����m�����;�
�hwZ�s�-R�z?�N�RKʤ��޸��-!�5\�đ�-�o�<<Rx�:�]\�`���p�i�;d-�@��t U�U�h4�F�mT���fz�,���8�?�c�qq۶��&;&&|5-�nW<aj}��������fz'8N1�H���I�p�фc9�aA��W,Րl_5O]J�PD����V��%Μ�X���UeZd5�G�d��ݥ����1�j���z�#ګo�}J��x���O� �ճ����� Tv� �?]�>D��H� 2f��u�;}������G����%8�<أ�+|G"F����K�`�8,�[�N"�?��Z�T�"����OA�zLG:Y����u�K�r�L���Q���tY��E(�­�� lF��01�g%tj#��	�p�⦢B�2��1�Q�C)?Q_1T�*��,z��erFHRS�N��L�]K�4%CgY��v�V	t�[O�������q`��"���!K�4��w�#bn���pm�C	�*�c�e/eʗO�E�p����jH���8��N%�T'㇡�%w@��n}��jj.����ԗ��+�~��b����U/րv��~��{�z-����񰰮x4%�\Y�!�(oE5iW5��do#"�U�*�(Nq�㢝���X)��(Wa-�fXSE��S �W���:����꫅�(�X4)����u��!K��u�O���K
�~HA_�S�ߡH.������ �
�l+~������R虲� �@Z�u�U-�V6�ŷ���N�����^��3c}��w��5��}�H���K�}rq�)2S�Qݲ�� �0���B<+i�g'��גșH4�v�~휖�T=_��.�g�h[qz�������qdb&�P�+���[m��H������za	n����dž�q� �p& i-]Rc>#�WS�����h/�s>b���h��D��n�����L�K��M��嚾�׫A�&�[�a�x:�`l�qmύ9O�S?�O��e4�uK��^���]!Lk��/��ϳD��(��A����rm{������l��q��g�=��l�yЙRb	]z���.��!Nu��j�=V��❮n"o�?�; �� �"��7e���g!k	�˘�U
'���وno&�^(��@�?��J<{�q����W] �"(�������l�r1����m�<o�̃��y%t���4a��2_��t�����3rpúIc�K��\���X,���� w��d��ܢ�o챰��@"����ʽ�@!�����sTˊǌ�B5��& �)��&����c��=<�ā�#��k��~�l6��%�w� 
ۭ'�s ��H�����Խj}IL�X7Jl3��(B�w�t�LΒv��ٝ>��S���v����'+Y���>��`�1怛		שT�p˓Bx�@�`�J���;L���/�cshT��:��[/e�lϗEK�Ӳ�?����c�#�:9b��%�)Z�	t2�'�zD��9�������c7��r�A���B�Y,�r�[_�
@� ������@�Z+���Y�^�Զ�Bq- �-N+�Y�G�B׷�)|)/0#���GA�"t4*e�b�>P�^_�c���0������+M�0�P$Yb�cԛ<U�y���g��؄�=�3L^��Z_�Aކ��rt�+:�6��l�L|�0��\h]E׹S�?�߹#;t%�ӞI;J �mJ��*�a$�zz����[!OJ��Ez�H�ܟ���!!�3����K���1<��@�v�v#��u�Fr�{smey��B����E���?�Ѿ��G�!}"ڐ��bDRp����W�
�ឈ8�
-Ôd�ߟ�>I��0��}ĥ���Z)���ۓRa]hpS���f�ƾA�5I+��eq���7��Eǆ�) ��jl�I�$��'�DU��EGF9�ף߬u�{��^2��j���`0�ڄ!��7�{`� N�����$#��\Ɲ�+�R3wIsm�iؚ6n�����l6�����$o������/Y���zL�" %F(�xE�OR��J����|�zq��NxD�`:'f�u�/D�jAo�_���$T�P)!�7۝�gmɔ̌	���ɡ�wܺ��㗯p`��zw��5��g'�Mymq���������긒�;&w��|�y�@�C�a�A�����������W� ���$���Rt̮BA�_���H���@���Ҭ�Nz��+ƕ?%����9�q*P[���|.��G���~G"�D�pO"*M�R�6�V�?U�8,Kx�'��(9_�ݐ�Wq�=A
q��;ǟP>a�M	�X�K: ��/z�Z;_E�x�J���v4؆t�-98���i�m�.h��5�����x��t��*���T��ڀ����e�p_������e���q����d�j��ߗr}�{�k�?�ǾP�'zUv÷d�Wi��V"�;Us������ o@yx�Mq��w���Q)������g���g��͑�33(����4���I�|c���[Á�//�-���t��V.H�M,�?���� @�_���"@�P�Q�FC8����ц��n�k�e	W��O.O�x}�k�_�W�HF���V�-;�h��v�r~\�'��rG?2�����x<V�yG��=�%�+�8]��
����,�������ߖ"�N�
b�'졉��5�6�O���P�]�ܱ���l��@ov�qX�� @u�)Z��4p���r��Y�D_)�F1���D,��3���h)�q����@��.L�S|r�΄x�jy?�$�u�ttZ;��'#��Q�h'�&��'U&n�Iy�F�.~���[\ܾ����Q�-?ӁK��U�,1�[��
>E�|Я	�4gX���i�a���Ƨ9�b!�;�0dr�N�>i���<2�QX���5���(���J�l�!ۛ9�H@G�M��q[bkV���+�Vj��
�/���\�n$E١YfE���D
��<�Op�V��u(�2�̇GU��>q_���AD�K�߷�H��|xQv:��vH��+�p�ϊ��HL�6Y|a�Ybs2GFM��˩Ͳ���*��؀��Q}VK׸��G�ax���8��̻j����M3)^��1U��)j��Eu4�i�� �����+�4%�۾}V�R���ӭ���&*���A�oB���˶��J1��W+�5���7ilBa}ԾFz�M�u`0��)=�T3F����t����u(u0�/����e�6�
r�vT�V<���T�\�o�^���r���0K���΅��
�����"1I�������'Ĭw�F~c�$�I�门�܈
�>�W���P' �S)��U7���},u�W��n8��Q�,'u��RĂ�р9��@W����;���*��(�B�u����y�,�j��ȳp�w��)*�)ѝ4%�Ѽ��S-��>��&�� �c ���֗KS�[�d��
����~z;�w^�xh��W�5RmE�\
@��1�V��l�۷_�Ƚ�M#f����B��0Z��f�e'&z��f^��,���)�xx��20��
ܚE����|u��Ap��"����L�ՠO��΍Em%��vH�	��� .y<�
������U��;����Y�l��V��*n(X����Ro�_D�٩�$U�-O�(Qj���q���D�d���Ut!�+�'S��2E"����N�����7\�,XN۳W�ɼ5���Lwvl����6�)�C~?i����ӣ��c��cVS��G�h�X���Yd���a���=���n�"e�p^D`ةx6vvP�7�^�x���ڋ_���:k�I5�X��f�^^T<dz�(�R��4O�����|/:w�6���O��}��@S�Ӕ����[8;���2�B�7�qa`��vtW�=�ِ��0��i��	
V�M#�3ẅ́fw+�W���U�J5K�+x�͸��6k�[R�g��]���<����"��������@�$��m'�s|\����^]��<�3�'0���y��O/sQP��u�P�,�&N-�������,�$�O��x���}�;����<�=_(f˰���7�Xܟ��6�~��
4����[�cһ���ySa����i�hL�A��eW���L���:NY���r85�ɠ�S0�:�{�X�#=dc��3�����AE�sq��.^��,�3��;G���.���m-S��f��Q�­��[V���ӬĐM�	�I������c���8�X|{�FT:]�}HE���p�Ugc��L�(i;h�:�xm��d�Tx����n�K��)RcgQT6����N\�\9��Dl"�ֳ���!�Tl�#X�A]�PuI<�Y�$#tYX
4��b@e��d��]\@�ʖ���_���1v-�h\�L2��C�ak���#]�Q�p�߯a���mjo��zX�2�d
���Q�Y�Y��%����e.}{oE�����ZV���!*W��M>��|�O}�0p���C�Z��7����w�j:2���,W������(��d|�<��彯g�l�O�.I�釂���K�U�_�lC�����Z��V%����{�Zip�����E=�Ӏ�I+={���JE��'�ы���؊�9�0g�fҀ_y�����Q�['qf8�r�RA��^�˫��f`�ݧ������-=ʮ%��8rm����,�åRW*�r�5��;�/7fBk�����fU3U�sc��f�*Ll�U\ u������d�v��5��'�qy�?)ːp���Cz�u)�Wq1�,�~� �b�����p��ic	9>�%D$v !m�>io.�YVC��ɋ���� ���ǽ'е�	 ���hR,ơ�!캌�&��"R��]j2��c��M��*�Gu �1R�-`���4��W�3�[�*�`f((B��0X�v<�g '��-X���tR�f��L	ó?:K�)��'��9H�3e#P�wa��-x@L�ed�a�_�;�����#�y��kH�]䘼;�x��tu�F���SO��-2�_Y	t�=��(��;2�ͽk?˴'rM-_WG_�CZ���ݟUŷ� ;|D�`vDI�h<�G��AN���Й�����0��(�z�q�_��!��6
I��=���BҔ2}+�>tf%u-���N���P"&��@"���/�萵&c���0�6A�, /�X��4�	��x6}˲=��x�˚~��5��U���������� ����j��t�������8^>�2�f���m��`�����~ͪ�
Y���W��u-�8�Bm`pH)n{�a��wݰ���֑{¿l�@b!.�{T@T�g��9r��8٬vJ��8�u���l�~3�P��=�
*�J*GB3Յ ��c����[!���gj�=Y�P���T�f��6�3L=��+�6�
��̊|�*�UԞjZ�?q��>G�a�g�}��_�(G�.��գ# �D��_�I���,=e���i|TK��N���d�O��P��i�$����}!t���ĭA�ȯ˄ �2vY��Je6��s�/͢d`��L��o8�~���I^����S=o�&h��[����Q@
2V�<��yʺoM��Yp��<��3SQ�ˁV��@�� b:���b���fXiT�1'��V~���<մ�C�z�ktE^�0��w}Yl�k<��S}����E@�2ow�7���� MF^��?��猫ķ��V��1Z��\L��~�����k���@�BN�?c}X�
U����n�K3Qv���*���	 a��6�̛sg�ԭ����%vy�k��f�L�,߷��+�)g��6L11;=R�}m��T0*Jd�UI���~�,���Ld��{k�o��+�u�m�/������}��k�^Oo�^�U*������ڍ"b��$Ow�R�]��$�J+���	�mL;0޵^L<��^|M�ى}$�Ǌ"�x��t`�I�E%M�j���ݐ���f>Q��
�42�T����:P��?h�h�xo۲T�O��ΉJSE�߲ϖ86@ӊ^º�8�V,!��[�1խ'ՕĢն�a1%����u��vۻ�t4|/�|��#�݄+M�l����dr�x����2l�0E;P�u���"�Yi[T�	4�Ԍ�k�('ʉ�M���t�g��p�>i��ÿ���˫5:��Xr|�.��;g�p�F���x��{[|m=�^e�璠�^�_q��h�g�.����= �*�/-�m��a�k�ߠJ�dרÅd���t��TzY�$�l��ޏ��1'ޝ��$��>�^Ql��Zπ�;��<?�66:0w�u�	��}s��Y>N��p�]"�UR��Z�3>�Z�z�`�޳b��:}�Ҫ�@5�C��S�kǨM��Bk����Wl�nF��5�C3ShV�S�6��.RF�憛���k�t�Pk�P>6�8u�}�C��$�4�y�e�N�O���)P�.��X �哥��=h�����D���q>$W'�C�x�\с �![��C%���|O��z�;Ə�{8�A,�@�°H�axd`��uNW�� �ş��{jt$Lӌ ���b��0:|��i��8)܉�k�D���U5���=�Ղ:�[[��M��-`�g�Jq��a�����D�ڇ%pr�%<g���,f�5Qx3��+3[]�eT �B�Nц~�_�2�lA�H�8�L�H�?���n���5<�~����4\�EU�Ń���;O�JS����X�5���Ђ�z�i�~�г�5Ff|�":y���Rlg��Y���h�g�T���������ͳ	&^�E�rjI���,[�������V!����Z�4��|�3���eQ�W��BR�9�M���d��x�~�{d2~�Cj�Pp���ˇP�i~3Q�)�N�2��n��%J� �,��Iuۊ,����� �����*q9�N�3��hRi4�V!8��;p�7����E�$���o�)������^e�7&+�NT��)��	鵫"������#W�XͶ�u���$���� W��P��<�#��xh��n*(H�=r�נPT�Fѡ
a񲀛���c�Dc���J���ƀl�j$pe^U)���ȯ�@��q�䧡���ގ ������BaZQf��(7m�k:��ش[<~����BvZD���cs��	&<�O�]�P��'��6ssBR�@�^�ˏB�� �������c�`va�x��_i�S꼗�"/q�>�����{�CQ�fx������L|���]j+f��|�=-j%�A��ϓ~�\�]Ӯ-�w�sI9��u/�B%����a�	�$̶K^i�5��ܓ�x+U��ǅ4n>�&� �j:�D3)2˦��9r���J~�j����*��\'�j�H��x��@�\D�C�}7�M�r0����?�&��2����^�PN7�6~���䅱 0�a¨_����ϸ1��]5y	�e���ʜ�n:�T*���V���~�mo��]3�S����
����!Y�׉,�����`3�)	�e���I.k�r�&3ukcO��5ʂ+>���
F��R���6��;V�g�˟�
SC� G�Pcd逘�#�j�Է@�̧��h��q��?��d	ї���ۈ�������uP8��F����p�vQB��v��nL6O��BoM�A���֓ S��XS޴�'�i� ��#�_�e��>�n@N�i8�^����Q���xh�>H�ʔ��v,��m��fW#`�ȅ��h�ణ��J�ɉu^_�`�y�z݂��Q�]\���m��#鿃��v��I9vʾ���&^a���%�^S��1p��U��`��>��ǝ�9=(d�N��s ����`���|���=g�tϒ���������|~C��+PZF9'��a��HT~(�39����i���b"*�˓ש����!�9�}TH�![��C]�Ϛ��]����F��y�G/�u�5YꉟPY���[R���M����v�ds|7�Q�@�MLBG �is�¢�H Xe"ӻUB6�Sd��P'����<{��,��>�M��C@��µI��2�@+g%��Kz ���:sY�~���⢱;HYU�V�6��}'@n Ox��a�~�F�`|�]K�ضS��ݼ@}�풷.���7�z3A@�~��,�g���Jq���8�������r�]��2�I\-���׈k����p��H����S,e�C��8L�;0��=W�:!-h�\�R���LߞQHʪtߕ����xc��,��e��cK���Ĩ�p=�)���� �BvOc;iCxS�L��;�np����+� ��+h�&R¹�<��W��.�W��.�6]&t�*��%�����{u�Ҳ�,L���22s���G ֚�������X��[�9��P��O�_�i[K"��4�u LZ�cѷ�;f+���C������w�Yo�F_.:@��I>įe��QՉS�.�nx�����K�<�;1}�f�1�G�,�����MX�j�GX��]T��ƣ�����W8����l������ZckMS!,�
j�2y�������v��%9_��S����n���|T�;��"��M>�w穆�z��wki�ۧ��2��4���>�e77��\&Ck{�@�pȬ��Ϩuc��T]*�V!��+�L֭��L����$��ĲS�J+q�YKW��(T:��F����
�?, �b��aIB����qKJ�r��p��e)�D)Ue��Iu�T��T�̄��	P��0@5��C\���oU��fQ�,h�ԼS�Hx4����k��ȿ,/�ag!խ,�p_���0���Ю~��{���=<3!��))�a�8��*H��h�4tvq@̑Ly9�l��d+��'%���D��
\����ox�j�8�2�G��A�f��o�+yE�� �s�<q,�m�u�gZ��:,N��ۀUC��U�����Q�ה�`\�+�O�wx���K �ާ�9^���*SWf-n�HHA��ܢd ��k4r
�����I���e�!5O�A�Mk�0m��;�F�zfo��f���&W<��3Ĺ���2T�&(ğX	x��I?�9G��uJ�]��ѹg{·�ư�­'�H	��o8���XT[���:�+�!�j!���MA��;�_���e�?2;"�y�D���0k�UI\e��Z�CPF´�ҍ�1��x�	��T�w�W0��h�8�/<s��KE��*,��F)N��v��ֶ��
�����̌�B�#\����*�����Y��Z����i{s�\�㙆;Z��"��@�?�<��Ǌ�ňy��ԧ���
"�����,+�;I�&��*��>+�䪑����fD�*qs6OҪ"*T�>H�9E�<�+aN}z��p��X��u�Q���l�R��$F��4a��s(a�}Zf��<�q�V4���CS(�ĖV3\o8}u��&��ܚ����N�$Z�� ��su�R��$d��߅�J�-��O�;�UT=m��nG�`#���Gd��(��"g��t�r`�{L @���u�s.���������z��t����i��vǄI+T?��� 8�����2]�2��a���~�� �r��?�%���`3���<͞@_���%�_�R�'��;Q	m�P��%������!1���QL�<'Wr��F/�Aԏ_*�U��"j�����X_�
�D��cC�@e�Pg�ps���3��J}#y�z�-<r����ԉ6-�d|�K��C�������Y��Dy�`��0���<u}?ʈO�FC�zXHо*>t7�}��4��/���=�o��_�T�Km�憕P�k�Od��xM���4�#-OG��j\��[_T|��l\�s%��Ӓ,��T��Z�y�������+��4[��(j����b[���{��k�^�|`Ξ�+��4܅�L�i9��20	0�鬜�9$��W0��88��Y9<�\<�`@S��
%t���T�A�E�����8��9ty5���]�S\.a�x-����2�ر��,�H��qUO�/�[��X�sD����_�Է�Xh�E���}_b!tOM����͢�I�Yu	��o� 1��WB�q7�b(�ѫō���m
O�c��gj��������9֘���ZƑw�B� ���-�jRv.��F-�?8�_��.؆FHq�t�T��D�~#TY(����[h?J�}���U$�=��r���� s��H���o;9��v�n#}�y䲹��5̅8���ؑ�G�������G���`�>z�~¥�_���U2S���\l�G�Xъ[��bQ[YV�3�=�!�PX1#�� ��}Y3����/$�̑����t���+d�(ρ���E�:k]�:O�wb�C�.���'���״�a}?�|�q
׽W�+��>m]N�Y~�*p� ��w���	$��]�q2�K��&,�YRg�w��J��6��L�L�����[f���@�X�'u��M���y�s��2�J1�9J��,�������U����np½D���ޜ�שnPǝ&�A�ebFe�)^�߱)fA��@u��_|�9�}|�o����=e�rMo쬶% {�ȡ�I���3HtĀ��ks��[]b�U�P�}�{Š4lb����`����*��G�����e`Ig��4��u��]!���v����>D��M��Y�z?���d;"<�� ��kW\oa?]Ȝ;���B&��Qy�ϔ�tȕ�/�h��� �x��8��R������ُfrD��&�*������H�
c }<]���Ӧ���$�j��4i�~�w#�I��3�d��89����]���!��U�������s��:�m��h�y^�]�i�\U}���%Y�j�Өٳ�n<G��$�JvX��f�@Y��	���2�b��mc�]��G�="K�9k�V5��¨A�[�ْu�`}?Sd�5i5"$�E����%�����Z:d�"N��mK*ï��X=�;�ͧ��_��5���*s@ꉢ�
@��h,�Y}Ag�vs}ܷ<=���f���bD��d:,�{��b޵����N���ƵQs������q�0S�Т5?����w@�Qv���}*i��J��Ɔ�m�-ǽ
�؋ۭ�t�ʰF��`���t�G�����2A���?�C�T�}�ω@q��,�uL�-�q.!�r���	�m�"��/p��a �;���RRyY�ί`ն��2C19��������M��歼�Btѡ�'ϋ�����\s�	l�(23����+��v_��E���
;���W�s����*>I?́{ӂW�d	�<�P��D�\���V��ͼ���,�n���i*3�j�]\��Y�[.Ut��W�
�0�mo̫)�������i%4ƫ�Yk;������і��[�,'t�TvF��g`���+S�n.��P����F�K�Wb���Y�Sv'���D�.�1�sK��� \���連z�*�f8h3�nw�����D%#�|9��:�%g=� 	����ot'm��SרL�#��s\b�Y�Ųt������zk���-n��g�B��G�q�x�	3�7������qW��/�C]����(wB�_�ƹ��Oqkφ�-Ol��vj���y�� �R�sv�:YS��
��9՘Pq�[<�J�b�>���:�s��G�fu">5�X���A�E�d��f qZ=E*��j�.����1*	�슑�T��L���E$���:s�n�MC,	l~�]j~b$_*<�Y�.g�;���GȀ 	�
ӂW<_D�# E}#=��1%X�
����Lp�Umr�F8̋HT��5z���q2W��1:��?����#V��d�y�l�L��A��v�ހ�
���I�S�9N��cό�D��N~�v�ʵzs������8�4��dY��5ˏNr�ș���H�$�n�C���Q�L&F�O~~���e.�;#������-�kd�Q9�&���Vw��}�g#���N��3���C%�GV3���`���Q�;|C���v�����]��H�"l��p�Cz�^�!X���ձ�y'�9�����eJ��X<;��v`�Á"�MZ@�9j �s��}8�yE3�Y)��BW�͖R/	x��B�p�c��u��T���"���V!� �˟��i�H��@������D�((!�7��tAO�P�o����w� s;��[�/���p��{�ay��F��V�\z�-e���} Nn�uh/ѧ�g�뀰�0�i闣`��::b�)H��� g��ʞ�����~0�4^���t9�a�U)�wj$r݌cՉ�K�FwwH ���<���p*�$�����d����a������"�2�n�AX�Y��l3������8O��n��#�͂�x�p�DAG�,xm��O
#{����k�W�O�*@��Qm�{�K�z3��ꚷ���,!�S�/�����I���ĂR$�3;2c�`��V��B�(`�{^�
D��S����G�^a�]�V���I�Ќv�C}���ca�M鳳Sԭc^�v�(i���Y��a+�����׉#�C��q�]]��x[����ϷъLD��m�~L��O���ݙ ����m��͸ʬ+��9�O�t|���K��A:���LҪ$��QQrp�Y&viV��]�U�z��G��ޟ�����M��'ك	,���5a���#�ҭ�	۟�N(�~hx�w����qLj[}��Bl���6m��I5���/��P�1U��N�D�l�υ��3��	 2d���2���@��!�/5iNp6(o�-jw8�ޅЀ�lbb;�R"����Q�C�pפ����c��gyF`�_)�-���	�~7�?�d���ܨ �j��m3���ū����ԓ��z�6G⥤{�pu� ����ȁ��g�L?��⹲U/�����;v�UJ�&���!�1ה���G:Tֵ_
	޸M�I|�_j��ҲU�g^�LW�����u�t��ӥ|1����!{��R�5����&���|��<!����;�К�'��q�S��/���.V [�S{P$����� _>PT_��r���5Q,:��6��A⵵�p��:���䀩��������y7���G��N2������̎^H�[\k�0�ծ�P������A��4.P��+f߈��n��|��S?�m��wd�b��v�n�C������(�pwR��&��?AH�à�v�%���".��9��x�q��JS>l�G� (�e�V�$��\��8y}�P5����C�$`*���;X����S�k�M�%�8�Xz�൤ޝe�(M@~Z�]D\����&tb�U����	H��`�?h����W�� l��R�Uf�.�b8�X��3V�XB\�<MF+c��rʍfg?M!��$����px �f^���5��X��
�nT \4Dl?�߲�b(x�%?��LH'-��Bkɦ��Q�,R��l��.)���wp�`��&;��C����Em'�U�\��,v�^�5ѠT/X�z��fc�Sk"���ݹ2}�|ꬿ-�Dg/+�Ꙇ�k5b�K��v�v�p̋���\�x�F���=�Ҽ�Gc�:�m3�>ŀ��Z�����Q�齥/Qx�'��Q#�v`�w�Y���O�.8�,_b��0�jY�|�g�nkܵD�\*0��M�KP+u�9�n��y��I��8�a4�<<�j�Ǽ}r�G0J�rt�?)���ޖ�Al�Z�]�u�z��eO<"H�l7Γ�L�El=jDq	��_��3 �D����Q)��Gm�����d���ЬTP���An'\D�� $�{����ؔ��3{�j�NS����y� S`�`���sPO�����^��	�6���^S�V�7�]y��^��3'�B���4$��K�K'��$NN`��{#�{���)�^T)�c Xt^���-M\8l�l��Z��� ���y��g�I��i��̍�t�~�K�U�=�g=!Ѭ�����53�'�����`���!rl�Ǯ�Z���[B�%ٍ+M'������=݈Օ�u���O���=��%Z��Ն���1�5FQ�M%M���!��$�OY�k�\�v���^�
�`"�F�mL�q�3o$�ev塯��)��2&��$I�}8�jh�����/��dY�:)x��M}2/ʚC	��������z96��%yA�U�Ve��y���#0�c?������L����#^����/��*h�S���«G���tN�����g��$�{�����oy��F->z���W	}�#��yQΥ��({��C�I�#�P�8�1�{UR�S�ˉ-{�YȲ/�2X�j�I ��B�S�%�`����*EB�n6KS��ɑ-;�1fͥ�A2�-�j���܉�e�!���E��*j���\�!`+H)���WI��(e	F	��������R	6!��Z��Iv[�����v��m%�/)�!iX�eT%��.���L����	N_�'2��_��#�sK�d��G�b�_����:m�&A�k��RE�y���͘�Z��\�hBs?#�4&��q0%G(Bp//����*�*Z��il�X'�09I۶�~�b����124 ��$�X��ڦ� ��)�<\F�z����IS�6�0�i?�fs��l�LQH
�\�s�n�+ m�M�d�Sj#�
�����]����`�ѼB~h��^�
�
k7��=HV�>u\����B^�^c=�eL�4������ Nls�n
�i�ȼ!��y����6kb�F�	0S�������X�W0�_�uiݷ"���O�	-A�.G��>�o/�!bD��Sª�s��Gld|�o'����izbf���w���pѴ/�y��$!]���T!����Hn�����/��ʴS�����s�9��9���I��N�$T6�	��*8�����H�)@Y(�6N"���f����
,�y��r��ͷX�����{P,�����
\�ށѢ���R�r^F�o�;r��e�V�����;	,�Zpg�^Du佹w#�0�޴��/��C��X���X�!'�n�;--�� -Ř��\%EH�����)���#r�0��|���T������&�YL�J;#�d'�.Q������c�\c��d�8���oT垷��|y!ѳ���#�-�㞂�G�k�χW���� ��ez2�G�&f��S+13,`Ŀ_M�)� ���A��F�ȹi��o�!��ŝjY���5e��tP�~���䰫sw�`t��&LXb����@a��5A8��fDhe���RL�A����@�]��J�>r\�z�m ��3{ءΔ[�%��O^�_]"�]>�v�R��q�`8�����`� �_�-$�iSh�Ӷv��V�qq"4QO�pO��!�*1W�: [r�v��N�D�BJ���q��/U��E�����J�x��1��@��d�3��%_y;�P�!�ey4]%��n�oF�DtsjZ�cX �?5����>���1� ��O/�a��DO���
A����D���i�s�ؓ�2yUT��8�{�\'���6�,̶#�岑���"����1���D*�o�s9��)ܯ}0Kw��$�1� ���@y�$�j8Jt6�N��zoH'P��?`�5��|�c��La�I$]�XA�<n\net�зȀ���_B�������Kӷ|	Y9kX�g�� �U�-����w������kQ��*	����u��� ��ы4lؘ�i1<U�`���.p���8�;���@��[�9X�����B�K]���th���.���;�uܗPL�}����ё��Y�(O(`ЎU ~��@ >K��
i�
���b|�+�g$rP�:��XI��!��2�@s]�=�W�L�VS�B�>Q,6�\�Pb�<#�q��� �i��\e5�O�湶��GP/"~�}�	� �H�FY�N����
��
A5=��!0<nZ��v�g�}/=j�l����Hss[��'CQ��Y:v4<����H�"?)J�!�bN�f���#�x��D�t�B��"��i���]�ƶ	�ʮ���h�ﶝ�J9�1��@Buz��2���G�v����転^ւ�A$�B�F��2]�B���18�ζ����}5V���H-�|J�v>�qB�\f�������- >��X��\4�>9�������1.�U=����7"�t�$*�Qϟ-�Gs���������Z��gq�b޻���У��!nqGxY\^�^��owf%Fx��pZ���*��Xj_\���qG�ɒ(N��s���bX^Օs�B �j?���a4�}�5S���[�������V�a^�1�6j�I3�|2c�#��_6Lg%����'p�|rz~��cy�����/���g���ɾo��V��Fn��/x~Wu�=ye(�̂��@�J��,y�F�iV�c@-4�>Mwh%5��OdPa�IE��w�$�2Ų�±k|�F�P��_7��� ݻk��X"G��T�i�#��+<�0�5���uB��s�a*�N�[N�u �L��W���̕\�k�W/,�����(:I�a�LKk�3���y6F�`�-���yaA�\�������#���@����򶚢͘lL&E���{, �2�D�dN���8K��)T�ϛ��}�xo�#���8 �LI{5�X_ʫ'�ё��	���h�r�|�2�a�����m� q�3��B�ˇ��?�.�jq�jZ����;���V�VV�������W����[/����R^�b�)Bi���@AU�JǸd ��A�B���7�U��ma�	�	q1� YL�di��K���cҚ��lCW��E�p��X,�/�`�����o�{уWڄQ�Q�ʯ�t���KO�w�v�"��<�+��SǾPFc~Fa�?z�Eͯ�d�G��H�hE�Ʃ5� �I�۷=�t���*4W��}�5Nˏ��n>a�����5R�-�k0m3�]��-��&�c�ˤJl�;7��7У]�M��d���"��Y�f��_8L�H��ol7`�:�U��0a�ɺ)s�.�L�s_1ϥ�[��(�FY�ZdK�[��-ym�Lj��ީ�pN�^�,1<c2�A={����3��R������磒b�˼�c ,�U�ͺ�O@�I=��V��9f��SÚ��2�b�,.����D�uD	��k�|vK�2��X��pk�`ZR�I���|/�y�+���܉-��UΒv��&@��b���(�ü+Ӹ^Ś��\K�i.9���$�E)���Ϣե:q��8�Z�YG�m�?��	�A]�d{V�Pg-�Z�=D��Y�h$X�A7�-d?,�{l`����7G�����]�6��5mH��y�[��7���f+���� ��b�5r|9�hGE���W��uF
�ӄ$��'�tVŎ�-�T��ԯx>I�R�Q�����^M;�綟AN.]���4�W�_t���\����C�s{�Ӗ8C��O�3�;A�0l����n�z 3��d�%e�W5*%S��-Eϑ�9�r�%%
�S�z�#�Py���	z:!sPrp�@�+���(>"�h�Q��3����������?��� 6_����ӽ�l��B"~�,kzč8�=A��|���)P�i1iT��3�hU7gܩ�3��);�S��X|Q��3��G�)�;k��]g�U�� �mZ���߳1�����J�|*���Ӧ�'��[yg��eQ�ܴ�M���C^�@�Rl�!��z��q�s\���.��%�)�#,e�R=�T�]��5���am�\�Ϗ��ݜ*���Kپg�i�38�����Ho���w�����_owOK6�Х�jT���\��mtk.����/l��\�����'�f�M����	��o�eQf�ZF)���M�X�d����I��ւ[����!/L��iR��[�@�P��t�j{00��>�I�P6���BF��`|t�LZ�U#�(��*�&����7F�`@���O���nH�Px�c����A
P�S�������u.��.��A;��������\�&Y7�E`��w�V�ݬ���KI`�e��]�u�b��q�:u��W�����]�2x�}�A߱Cݔ�(����zBN��つ�k����Ҋ��^Kh���	�x��������zR��ξ�F5[�	� g�l?"	�Bl;�f����m	�n�U���O{�o�K���W��Q��r����]��gd�F��L~�l����n�������kc�Q5�]�h���]�*E$�'}KO pO50�M���4m6-x<£��H<�YP�FF��T8�u�{%;��V6EVy=ٙ8�+�5�S��E�uH�y5x�~o�����G:��|W ���O�%�R >ͯZw?8i-�����ցX��빫/~V��t]�$Hk�r��75��_&�
yO�!�}�^*��R\c�)5g62��[�x���,AF=�J�,"�wnL9����x���C�*m<>F�ԟ�6�M}���F�%W�C��Ƭ��G.H��\�i�wwF��<&p�,}�����_�Z]ت�Sʾ��+���ּ�����x�"�H���D�P�-Zo��i~�9n�O<:�:���\q�+� ���}���x����ݟ�E+�
�Wͤb��[Ѹ/k�i�[@��e��ԑ,*q���y:̀�墈��ǚF)]�x�$ ��wV���������݈�u���q<���L��~�^��t
�#��=�3��j��[T�)y�I��|O�,֚���I��ٰ\͏��n��
]��䝷gvV��.O$�����"N^T���2ʘ��8�ǽ�ɤ�)Hs�	����ɷ���V��ݲA5S��ĸ����Bc���n:?���be G"aN-�m�ʦj�O�R��������	o����>�`l�G2�WQ_����_h����6h��4�{���dY=4��6���n�g�y�o�����d����R[w;���ԉO�9�ګ�?���� ^��D_���beI葲@Y���`�~bĲ0����b�T��d1�x�ZT��ļsF�=8
����ހ��5�^�Ԣ�>[
?�
J$����������w&kI`��.P����sHM��%�)�n�܏�%q'�,)�o�
�+e(�;q<���S;��3r�,CP�s+--?�i]��lW�^K��[�"A��=Qs������.R��T��K%!	��NY���؍��H] g�A�}��k�Yv�i�Dq��p��W�|�m�/�5�z�.q��Ŵ�3)�1������GvA���iꁾ�+�)�j���˳x���B�&���p�MEN��9��Y ޯ�X��w�A�Ҟ�-HB��p����<ׇc�4H���\��!^�FN�jL�Fl+υ� c�PQ��w����~�(��-��?�@`�����N@&��w��U�	G{a3���)����#G�Әه1���B�?�Q�*�L���n]�X�0'Yt\�p��Cw�M_"<;�=��p�����I6:ИgG��[�UN3w��E�6��}
 aȵ�߫�|]�����Y|�RO6cV��0�_/���`����=�0�A�kd���b��� =.U�
�C"j̻���x6jv�],����l�B��`3���ۍ��������r�x��j���4���LcRa�:�iѮ5p&I/ԒE՞�S�2�q5�����0�`��q4�5�sa����n 0)�2�SX�&�}ttcí�?���$ϡR�'k��㇦���ǵh1_z�I����Hw����D�6c+���O��(	�����R (9Px��v��^��ч�.v�h��kS�����e��P#^^�.2д5ԣ֛uUc� 4s���N;R��`�n�	��ړ�۸%�B+�EBIT]��˼��Х's`���uom�Au~�o�d�涏f(�n���o+�ь�L�,m,�����i��8°��z`m]3�	�����3n���+j�(n�+�5������z���S�@�nΌsP�}cqf�����!i���Z�G| �>�=��*p�bG?�(t�<K�=�V�έʹ����F@�֪L��(:տ�����eYd|��=��1�2���>�ĸ��?� #�ϩӻG���]�JZ�L4�f��(6҉G_�hK��L �a�}��}O�:��b(`��=�y)���my�h�������ژ)����i����Ŭ^������re!��t�����k?��'�aǯ8w9�;]A��{�`!��=m�xm=WB�q+�,+ssڍq���'i҅��3�?O�����e�j�[cׄ�g��i��4Wuck�	l��mB��4�� ���5O�֛-��
ϕ�	Rӏ���4�����.��x�G5��.�fl ��j��6� .{�D����니-*�ǂ�W�U|����Z; �LȰ�H|��pveS޴��g��M���\B=��P�'�֭�U�>&�䋒����'m��I�8��F4@0�|��)TL������ʖ��Yqn���m�LޡgGMo_�Lw��	Փ�-�~8}��/����� Fz��)&�^�'�����@���5��e���2/��*�~��w()�4P?��EϿ#�x�!���a�֬&��8�hr����p�O��攥��>	js@�0�Y(�[�[3��>Q�^&��'��5��8�j��q�Nif��:�$�xZ1oe�[��ց�GkL��7j���5��_X��\T �V*H=d��:����x	F͢��vu��sƈ����f��B�"Jl �E2'V��տ�F�������[A�fY�Y��s�Ȫ_[<�鑣ϟ�-��|H��z~��Qm.W��2\*5�Qe�"�kx�:���_��	/�HX�q���v<�r4��lj�.���p��&@��5�~����(r�WT�7Νu��*��8Ԋp��?U[�p��=��)1��{���Ϊ��D�4����˭赂zR�!ޕ0Z���׌���y�l�,�9kCC���b����n<<��p��L�h'z��m���k�E�wN