��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� 8P�?�bj���H��G���+'���3�lUK���?�>SJCu:���A��:�Q)s�.��H���>�j�<I��Ef?����3�"x�lc�P#'�1;�B�h`�H}H|��ɋ#U�)ļ�MY�?�3�J\��и�ȯ�Rb�#w:��c����~��*`z�Ui��i�b/p;KK����∋MgT�����T-5AA���Y�J?�� 1m��N,�=6r�΍���RC5�|�鄻���ݡ�f��eA����zt��6	W���)�%s��n�#[e�k�ÐL��݊�-�9�3��s�=����c������q!��͖
e$h#��˚J����v��qL
4�O�UiT��2���B͒����ZNK�R��Zl��Y�o4P]���,�|�n��w�{�&�D���Re��N�� 0�ۖ�sJ��?k�؇��!)'	&�K˜\(��xM�G|��+	�,֦[�IsZ#���Xnn�mnJ�i�
�5i�?�(|G�L�A^���U�Jm�V45�<�]2��6�=n(Չj�ʡ1u(ϊ=�u��ӄ������c��}���C{B$A���|�
���$��!Ұ�Tؖܭ�"�**@N͜���c�}%��l�غ>�i�1��<����/l�}7 ��b[�%:�`�\���lj�8��E�b=��E�+�H��gJ�0B/�F�rU��z5U��P�4�c{����	�[�OHJ��@Xg�av;�l�u�du��b��C^����A�g���,r�Q��L�O�g�#xp���v�MdF����2��a`��X���^_A�6��S�S���y�Gn-��4D�ӌG�z�^�~����C�:bއ�1���@C�I��N�pptO�Lͳ�@%I�/�Bx�\��x�`,�ئvO���mE�Q:���v��@�M��M��DY�Os�H�v�dT��4�j��o�s������%.���=��Fk��K���e��k����F�C�rʆ&���FT�Na^�hi_�i���HHo��Q�R oj]E���Sꋅ�!O,N��䬘��$)��z���(P�?	���;��gI��o��C	,"��T�H�Wo9���a(��İ@{��nM�K�$�4�g&�Z=/�yP>�M��2�!�v���>#V�(���n�l-VAé���?Q>�u�qŘ�Y	�9�^��{
]�5Vc��(��Ա��*�Z4s�)�GaJDa�|�e�?����57�]&�[*�|�B��/��p1g�Ki�bQuDnL$	vG�*�Ξ$��\��$�Td�4����0O��t0{ �cK�`74z���K�>(������1Tm�4�U��gM�_e��Sb� ڶ���k�N������j�Y%8�c�%*���|C*X	�uI���_�i�P�����r��ohaxB��
f����l,�khX���}J�պ/� 8����l�CjӜ���������7�z"�]���?~���%����w$@H�qv}�R��5A	eXS2$û��F$T�RB��ͩ�h�|�P��1tdC.��\�oM��3_ę 17�cΈ����R��[��[�0R�T-�M���2h�Q��v���=lt~���-,
�m(��>"@���GT5 UTD��+O^�"}�>�	�M�E��-7���kŹ*���`/�����'E+��33D�\*��O\˭��M}�ֳ�˅,�,\��De;=$01s^����:�ߥ=��[XB���ϗ�!X�:����g�8��\X�g�{\u�
�<\S��>
����ӒF]Ei�:vN�����ֶ��nNڷ����r��c~���抇�9�d�9��d����UKy{��"�mX�N��@#���ǎ��)Dљ�fW����oyC� �a}1���9�`fvK� ���&Z���'!�jw���۟ū���,�E���[b�V5���Х��Bsxђ��kaw�	5�l�ט47���s��R�0A>�U��j�²��rx	C��d�[�@c�S���b:��`ٚ�7�HsA�����g���w�g�놦����"�T
ݒ���}�gEb)Q>/�� �W��5�o"��&/�����Jn��!68��s����"W�gT��ڟ�J
�B
�Hn��	�}��R�M�H�-�+�򒛑����-��S�uD�� �8Tk��1����ꖥ�Ў���/^�^ղ����T:8il��s-o�!?o�d� �Ϫ!F���F*���q���J���k�3����=���h�!��7V���S�R�ӷ�_4C�
<��t�b��Ui������8.��TV��0���=ߋ_V�����h�?w����/^Z��-b뀚뛽K�����F	�_��\��bAº�1���k��h��	��5���t�J����Ǉ����	��Ie;6FN�Z��0����C��7�7�Y���4�O@�6*�������W�}�Y-�ǥ	��*��z�Rdb{|���H`�Á�WR����m �L��|ۆ#Q54�6����u�y��s%��&�d�Jȩ<��Y��,�̶<^u	���@�� ��$Db��h;GC5w�ڭ��~�g�ws)�������45�x�����F渚�B���% �	��eⴔR�mq�`G���n������u�b�Z�r�/&�26��h����FQ��I�X5C`���{�E�ʷ�!�B��%��_�%`�臤t~���<��^��V`�p���<���Ѐ� LQ����O�d�5	�a���p��!���\5+��F����Lbt@��Aa�+;���IW\W;�P�6Ӟۄ_�p������v¿����Ҁ��5�k��ó�����N�F�酇gbd��Uk�-NX��n(4!�l}H�<`9b�1S��4PO�	�O�fV2z�p��wMI�g����*�9x`Sͱ����ɽ�^�O,�����6GL�	���[o�o�E]D��A�#n�
2�!%N]�_���`?���uH-ӳ�|��� <��F@Ǌ��a"�|�q�6�D���3n�[Q�R���7��؟��mxHxPQV5�,o;��զ���Y^�B��m�٨�+��o�7���݌�z���ȫ�'E"7� ���&��
�0����g�<��Biӛ�#B�=��_�,�+���/P�{��fPp=0����Uiޛ5Aњ������8�����_s�H,�Jَ�ϋ����͆H���M؛�ѯ+�k�:I�q���)����=R�PB)���ĺ�����T�2Y%��Gb����ݨ5C�%���*�S����d��H�P�E�qaK���֒����%�2ٽ�cK���
�X��?5R�LNYq�n�1��ģ݊�}y?�>��(�r��z�b :��Z��E�6��@y**���TM�2�^�&�
�Ԩف�:����iƻ�Ao���t�ן�Á����n҄a��۪>�~�\�u��Q�#M�W��ֻ�%�%d�hpe�f���$vfj;�dZx��c���11�
(0�]v/_^V��zGm�sH;)����vsP�E�	D���Z���J7�Y�~!ӱ_ 2���#���^ځ,U�kw=ߑ�L���!-%g�Q��O�Ҩ�D�e��;V�.�m<��VF�	W&�勤I�c��`�#i!���:������M��U;)�,f�g:��u}����ڕ��b�,5���Pe:�����:K��&;��F�g�,�zMO�)Ww������������L[J�@�4_b�=���ܒ)��]0޼��i���0E�u������;��eJ0M�2�{��u�Q�$1h�o��aj�=���(\�9>��I!���`��a��j���U/�O���Ed
N�����g}g+����ʚ�	���)r�S�i�K@ی���49ތ�<3�W��⫈38W��s�l������x��d<gѥ�"Xz[y̺�|t�Љ��I[�m�P1]�Ī��R�b３�R�i�߰�2� �hY\�9�(x���
,�A�Wx��8��|��,�>d}�bo
��7�G���L�� �]�4yή�u��}!p��T�<�dk�ɱU�C/��Ɓ13����l�kV����C�S� ���(H��ŲV����ft`���x]�Mn�}Jᡪ�f>˦"l�A�*1� k�%�4bL�̀���h*۸gN��|�vn��i�\�ϝ����c���'����<�*=q�Z ĎV��q�՚mf�l�r_���"5Xd�dO���0��L�E�(�VTvA'j���v����9���C"���7=Eu���g��(�w���Y��
q��`~�.<'p�0\��e;y=1-̋\g� �H\NYfr��m��ID�''f}Y����隈�"�aQ �m�A�a3�ctS����&a{�?D�7^�m�y2hIV�fd��ц���9'sE�
��E���|
�G��$�o8�<�#*.2K#V�;e